`ifndef BSG_DEFINES_V
`define BSG_DEFINES_V

`define BSG_MAX(x,y) (((x)>(y)) ? (x) : (y))
`define BSG_MIN(x,y) (((x)<(y)) ? (x) : (y))

`define BSG_SIGN_EXTEND(sig, width) \
  ({{`BSG_MAX(width-$bits(sig),0){sig[$bits(sig)-1]}}, sig[0+:`BSG_MIN(width, $bits(sig))]})
`define BSG_ZERO_EXTEND(sig, width) \
  ({{`BSG_MAX(width-$bits(sig),0){1'b0}}, sig[0+:`BSG_MIN(width, $bits(sig))]})

// place this macro at the end of a verilog module file if that module has invalid parameters
// that must be specified by the user. this will prevent that module from becoming a top-level
// module per the discussion here: https://github.com/SymbiFlow/sv-tests/issues/1160 and the
// SystemVerilog Standard

//    "Top-level modules are modules that are included in the SystemVerilog
//    source text, but do not appear in any module instantiation statement, as
//    described in 23.3.2. This applies even if the module instantiation appears
//    in a generate block that is not itself instantiated (see 27.3). A design
//    shall contain at least one top-level module. A top-level module is
//    implicitly instantiated once, and its instance name is the same as the
//    module name. Such an instance is called a top-level instance."
//  

`define BSG_ABSTRACT_MODULE(fn) \
    /*verilator lint_off DECLFILENAME*/ \
    /*verilator lint_off PINMISSING*/ \
    module fn``__abstract(); if (0) begin : abstract fn not_used(); end endmodule \
    /*verilator lint_on PINMISSING*/ \
    /*verilator lint_on DECLFILENAME*/

// macro for defining invalid parameter; with the abstract module declaration
// it should be sufficient to omit the "inv" but we include this for tool portability
// if later we find that all tools are compatible, we can remove the use of this from BaseJump STL

`ifdef XCELIUM // Bare default parameters are incompatible as of 20.09.012
               // = "inv" causes type inference mismatch as of 20.09.012
`define BSG_INV_PARAM(param) param = -1
`elsif YOSYS // Bare default parameters are incompatible as of 0.9
`define BSG_INV_PARAM(param) param = "inv"
`else // VIVADO, DC, VERILATOR, GENUS, SURELOG
`define BSG_INV_PARAM(param) param
`endif


// maps 1 --> 1 instead of to 0
`define BSG_SAFE_CLOG2(x) ( (((x)==1) || ((x)==0))? 1 : $clog2((x)))
`define BSG_IS_POW2(x) ( (1 << $clog2(x)) == (x))
`define BSG_WIDTH(x) ($clog2(x+1))
`define BSG_SAFE_MINUS(x, y) (((x)<(y))) ? 0 : ((x)-(y))

// calculate ceil(x/y) 
`define BSG_CDIV(x,y) (((x)+(y)-1)/(y))

`ifdef SYNTHESIS
`define BSG_UNDEFINED_IN_SIM(val) (val)
`else
`define BSG_UNDEFINED_IN_SIM(val) ('X)
`endif

`ifdef VERILATOR
`define BSG_HIDE_FROM_VERILATOR(val)
`else
`define BSG_HIDE_FROM_VERILATOR(val) val
`endif

`ifdef SYNTHESIS
`define BSG_DISCONNECTED_IN_SIM(val) (val)
`elsif VERILATOR
`define BSG_DISCONNECTED_IN_SIM(val) (val)
`else
`define BSG_DISCONNECTED_IN_SIM(val) ('z)
`endif

// Ufortunately per the Xilinx forums, Xilinx does not define
// any variable that indicates that Vivado Synthesis is running
// so as a result we identify Vivado merely as the exclusion of
// Synopsys Design Compiler (DC). Support beyond DC and Vivado
// will require modification of this macro.

`ifdef SYNTHESIS
  `ifdef DC
  `define BSG_VIVADO_SYNTH_FAILS
  `elsif CDS_TOOL_DEFINE
  `define BSG_VIVADO_SYNTH_FAILS
  `elsif SURELOG
  `define BSG_VIVADO_SYNTH_FAILS
  `elsif YOSYS
  `define BSG_VIVADO_SYNTH_FAILS
  `else
  `define BSG_VIVADO_SYNTH_FAILS this_module_is_not_synthesizeable_in_vivado
  `endif
`else
`define BSG_VIVADO_SYNTH_FAILS
`endif

// macro for denoting that a code snippet is unsynthesiable

`ifdef SYNTHESIS
  `define BSG_HIDE_FROM_SYNTHESIS
`endif

`define BSG_STRINGIFY(x) `"x`"


// For the modules that must be hardened, add this macro at the top.
`ifdef SYNTHESIS
`define BSG_SYNTH_MUST_HARDEN this_module_must_be_hardened
`else
`define BSG_SYNTH_MUST_HARDEN
`endif


// using C-style shifts instead of a[i] allows the parameter of BSG_GET_BIT to be a parameter subrange                                                                                                                                                                               
// e.g., parameter[4:1][1], which DC 2016.12 does not allow                                                                                                                                                                                                                          

`define BSG_GET_BIT(X,NUM) (((X)>>(NUM))&1'b1)

// This version of countones works in synthesis, but only up to 64 bits                                                                                                                                                                                                              
// we do a funny thing where we propagate X's in simulation if it is more than 64 bits                                                                                                                                                                                               
// and in synthesis, go ahead and ignore the high bits                                                                                                                                                                      

`define BSG_COUNTONES_SYNTH(y) (($bits(y) < 65) ? 1'b0 : `BSG_UNDEFINED_IN_SIM(1'b0)) + (`BSG_GET_BIT(y,0) +`BSG_GET_BIT(y,1) +`BSG_GET_BIT(y,2) +`BSG_GET_BIT(y,3) +`BSG_GET_BIT(y,4) +`BSG_GET_BIT(y,5) +`BSG_GET_BIT(y,6)+`BSG_GET_BIT(y,7) +`BSG_GET_BIT(y,8)+`BSG_GET_BIT(y,9) \
                                                                                       +`BSG_GET_BIT(y,10)+`BSG_GET_BIT(y,11)+`BSG_GET_BIT(y,12)+`BSG_GET_BIT(y,13)+`BSG_GET_BIT(y,14)+`BSG_GET_BIT(y,15)+`BSG_GET_BIT(y,16)+`BSG_GET_BIT(y,17)+`BSG_GET_BIT(y,18)+`BSG_GET_BIT(y,19) \
                                                                                       +`BSG_GET_BIT(y,20)+`BSG_GET_BIT(y,21)+`BSG_GET_BIT(y,22)+`BSG_GET_BIT(y,23)+`BSG_GET_BIT(y,24)+`BSG_GET_BIT(y,25)+`BSG_GET_BIT(y,26)+`BSG_GET_BIT(y,27)+`BSG_GET_BIT(y,28)+`BSG_GET_BIT(y,29) \
                                                                                       +`BSG_GET_BIT(y,30)+`BSG_GET_BIT(y,31)+`BSG_GET_BIT(y,32)+`BSG_GET_BIT(y,33)+`BSG_GET_BIT(y,34)+`BSG_GET_BIT(y,35)+`BSG_GET_BIT(y,36)+`BSG_GET_BIT(y,37)+`BSG_GET_BIT(y,38)+`BSG_GET_BIT(y,39) \
                                                                                       +`BSG_GET_BIT(y,40)+`BSG_GET_BIT(y,41)+`BSG_GET_BIT(y,42)+`BSG_GET_BIT(y,43)+`BSG_GET_BIT(y,44)+`BSG_GET_BIT(y,45)+`BSG_GET_BIT(y,46)+`BSG_GET_BIT(y,47)+`BSG_GET_BIT(y,48)+`BSG_GET_BIT(y,49) \
                                                                                       +`BSG_GET_BIT(y,50)+`BSG_GET_BIT(y,51)+`BSG_GET_BIT(y,52)+`BSG_GET_BIT(y,53)+`BSG_GET_BIT(y,54)+`BSG_GET_BIT(y,55)+`BSG_GET_BIT(y,56)+`BSG_GET_BIT(y,57)+`BSG_GET_BIT(y,58)+`BSG_GET_BIT(y,59) \
                                                                                       +`BSG_GET_BIT(y,60)+`BSG_GET_BIT(y,61)+`BSG_GET_BIT(y,62)+`BSG_GET_BIT(y,63))

// nullify rpgroups
`ifndef rpgroup
`define rpgroup(x)
`endif

// verilog preprocessing -> if defined(A) && defined(B) then define C
`define BSG_DEFIF_A_AND_B(A,B,C) \
    `undef C \
    `ifdef A \
        `ifdef B \
            `define C \
        `endif \
    `endif

// verilog preprocessing -> if defined(A) && !defined(B) then define C
`define BSG_DEFIF_A_AND_NOT_B(A,B,C) \
    `undef C \
    `ifdef A \
        `ifndef B \
            `define C \
        `endif \
    `endif

// verilog preprocessing -> if !defined(A) && defined(B) then define C
`define BSG_DEFIF_NOT_A_AND_B(A,B,C) `BSG_DEFIF_A_AND_NOT_B(B,A,C)

// verilog preprocessing -> if !defined(A) && !defined(B) then define C
`define BSG_DEFIF_NOT_A_AND_NOT_B(A,B,C) \
    `undef C \
    `ifndef A \
        `ifndef B \
            `define C \
        `endif \
    `endif

// verilog preprocessing -> if defined(A) || defined(B) then define C
`define BSG_DEFIF_A_OR_B(A,B,C) \
    `undef C \
    `ifdef A \
        `define C \
    `endif \
    `ifdef B \
        `define C \
    `endif

// verilog preprocessing -> if defined(A) || !defined(B) then define C
`define BSG_DEFIF_A_OR_NOT_B(A,B,C) \
    `undef C \
    `ifdef A \
        `define C \
    `endif \
    `ifndef B \
        `define C \
    `endif

// verilog preprocessing -> if !defined(A) || defined(B) then define C
`define BSG_DEFIF_NOT_A_OR_B(A,B,C) `BSG_DEFIF_A_OR_NOT_B(B,A,C)

// verilog preprocessing -> if !defined(A) || !defined(B) then define C
`define BSG_DEFIF_NOT_A_OR_NOT_B(A,B,C) \
    `undef C \
    `ifndef A \
        `define C \
    `endif \
    `ifndef B \
        `define C \
    `endif

`endif
// MBT 7/7/2016
//
// 1 read-port, 1 write-port ram
//
// reads are synchronous
//
// NOTE: Users of BaseJump STL should not instantiate this module directly
// they should use bsg_mem_1r1w_sync_mask_write_bit.


//`include "bsg_defines.sv"

module bsg_mem_1r1w_sync_mask_write_bit_synth #(parameter `BSG_INV_PARAM(width_p)
						, parameter `BSG_INV_PARAM(els_p)
						, parameter read_write_same_addr_p=0
						, parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
                                                , parameter latch_last_read_p=0
                                                , parameter disable_collision_warning_p=1
                                        )
   (input   clk_i
    , input reset_i

    , input                     w_v_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0]       w_mask_i
    , input [addr_width_lp-1:0] w_addr_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0]       w_data_i

    // currently unused
    , input                      r_v_i
    , input [addr_width_lp-1:0]  r_addr_i

    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r_data_o
    );

   wire                   unused = reset_i;

   if (width_p == 0)
    begin: z
      wire unused0 = &{clk_i, w_v_i, w_mask_i, w_addr_i, r_v_i, r_addr_i};
      assign r_data_o = '0;
    end
   else
    begin: nz

   logic [width_p-1:0]    mem [els_p-1:0];
   logic read_en;
   logic [width_p-1:0] data_out;

   // this treats the ram as an array of registers for which the
   // read addr is latched on the clock, the write
   // is done on the clock edge, and actually multiplexing
   // of the registers for reading is done after the clock edge.

   // logically, this means that reads happen in time after
   // the writes, and "simultaneous" reads and writes to the
   // register file are allowed -- IF read_write_same_addr is set.

   // note that this behavior is generally incompatible with
   // hardened 1r1w rams, so it's better not to take advantage
   // of it if not necessary

   // we explicitly 'X out the read address if valid is not set
   // to avoid accidental use of data when the valid signal was not
   // asserted. without this, the output of the register file would
   // "auto-update" based on new writes to the ram, a spooky behavior
   // that would never correspond to that of a hardened ram.

   logic [addr_width_lp-1:0] r_addr_r;

   assign read_en = r_v_i;
   assign data_out = mem[r_addr_r];


   always_ff @(posedge clk_i)
     begin
        if (r_v_i)
          r_addr_r <= r_addr_i;

`ifndef BSG_HIDE_FROM_SYNTHESIS
        else
          r_addr_r <= 'X;

        // if addresses match and this is forbidden, then nuke the read address

        if (r_addr_i == w_addr_i && w_v_i && r_v_i && !read_write_same_addr_p)
          begin
             if (!disable_collision_warning_p)
               begin
                 $error("X'ing matched read address %x (%m)",r_addr_i);
               end
             r_addr_r <= 'X;
          end
`endif

     end

  if (latch_last_read_p)
    begin: llr
      logic read_en_r; 

      bsg_dff #(
        .width_p(1)
      ) read_en_dff (
        .clk_i(clk_i)
        ,.data_i(read_en)
        ,.data_o(read_en_r)
      );

      bsg_dff_en_bypass #(
        .width_p(width_p)
      ) dff_bypass (
        .clk_i(clk_i)
        ,.en_i(read_en_r)
        ,.data_i(data_out)
        ,.data_o(r_data_o)
      );
    end
  else
    begin: no_llr
      assign r_data_o = data_out;
    end

   genvar                       i;
   for (i = 0; i < width_p; i=i+1)
     begin
	always_ff @(posedge clk_i)

	  if (w_v_i && w_mask_i[i])
            mem[w_addr_i][i] <= w_data_i[i];
     end
  end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_1r1w_sync_mask_write_bit_synth)
// MBT 7/7/2016
//
// 1 read-port, 1 write-port ram
//
// reads are synchronous
//
// NOTE: Users of BaseJump STL should not instantiate this module directly
// they should use bsg_mem_1r1w_sync_mask_write_bit.


//`include "bsg_defines.sv"

module bsg_mem_1r1w_sync_mask_write_byte_synth #(parameter `BSG_INV_PARAM(width_p)
						, parameter `BSG_INV_PARAM(els_p)
						, parameter read_write_same_addr_p=0
						, parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
                                                , parameter latch_last_read_p=0
                                                , parameter write_mask_width_lp = width_p>>3
						, parameter harden_p=0
                                                , parameter disable_collision_warning_p=1
                                        )
   (input   clk_i
    , input reset_i

    , input                     w_v_i
    // for each bit set in the mask, a byte is written
    , input [`BSG_SAFE_MINUS(write_mask_width_lp, 1):0] w_mask_i
    , input [addr_width_lp-1:0] w_addr_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0]       w_data_i

    // currently unused
    , input                      r_v_i
    , input [addr_width_lp-1:0]  r_addr_i

    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r_data_o
    );

   wire                   unused = reset_i;

   if (width_p == 0)
    begin: z
      wire unused0 = &{clk_i, w_v_i, w_mask_i, w_addr_i, r_v_i, r_addr_i};
      assign r_data_o = '0;
    end
   else
    begin: nz

  for(genvar i=0; i<write_mask_width_lp; i=i+1)
  begin: bk
    bsg_mem_1r1w_sync #( .width_p      (8)
                        ,.els_p        (els_p)
                        ,.addr_width_lp(addr_width_lp)
                        ,.latch_last_read_p(latch_last_read_p)
			,.verbose_if_synth_p(0) // don't print out details of ram if breaks into synth srams
                      ) mem_1r1w_sync
                      ( .clk_i  (clk_i)
                       ,.reset_i(reset_i)
                       ,.w_v_i    (w_v_i & w_mask_i[i])
                       ,.w_data_i (w_data_i[(i*8)+:8])
                       ,.w_addr_i (w_addr_i)
                       ,.r_v_i    (r_v_i)
                       ,.r_addr_i (r_addr_i)
                       ,.r_data_o (r_data_o[(i*8)+:8])
                      );
  end
   end

endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_1r1w_sync_mask_write_byte_synth)

// MBT 7/7/2016
//
// 1 read-port, 1 write-port ram
//
// reads are synchronous
//
// although we could merge this with normal bsg_mem_1r1w
// and select with a parameter, we do not do this because
// it's typically a very big change to the instantiating code
// to move to/from sync/async, and we want to reflect this.
//
// NOTE: Users of BaseJump STL should not instantiate this module directly
// they should use bsg_mem_1r1w_sync.

//`include "bsg_defines.sv"

module bsg_mem_1r1w_sync_synth #(parameter `BSG_INV_PARAM(width_p)
				 , parameter `BSG_INV_PARAM(els_p)
				 , parameter read_write_same_addr_p=0
				 , parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
                                 , parameter latch_last_read_p=0
                 , parameter verbose_p=1
				 )
   (input   clk_i
    , input reset_i

    , input                     w_v_i
    , input [addr_width_lp-1:0] w_addr_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0]       w_data_i

    // currently unused
    , input                      r_v_i
    , input [addr_width_lp-1:0]  r_addr_i

    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r_data_o
    );

   wire                   unused = reset_i;

   if (width_p == 0 || els_p == 0)
    begin: z
      wire unused0 = &{clk_i, w_v_i, w_addr_i, r_v_i, r_addr_i};
      assign r_data_o = '0;
    end
   else
    begin: nz

   logic [width_p-1:0]    mem [els_p-1:0];
   logic read_en;
   logic [width_p-1:0] data_out;

   // this treats the ram as an array of registers for which the
   // read addr is latched on the clock, the write
   // is done on the clock edge, and actually multiplexing
   // of the registers for reading is done after the clock edge.

   // logically, this means that reads happen in time after
   // the writes, and "simultaneous" reads and writes to the
   // register file are allowed -- IF read_write_same_addr is set.

   // note that this behavior is generally incompatible with
   // hardened 1r1w rams, so it's better not to take advantage
   // of it if not necessary

   // we explicitly 'X out the read address if valid is not set
   // to avoid accidental use of data when the valid signal was not
   // asserted. without this, the output of the register file would
   // "auto-update" based on new writes to the ram, a spooky behavior
   // that would never correspond to that of a hardened ram.

   logic [addr_width_lp-1:0] r_addr_r;
   wire [addr_width_lp-1:0] r_addr_li = (els_p > 1) ? r_addr_i:'0;
   wire [addr_width_lp-1:0] w_addr_li = (els_p > 1) ? w_addr_i:'0;

   assign read_en = r_v_i;
   assign data_out = mem[r_addr_r];

   always_ff @(posedge clk_i)
     if (r_v_i)
       r_addr_r <= r_addr_li;
     else
       r_addr_r <= 'X;

  if (latch_last_read_p)
    begin: llr
      logic read_en_r; 

      bsg_dff #(
        .width_p(1)
      ) read_en_dff (
        .clk_i(clk_i)
        ,.data_i(read_en)
        ,.data_o(read_en_r)
      );

      bsg_dff_en_bypass #(
        .width_p(width_p)
      ) dff_bypass (
        .clk_i(clk_i)
        ,.en_i(read_en_r)
        ,.data_i(data_out)
        ,.data_o(r_data_o)
      );
    end
  else
    begin: no_llr
      assign r_data_o = data_out;
    end

   always_ff @(posedge clk_i)
     if (w_v_i)
       mem[w_addr_li] <= w_data_i;

   end

`ifndef BSG_HIDE_FROM_SYNTHESIS
   initial
     begin
        if (verbose_p)
      $display("## %L: instantiating width_p=%d, els_p=%d (%m)",width_p,els_p);
     end
`endif

endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_1r1w_sync_synth)// MBT
//
// 1 read-port, 1 write-port ram
//
// reads are asynchronous
//
// for synthesizable internal version, we omit assertions
// these should be placed in the outer wrapper
//

//`include "bsg_defines.sv"

module bsg_mem_1r1w_synth #(parameter `BSG_INV_PARAM(width_p)
			    ,parameter `BSG_INV_PARAM(els_p)
			    ,parameter read_write_same_addr_p=0
			    ,parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p))
(
  input w_clk_i
  ,input w_reset_i

  ,input w_v_i
  ,input [addr_width_lp-1:0] w_addr_i
  ,input [`BSG_SAFE_MINUS(width_p, 1):0] w_data_i

  // currently unused
  ,input r_v_i
  ,input [addr_width_lp-1:0]  r_addr_i

  ,output logic [`BSG_SAFE_MINUS(width_p, 1):0] r_data_o
);

  wire unused0 = w_reset_i;
  wire unused1 = r_v_i;

  if (width_p == 0 || els_p == 0)
   begin: z
     wire unused2 = &{w_clk_i, w_addr_i, w_data_i, r_addr_i};
     assign r_data_o = '0;
   end
  else
   begin: nz

  logic [width_p-1:0] mem [els_p-1:0];

  wire [addr_width_lp-1:0] r_addr_li = (els_p > 0) ? r_addr_i:'0;
  wire [addr_width_lp-1:0] w_addr_li = (els_p > 0) ? w_addr_i:'0;

  // this implementation ignores the r_v_i
  assign r_data_o = mem[r_addr_li];

  always_ff @(posedge w_clk_i) begin
    if (w_v_i) begin
      mem[w_addr_li] <= w_data_i;
    end
  end
   end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_1r1w_synth)
// MBT 11/9/2014
//
// Synchronous 1-port ram.
// Only one read or one write may be done per cycle.
//
// NOTE: Users of BaseJump STL should not instantiate this module directly
// they should use bsg_mem_1rw_sync_mask_write_bit.
//

//`include "bsg_defines.sv"

module bsg_mem_1rw_sync_mask_write_bit_synth
  #(parameter `BSG_INV_PARAM(width_p)
    , parameter `BSG_INV_PARAM(els_p)
    , parameter latch_last_read_p=0
    , parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
   )
   (input   clk_i
    , input reset_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0] data_i
    , input [addr_width_lp-1:0] addr_i
    , input v_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0] w_mask_i
    , input w_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0]  data_o
    );

   wire unused = reset_i;

   if (width_p == 0 || els_p == 0)
    begin: z
      wire unused0 = &{clk_i, data_i, addr_i, v_i, w_mask_i, w_i};
      assign data_o = '0;
    end
   else
    begin: nz

   logic [addr_width_lp-1:0] addr_r;
   logic [width_p-1:0] mem [els_p-1:0];
   logic read_en;
   
   wire [addr_width_lp-1:0] addr_li = (els_p>1) ? addr_i:'0;
   
   assign read_en = v_i & ~w_i;

   always_ff @(posedge clk_i)
     if (read_en)
       addr_r <= addr_li;
     else
       addr_r <= 'X;

   logic [width_p-1:0] data_out;

   assign data_out = mem[addr_r];

   if (latch_last_read_p)
     begin: llr
      logic read_en_r; 

      bsg_dff #(
        .width_p(1)
      ) read_en_dff (
        .clk_i(clk_i)
        ,.data_i(read_en)
        ,.data_o(read_en_r)
      );

      bsg_dff_en_bypass #(
        .width_p(width_p)
      ) dff_bypass (
        .clk_i(clk_i)
        ,.en_i(read_en_r)
        ,.data_i(data_out)
        ,.data_o(data_o)
      );
     end
   else
     begin: no_llr
       assign data_o = data_out;
     end



// The Verilator and non-Verilator models are functionally equivalent. However, Verilator
//   cannot handle an array of non-blocking assignments in a for loop. It would be nice to 
//   see if these two models synthesize the same, because we can then reduce to the Verilator
//   model and avoid double maintenence. One could also add this feature to Verilator...
//   (Identified in Verilator 4.011)
`ifdef VERILATOR
   logic [width_p-1:0] data_n;

   for (genvar i = 0; i < width_p; i++)
     begin : rof1
       assign data_n[i] = w_mask_i[i] ? data_i[i] : mem[addr_li][i];
     end // rof1

   always_ff @(posedge clk_i)
     if (v_i & w_i)
       mem[addr_li] <= data_n;

`else
 
// this code does not map correctly with Xilinx Ultrascale FPGAs 
// in Vivado, substitute this file with hard/ultrascale_plus/bsg_mem/bsg_mem_1rw_sync_mask_write_bit.sv
      
`BSG_VIVADO_SYNTH_FAILS
      
   always_ff @(posedge clk_i)
     if (v_i & w_i)
       for (integer i = 0; i < width_p; i=i+1)
         if (w_mask_i[i])
           mem[addr_li][i] <= data_i[i];
`endif
   end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_1rw_sync_mask_write_bit_synth)
// NOTE: Users of BaseJump STL should not instantiate this module directly
// they should use bsg_mem_1r1w_sync_mask_write_byte.

//`include "bsg_defines.sv"

module bsg_mem_1rw_sync_mask_write_byte_synth
  #(parameter `BSG_INV_PARAM(els_p)
    , parameter addr_width_lp = `BSG_SAFE_CLOG2(els_p)
    , parameter latch_last_read_p=0

    , parameter `BSG_INV_PARAM(data_width_p )
    , parameter write_mask_width_lp = data_width_p>>3
  )
  ( input clk_i
   ,input reset_i

   ,input v_i
   ,input w_i

   ,input [addr_width_lp-1:0]       addr_i
   ,input [`BSG_SAFE_MINUS(data_width_p, 1):0]        data_i
    // for each bit set in the mask, a byte is written
   ,input [`BSG_SAFE_MINUS(write_mask_width_lp, 1):0] write_mask_i

   ,output [`BSG_SAFE_MINUS(data_width_p, 1):0] data_o
  );

  genvar i;

  if (data_width_p == 0 || els_p == 0)
   begin: z
     wire unused0 = &{clk_i, reset_i, v_i, w_i, addr_i, data_i, write_mask_i};
     assign data_o = '0;
   end
  else
   begin: nz

  for(i=0; i<write_mask_width_lp; i=i+1)
  begin: bk
    bsg_mem_1rw_sync #( .width_p      (8)
                        ,.els_p        (els_p)
                        ,.addr_width_lp(addr_width_lp)
                        ,.latch_last_read_p(latch_last_read_p)
			,.verbose_if_synth_p(0) // don't print out details of ram if breaks into synth srams
                      ) mem_1rw_sync
                      ( .clk_i  (clk_i)
                       ,.reset_i(reset_i)
                       ,.data_i (data_i[(i*8)+:8])
                       ,.addr_i (addr_i)
                       ,.v_i    (v_i & (w_i ? write_mask_i[i] : 1'b1))
                       ,.w_i    (w_i & write_mask_i[i])
                       ,.data_o (data_o[(i*8)+:8])
                      );
  end
   end

endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_1rw_sync_mask_write_byte_synth)
// MBT 11/9/2014
//
// Synchronous 1-port ram.
// Only one read or one write may be done per cycle.
//
// NOTE: Users of BaseJump STL should not instantiate this module directly
// they should use bsg_mem_1rw_sync.

//`include "bsg_defines.sv"

module bsg_mem_1rw_sync_synth
  #(parameter `BSG_INV_PARAM(width_p)
    , parameter `BSG_INV_PARAM(els_p)
    , parameter latch_last_read_p=0
    , parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
    , parameter verbose_p=1
   )
   (input   clk_i
	 	, input v_i
		, input reset_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0] data_i
    , input [addr_width_lp-1:0] addr_i
    , input w_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0]  data_o
    );

  wire unused = reset_i;

  if (width_p == 0 || els_p == 0)
   begin: z
     wire unused0 = &{clk_i, v_i, data_i, addr_i, w_i};
     assign data_o = '0;
   end
  else
   begin: nz

    logic [addr_width_lp-1:0] addr_r;
    logic [width_p-1:0]    mem [els_p-1:0];
    logic read_en;
    logic [width_p-1:0] data_out;

    wire [addr_width_lp-1:0] addr_li = (els_p>0) ? addr_i:'0;

    assign read_en = v_i & ~w_i;
    assign data_out = mem[addr_r];

    always_ff @ (posedge clk_i) 
      if (read_en)
        addr_r <= addr_li;
      else
        addr_r <= 'X;

    if (latch_last_read_p)
      begin: llr
        logic read_en_r; 

        bsg_dff #(
          .width_p(1)
        ) read_en_dff (
          .clk_i(clk_i)
          ,.data_i(read_en)
          ,.data_o(read_en_r)
        );

        bsg_dff_en_bypass #(
          .width_p(width_p)
        ) dff_bypass (
          .clk_i(clk_i)
          ,.en_i(read_en_r)
          ,.data_i(data_out)
          ,.data_o(data_o)
        );
      end
    else
      begin: no_llr
        assign data_o = data_out;
      end


    always_ff @(posedge clk_i)
      if (v_i & w_i) 
        mem[addr_li] <= data_i;
   end // non_zero_width
`ifndef BSG_HIDE_FROM_SYNTHESIS
   initial
     begin
        if (verbose_p)
	  $display("## %L: instantiating width_p=%d, els_p=%d (%m)",width_p,els_p);
     end
   

   always_ff @(negedge clk_i)
     if (v_i)
       assert ( (v_i !== 1'b1) || (reset_i === 'X) || (reset_i === 1'b1) || (addr_i < els_p) || (els_p <= 1))
         else $error("Invalid address %x to %m of size %x (reset_i = %b, v_i = %b, clk_i = %b)\n", addr_i, els_p, reset_i, v_i, clk_i);
`endif

endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_1rw_sync_synth)
// MBT 7/7/2016
//
// 2 read-port, 1 write-port ram
//
// reads are synchronous
//
// although we could merge this with normal bsg_mem_1r1w
// and select with a parameter, we do not do this because
// it's typically a very big change to the instantiating code
// to move to/from sync/async, and we want to reflect this.
//
// NOTE: Users of BaseJump STL should not instantiate this module directly
// they should use bsg_mem_2r1w_sync.

//`include "bsg_defines.sv"

module bsg_mem_2r1w_sync_synth #(parameter `BSG_INV_PARAM(width_p)
				 , parameter `BSG_INV_PARAM(els_p)
				 , parameter read_write_same_addr_p=0
				 , parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
				 )
   (input   clk_i
    , input reset_i

    , input                     w_v_i
    , input [addr_width_lp-1:0] w_addr_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0]       w_data_i

    // currently unused
    , input                      r0_v_i
    , input [addr_width_lp-1:0]  r0_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r0_data_o

    , input                      r1_v_i
    , input [addr_width_lp-1:0]  r1_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r1_data_o
    );

   wire                   unused = reset_i;

   if (width_p == 0)
    begin: z
      wire unused0 = &{clk_i, w_v_i, w_addr_i, w_data_i, r0_v_i, r0_addr_i, r1_v_i, r1_addr_i};
      assign r0_data_o = '0;
      assign r1_data_o = '0;
    end
   else
    begin: nz

   logic [width_p-1:0]    mem [els_p-1:0];

   // keep consistent with bsg_ip_cores/bsg_mem/bsg_mem_2r1w_sync.sv
   // keep consistent with bsg_ip_cores/hard/bsg_mem/bsg_mem_2r1w_sync.sv
   
   // this treats the ram as an array of registers for which the
   // read addr is latched on the clock, the write
   // is done on the clock edge, and actually multiplexing
   // of the registers for reading is done after the clock edge.

   // logically, this means that reads happen in time after
   // the writes, and "simultaneous" reads and writes to the
   // register file are allowed -- IF read_write_same_addr is set.

   // note that this behavior is generally incompatible with
   // hardened 1r1w rams, so it's better not to take advantage
   // of it if not necessary

   // we explicitly 'X out the read address if valid is not set
   // to avoid accidental use of data when the valid signal was not
   // asserted. without this, the output of the register file would
   // "auto-update" based on new writes to the ram, a spooky behavior
   // that would never correspond to that of a hardened ram.
   
   //the read logic, register the input
   logic [addr_width_lp-1:0]  r0_addr_r, r1_addr_r;

   always_ff @(posedge clk_i)
     if (r0_v_i)
       r0_addr_r <= r0_addr_i;
     else
       r0_addr_r <= 'X;

   always_ff @(posedge clk_i)
     if (r1_v_i)
       r1_addr_r <= r1_addr_i;
     else
       r1_addr_r <= 'X;

   assign r0_data_o = mem[ r0_addr_r ];
   assign r1_data_o = mem[ r1_addr_r ];

   //the write logic, the memory is treated as dff array
   always_ff @(posedge clk_i)
     if (w_v_i)
       mem[w_addr_i] <= w_data_i;

   end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_2r1w_sync_synth)
// MBT 4/1/2014
//
// 2 read-port, 1 write-port ram
//
// reads are asynchronous
//
// this file should not be directly instantiated by end programmers
// use bsg_mem_2r1w instead
//

//`include "bsg_defines.sv"

module bsg_mem_2r1w_synth #(parameter `BSG_INV_PARAM(width_p)
			    , parameter `BSG_INV_PARAM(els_p)
			    , parameter read_write_same_addr_p=0
			    , parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
			    )
   (input   w_clk_i
    , input w_reset_i

    , input                     w_v_i
    , input [addr_width_lp-1:0] w_addr_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0]       w_data_i

    , input                      r0_v_i
    , input [addr_width_lp-1:0]  r0_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r0_data_o

    , input                      r1_v_i
    , input [addr_width_lp-1:0]  r1_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r1_data_o

    );

   wire                   unused = w_reset_i;

   if (width_p == 0 || els_p == 0)
    begin: z
      wire unused0 = &{w_clk_i, w_v_i, w_addr_i, w_data_i, r0_v_i, r0_addr_i, r1_v_i, r1_addr_i};
      assign r0_data_o = '0;
      assign r1_data_o = '0;
    end
   else
    begin: nz

   logic [width_p-1:0]    mem [els_p-1:0];

   // this implementation ignores the r_v_i
   wire [addr_width_lp-1:0]  r0_addr_li = (els_p>1) ? r0_addr_i:'0;
   wire [addr_width_lp-1:0]  r1_addr_li = (els_p>1) ? r1_addr_i:'0;

   assign r1_data_o = mem[r1_addr_li];
   assign r0_data_o = mem[r0_addr_li];
   
   wire [addr_width_lp-1:0]  w_addr_li = (els_p>1) ? w_addr_i:'0;

   always_ff @(posedge w_clk_i)
     if (w_v_i)
       begin
          mem[w_addr_li] <= w_data_i;
       end
   end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_2r1w_synth)

//`include "bsg_defines.sv"

module bsg_mem_2rw_sync_mask_write_bit_synth #( parameter `BSG_INV_PARAM(width_p )
                         , parameter `BSG_INV_PARAM(els_p )
                         , parameter read_write_same_addr_p = 0
                         , parameter disable_collision_warning_p = 0
                         , parameter addr_width_lp = `BSG_SAFE_CLOG2(els_p)
                         , parameter harden_p = 1
                         )
  ( input                      clk_i
  , input                      reset_i

  , input [width_p-1:0]        a_data_i
  , input [width_p-1:0]        a_w_mask_i
  , input [addr_width_lp-1:0]  a_addr_i
  , input                      a_v_i
  , input                      a_w_i

  , input [width_p-1:0]        b_data_i
  , input [width_p-1:0]        b_w_mask_i
  , input [addr_width_lp-1:0]  b_addr_i
  , input                      b_v_i
  , input                      b_w_i

  , output logic [width_p-1:0] a_data_o
  , output logic [width_p-1:0] b_data_o
  );

   wire                   unused = reset_i;

   if (width_p == 0)
    begin: z
      wire unused0 = &{clk_i, a_data_i, a_w_mask_i, a_addr_i, a_v_i, a_w_i};
      wire unused1 = &{clk_i, b_data_i, b_w_mask_i, b_addr_i, b_v_i, b_w_i};
      assign a_data_o = '0;
      assign b_data_o = '0;
    end
   else
    begin: nz

   logic [width_p-1:0]    mem [els_p-1:0];

   // this treats the ram as an array of registers for which the
   // read addr is latched on the clock, the write
   // is done on the clock edge, and actually multiplexing
   // of the registers for reading is done after the clock edge.

   // logically, this means that reads happen in time after
   // the writes, and "simultaneous" reads and writes to the
   // register file are allowed -- IF read_write_same_addr is set.

   // note that this behavior is generally incompatible with
   // hardened 1r1w rams, so it's better not to take advantage
   // of it if not necessary

   // we explicitly 'X out the read address if valid is not set
   // to avoid accidental use of data when the valid signal was not
   // asserted. without this, the output of the register file would
   // "auto-update" based on new writes to the ram, a spooky behavior
   // that would never correspond to that of a hardened ram.

   logic [addr_width_lp-1:0] a_addr_r, b_addr_r;

   always_ff @(posedge clk_i)
     begin
        if (a_v_i)
            a_addr_r <= a_addr_i;
        else
            a_addr_r <= 'X;
          
        if (b_v_i)
            b_addr_r <= b_addr_i;
        else
            b_addr_r <= 'X;

`ifndef BSG_HIDE_FROM_SYNTHESIS
        // if addresses match and this is forbidden, then nuke the read address

        if (a_addr_i == b_addr_i && a_v_i && b_v_i && (a_w_i || b_w_i) && !read_write_same_addr_p)
          begin
             if (!disable_collision_warning_p)
               begin
                 $error("X'ing matched read addresses %x %x (%m)",a_addr_i, b_addr_i);
               end
             a_addr_r <= 'X;
             b_addr_r <= 'X;
          end
`endif

     end

   assign a_data_o = mem[a_addr_r];
   assign b_data_o = mem[b_addr_r];


   genvar                       i;
   for (i = 0; i < width_p; i=i+1)
     begin
	always_ff @(posedge clk_i)
      begin

	  if (a_v_i & a_w_i && a_w_mask_i[i])
            mem[a_addr_i][i] <= a_data_i[i];
	  if (b_v_i & b_w_i && b_w_mask_i[i])
            mem[b_addr_i][i] <= b_data_i[i];
      end
     end
  end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_2rw_sync_mask_write_bit_synth)

//`include "bsg_defines.sv"

module bsg_mem_2rw_sync_mask_write_byte_synth #( parameter `BSG_INV_PARAM(width_p )
                         , parameter `BSG_INV_PARAM(els_p )
                         , parameter read_write_same_addr_p=0
                         , parameter addr_width_lp = `BSG_SAFE_CLOG2(els_p)
                         , parameter harden_p = 1
                         , parameter disable_collision_warning_p=0     
                         , parameter write_mask_width_lp=(width_p>>3)              
                         )
  ( input                      clk_i
  , input                      reset_i

  , input [width_p-1:0]        a_data_i
  , input [write_mask_width_lp-1:0] a_w_mask_i
  , input [addr_width_lp-1:0]  a_addr_i
  , input                      a_v_i
  , input                      a_w_i

  , input [width_p-1:0]        b_data_i
  , input [write_mask_width_lp-1:0] b_w_mask_i
  , input [addr_width_lp-1:0]  b_addr_i
  , input                      b_v_i
  , input                      b_w_i

  , output logic [width_p-1:0] a_data_o
  , output logic [width_p-1:0] b_data_o
  );

   wire                   unused = reset_i;

   if (width_p == 0)
    begin: z
      wire unused0 = &{clk_i, a_data_i, a_w_mask_i, a_addr_i, a_v_i, a_w_i};
      wire unused1 = &{clk_i, b_data_i, b_w_mask_i, b_addr_i, b_v_i, b_w_i};
      assign a_data_o = '0;
      assign b_data_o = '0;
    end
   else
    begin: nz

  genvar i;
  for(i=0; i<write_mask_width_lp; i=i+1)
  begin: bk
    bsg_mem_2rw_sync #( .width_p      (8)
                        ,.els_p        (els_p)
                        ,.addr_width_lp(addr_width_lp)
                        ,.disable_collision_warning_p(disable_collision_warning_p)
                        ,.harden_p(harden_p)
                      ) mem_2rw_sync
                      ( .clk_i  (clk_i)
                       ,.reset_i(reset_i)
                       ,.a_data_i (a_data_i[(i*8)+:8])
                       ,.a_addr_i (a_addr_i)
                       ,.a_v_i    (a_v_i & (a_w_i ? a_w_mask_i[i] : 1'b1))
                       ,.a_w_i    (a_w_i & a_w_mask_i[i])
                       ,.a_data_o (a_data_o[(i*8)+:8])
                       ,.b_data_i (b_data_i[(i*8)+:8])
                       ,.b_addr_i (b_addr_i)
                       ,.b_v_i    (b_v_i & (b_w_i ? b_w_mask_i[i] : 1'b1))
                       ,.b_w_i    (b_w_i & b_w_mask_i[i])
                       ,.b_data_o (b_data_o[(i*8)+:8])
                      );
  end
    end

endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_2rw_sync_mask_write_byte_synth)


//`include "bsg_defines.sv"

module bsg_mem_2rw_sync_synth #( parameter `BSG_INV_PARAM(width_p )
                         , parameter `BSG_INV_PARAM(els_p )
                         , parameter read_write_same_addr_p=0
                         , parameter addr_width_lp = `BSG_SAFE_CLOG2(els_p)
                         , parameter harden_p = 1
                         , parameter disable_collision_warning_p=0                   
                         )
  ( input                      clk_i
  , input                      reset_i

  , input [width_p-1:0]        a_data_i
  , input [addr_width_lp-1:0]  a_addr_i
  , input                      a_v_i
  , input                      a_w_i

  , input [width_p-1:0]        b_data_i
  , input [addr_width_lp-1:0]  b_addr_i
  , input                      b_v_i
  , input                      b_w_i

  , output logic [width_p-1:0] a_data_o
  , output logic [width_p-1:0] b_data_o
  );

   wire                   unused = reset_i;

   if (width_p == 0)
    begin: z
      wire unused0 = &{clk_i, a_data_i, a_addr_i, a_v_i, a_w_i};
      wire unused1 = &{clk_i, b_data_i, b_addr_i, b_v_i, b_w_i};
      assign a_data_o = '0;
      assign b_data_o = '0;
    end
   else
    begin: nz

   logic [width_p-1:0]    mem [els_p-1:0];

   // this treats the ram as an array of registers for which the
   // read addr is latched on the clock, the write
   // is done on the clock edge, and actually multiplexing
   // of the registers for reading is done after the clock edge.

   // logically, this means that reads happen in time after
   // the writes, and "simultaneous" reads and writes to the
   // register file are allowed -- IF read_write_same_addr is set.

   // note that this behavior is generally incompatible with
   // hardened 1r1w rams, so it's better not to take advantage
   // of it if not necessary

   // we explicitly 'X out the read address if valid is not set
   // to avoid accidental use of data when the valid signal was not
   // asserted. without this, the output of the register file would
   // "auto-update" based on new writes to the ram, a spooky behavior
   // that would never correspond to that of a hardened ram.

   logic [addr_width_lp-1:0] a_addr_r, b_addr_r;

   always_ff @(posedge clk_i)
     begin
        if (a_v_i)
            a_addr_r <= a_addr_i;
        else
            a_addr_r <= 'X;
          
        if (b_v_i)
            b_addr_r <= b_addr_i;
        else
            b_addr_r <= 'X;

`ifndef BSG_HIDE_FROM_SYNTHESIS
        // if addresses match and this is forbidden, then nuke the read address

        if (a_addr_i == b_addr_i && a_v_i && b_v_i && (a_w_i || b_w_i) && !read_write_same_addr_p)
          begin
             if (!disable_collision_warning_p)
               begin
                 $error("X'ing matched read address %x (%m)",a_addr_i);
               end
             a_addr_r <= 'X;
             b_addr_r <= 'X;
          end
`endif

     end

   assign a_data_o = mem[a_addr_r];
   assign b_data_o = mem[b_addr_r];

	always_ff @(posedge clk_i)
    begin
	  if (a_v_i & a_w_i)
            mem[a_addr_i] <= a_data_i;
	  if (b_v_i & b_w_i)
            mem[b_addr_i] <= b_data_i;
    end
  end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_2rw_sync_synth)

// MBT 7/7/2016
// DWP 11/27/2019
//
// 3 read-port, 1 write-port ram
//
// reads are synchronous
//
// although we could merge this with normal bsg_mem_1r1w
// and select with a parameter, we do not do this because
// it's typically a very big change to the instantiating code
// to move to/from sync/async, and we want to reflect this.
//
// NOTE: Users of BaseJump STL should not instantiate this module directly
// they should use bsg_mem_3r1w_sync.

//`include "bsg_defines.sv"

module bsg_mem_3r1w_sync_synth #(parameter `BSG_INV_PARAM(width_p)
				 , parameter `BSG_INV_PARAM(els_p)
				 , parameter read_write_same_addr_p=0
				 , parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
				 )
   (input   clk_i
    , input reset_i

    , input                     w_v_i
    , input [addr_width_lp-1:0] w_addr_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0]       w_data_i

    // currently unused
    , input                      r0_v_i
    , input [addr_width_lp-1:0]  r0_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r0_data_o

    , input                      r1_v_i
    , input [addr_width_lp-1:0]  r1_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r1_data_o

    , input                      r2_v_i
    , input [addr_width_lp-1:0]  r2_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r2_data_o
    );

   wire                   unused = reset_i;

   if (width_p == 0)
    begin: z
      wire unused0 = &{clk_i, w_v_i, w_addr_i, w_data_i, r0_v_i, r0_addr_i, r1_v_i, r1_addr_i, r2_v_i, r2_addr_i};
      assign r0_data_o = '0;
      assign r1_data_o = '0;
      assign r2_data_o = '0;
    end
   else
    begin: nz

   logic [width_p-1:0]    mem [els_p-1:0];

   // keep consistent with bsg_ip_cores/bsg_mem/bsg_mem_3r1w_sync.sv
   // keep consistent with bsg_ip_cores/hard/bsg_mem/bsg_mem_3r1w_sync.sv

   // this treats the ram as an array of registers for which the
   // read addr is latched on the clock, the write
   // is done on the clock edge, and actually multiplexing
   // of the registers for reading is done after the clock edge.

   // logically, this means that reads happen in time after
   // the writes, and "simultaneous" reads and writes to the
   // register file are allowed -- IF read_write_same_addr is set.

   // note that this behavior is generally incompatible with
   // hardened 1r1w rams, so it's better not to take advantage
   // of it if not necessary

   // we explicitly 'X out the read address if valid is not set
   // to avoid accidental use of data when the valid signal was not
   // asserted. without this, the output of the register file would
   // "auto-update" based on new writes to the ram, a spooky behavior
   // that would never correspond to that of a hardened ram.

   //the read logic, register the input
   logic [addr_width_lp-1:0]  r0_addr_r, r1_addr_r, r2_addr_r;

   always_ff @(posedge clk_i)
     if (r0_v_i)
       r0_addr_r <= r0_addr_i;
     else
       r0_addr_r <= 'X;

   always_ff @(posedge clk_i)
     if (r1_v_i)
       r1_addr_r <= r1_addr_i;
     else
       r1_addr_r <= 'X;

   always_ff @(posedge clk_i)
     if (r2_v_i)
       r2_addr_r <= r2_addr_i;
     else
       r2_addr_r <= 'X;

   assign r0_data_o = mem[ r0_addr_r ];
   assign r1_data_o = mem[ r1_addr_r ];
   assign r2_data_o = mem[ r2_addr_r ];

   //the write logic, the memory is treated as dff array
   always_ff @(posedge clk_i)
     if (w_v_i)
       mem[w_addr_i] <= w_data_i;

    end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_3r1w_sync_synth)
// MBT 4/1/2014
// DWP 11/27/2019
//
// 3 read-port, 1 write-port ram
//
// reads are asynchronous
//
// this file should not be directly instantiated by end programmers
// use bsg_mem_3r1w instead
//

//`include "bsg_defines.sv"

module bsg_mem_3r1w_synth #(parameter `BSG_INV_PARAM(width_p)
			    , parameter `BSG_INV_PARAM(els_p)
			    , parameter read_write_same_addr_p=0
			    , parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
			    )
   (input   w_clk_i
    , input w_reset_i

    , input                     w_v_i
    , input [addr_width_lp-1:0] w_addr_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0]       w_data_i

    , input                      r0_v_i
    , input [addr_width_lp-1:0]  r0_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r0_data_o

    , input                      r1_v_i
    , input [addr_width_lp-1:0]  r1_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r1_data_o

    , input                      r2_v_i
    , input [addr_width_lp-1:0]  r2_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r2_data_o
    );

   wire                   unused = w_reset_i;

   if (width_p == 0)
    begin: z
      wire unused0 = &{w_clk_i, w_v_i, w_addr_i, w_data_i, r0_v_i, r0_addr_i, r1_v_i, r1_addr_i, r2_v_i, r2_addr_i};
      assign r0_data_o = '0;
      assign r1_data_o = '0;
      assign r2_data_o = '0;
    end
   else
    begin: nz

   logic [width_p-1:0]    mem [els_p-1:0];

   // this implementation ignores the r_v_i
   assign r2_data_o = mem[r2_addr_i];
   assign r1_data_o = mem[r1_addr_i];
   assign r0_data_o = mem[r0_addr_i];

   wire                   unused = w_reset_i;

   always_ff @(posedge w_clk_i)
     if (w_v_i)
       begin
          mem[w_addr_i] <= w_data_i;
       end
    end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_3r1w_synth)


module bsg_dff_reset_en_width_p2_reset_val_p0_harden_p0
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [1:0] data_i;
  output [1:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [1:0] data_o;
  wire N0,N1,N2;
  reg data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_en_bypass_width_p2
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [1:0] data_i;
  output [1:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [1:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_reset_en_width_p2_reset_val_p0_harden_p0
  dff
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(en_i),
    .data_i(data_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_dff_reset_en_width_p1_reset_val_p0_harden_p0
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [0:0] data_o;
  wire N0,N1,N2;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_en_bypass_width_p1
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [0:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_reset_en_width_p1_reset_val_p0_harden_p0
  dff
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(en_i),
    .data_i(data_i[0]),
    .data_o(data_r[0])
  );

  assign data_o[0] = (N0)? data_i[0] : 
                     (N1)? data_r[0] : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_counter_clear_up_max_val_p64_init_val_p0
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [6:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire [6:0] count_o;
  wire N0,N1,N4,N5,N6,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N2,N3,N7,N30,N20;
  reg count_o_6_sv2v_reg,count_o_5_sv2v_reg,count_o_4_sv2v_reg,count_o_3_sv2v_reg,
  count_o_2_sv2v_reg,count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[6] = count_o_6_sv2v_reg;
  assign count_o[5] = count_o_5_sv2v_reg;
  assign count_o[4] = count_o_4_sv2v_reg;
  assign count_o[3] = count_o_3_sv2v_reg;
  assign count_o[2] = count_o_2_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign N20 = reset_i | clear_i;
  assign { N12, N11, N10, N9, N8, N6, N5 } = count_o + 1'b1;
  assign N13 = (N0)? 1'b1 : 
               (N7)? 1'b1 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = clear_i;
  assign N15 = (N1)? 1'b1 : 
               (N30)? 1'b0 : 1'b0;
  assign N1 = up_i;
  assign N14 = (N0)? up_i : 
               (N7)? N5 : 1'b0;
  assign N4 = N19;
  assign N16 = ~reset_i;
  assign N17 = ~clear_i;
  assign N18 = N16 & N17;
  assign N19 = up_i & N18;
  assign N2 = up_i | clear_i;
  assign N3 = ~N2;
  assign N7 = up_i & N17;
  assign N30 = ~up_i;

  always @(posedge clk_i) begin
    if(N20) begin
      count_o_6_sv2v_reg <= 1'b0;
      count_o_5_sv2v_reg <= 1'b0;
      count_o_4_sv2v_reg <= 1'b0;
      count_o_3_sv2v_reg <= 1'b0;
      count_o_2_sv2v_reg <= 1'b0;
      count_o_1_sv2v_reg <= 1'b0;
    end else if(N15) begin
      count_o_6_sv2v_reg <= N12;
      count_o_5_sv2v_reg <= N11;
      count_o_4_sv2v_reg <= N10;
      count_o_3_sv2v_reg <= N9;
      count_o_2_sv2v_reg <= N8;
      count_o_1_sv2v_reg <= N6;
    end 
    if(reset_i) begin
      count_o_0_sv2v_reg <= 1'b0;
    end else if(N13) begin
      count_o_0_sv2v_reg <= N14;
    end 
  end


endmodule



module bsg_mem_1r1w_sync_width_p50_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [5:0] w_addr_i;
  input [49:0] w_data_i;
  input [5:0] r_addr_i;
  output [49:0] r_data_o;
  input clk_i;
  input reset_i;
  input w_v_i;
  input r_v_i;
  wire [49:0] r_data_o;

  bsg_mem_1r1w_sync_synth
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_dff_reset_set_clear_width_p1
(
  clk_i,
  reset_i,
  set_i,
  clear_i,
  data_o
);

  input [0:0] set_i;
  input [0:0] clear_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  wire [0:0] data_o;
  wire N0,N1,N2;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N0 = N2 | set_i[0];
  assign N2 = data_o[0] & N1;
  assign N1 = ~clear_i[0];

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_0_sv2v_reg <= N0;
    end 
  end


endmodule



module bsg_dff_reset_en_0000000f
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [14:0] data_i;
  output [14:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [14:0] data_o;
  wire N0,N1,N2;
  reg data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bp_fe_btb_00
(
  clk_i,
  reset_i,
  init_done_o,
  r_addr_i,
  r_v_i,
  r_tag_o,
  r_idx_o,
  r_tgt_o,
  r_tgt_v_o,
  r_tgt_jmp_o,
  w_v_i,
  w_force_i,
  w_clr_i,
  w_jmp_i,
  w_tag_i,
  w_idx_i,
  w_tgt_i,
  w_yumi_o
);

  input [38:0] r_addr_i;
  output [8:0] r_tag_o;
  output [5:0] r_idx_o;
  output [38:0] r_tgt_o;
  input [8:0] w_tag_i;
  input [5:0] w_idx_i;
  input [38:0] w_tgt_i;
  input clk_i;
  input reset_i;
  input r_v_i;
  input w_v_i;
  input w_force_i;
  input w_clr_i;
  input w_jmp_i;
  output init_done_o;
  output r_tgt_v_o;
  output r_tgt_jmp_o;
  output w_yumi_o;
  wire [8:0] r_tag_o;
  wire [5:0] r_idx_o,w_addr_li;
  wire [38:0] r_tgt_o;
  wire init_done_o,r_tgt_v_o,r_tgt_jmp_o,w_yumi_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,
  N11,N12,rw_same_addr,suppress_read,suppress_write,w_v_li,N13,N14,N15,N16,r_v_li,
  N17,r_data_lo_v_,r_data_lo_jmp_,r_data_lo_tag__8_,r_data_lo_tag__7_,
  r_data_lo_tag__6_,r_data_lo_tag__5_,r_data_lo_tag__4_,r_data_lo_tag__3_,r_data_lo_tag__2_,
  r_data_lo_tag__1_,r_data_lo_tag__0_,r_v_r,N18,N19,N20,N22,N23,N24,N25,N26,N27,N28,
  N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45;
  wire [1:0] state_r,state_n;
  wire [6:0] init_cnt;
  wire [49:0] w_data_li;
  wire [0:0] r_idx_li;
  reg state_r_1_sv2v_reg,state_r_0_sv2v_reg;
  assign state_r[1] = state_r_1_sv2v_reg;
  assign state_r[0] = state_r_0_sv2v_reg;

  bsg_counter_clear_up_max_val_p64_init_val_p0
  init_counter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(1'b0),
    .up_i(N24),
    .count_o(init_cnt)
  );

  assign N6 = state_r[1] | N22;
  assign N8 = N19 | state_r[0];
  assign N10 = state_r[1] & state_r[0];
  assign N11 = N19 & N22;
  assign N17 = { r_addr_i[7:3], r_idx_li[0:0] } == w_idx_i;

  bsg_mem_1r1w_sync_width_p50_els_p64_latch_last_read_p1
  btb_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(w_v_li),
    .w_addr_i(w_addr_li),
    .w_data_i(w_data_li),
    .r_v_i(r_v_li),
    .r_addr_i({ r_addr_i[7:3], r_idx_li[0:0] }),
    .r_data_o({ r_data_lo_v_, r_data_lo_jmp_, r_data_lo_tag__8_, r_data_lo_tag__7_, r_data_lo_tag__6_, r_data_lo_tag__5_, r_data_lo_tag__4_, r_data_lo_tag__3_, r_data_lo_tag__2_, r_data_lo_tag__1_, r_data_lo_tag__0_, r_tgt_o })
  );


  bsg_dff_reset_set_clear_width_p1
  r_v_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .set_i(r_v_li),
    .clear_i(r_v_i),
    .data_o(r_v_r)
  );


  bsg_dff_reset_en_0000000f
  tag_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(r_v_i),
    .data_i({ r_addr_i[7:3], r_idx_li[0:0], r_addr_i[16:8] }),
    .data_o({ r_idx_o, r_tag_o })
  );

  assign N18 = { r_data_lo_tag__8_, r_data_lo_tag__7_, r_data_lo_tag__6_, r_data_lo_tag__5_, r_data_lo_tag__4_, r_data_lo_tag__3_, r_data_lo_tag__2_, r_data_lo_tag__1_, r_data_lo_tag__0_ } == r_tag_o;
  assign N19 = ~state_r[1];
  assign N20 = state_r[0] | N19;
  assign init_done_o = ~N20;
  assign N22 = ~state_r[0];
  assign N23 = N22 | state_r[1];
  assign N24 = ~N23;
  assign N25 = ~init_cnt[5];
  assign N26 = ~init_cnt[4];
  assign N27 = ~init_cnt[3];
  assign N28 = ~init_cnt[2];
  assign N29 = ~init_cnt[1];
  assign N30 = ~init_cnt[0];
  assign N31 = N25 | init_cnt[6];
  assign N32 = N26 | N31;
  assign N33 = N27 | N32;
  assign N34 = N28 | N33;
  assign N35 = N29 | N34;
  assign N36 = N30 | N35;
  assign N37 = ~N36;
  assign state_n = (N0)? { N37, N36 } : 
                   (N1)? { 1'b1, 1'b0 } : 
                   (N2)? { 1'b0, 1'b1 } : 1'b0;
  assign N0 = N7;
  assign N1 = N9;
  assign N2 = N12;
  assign w_addr_li = (N3)? init_cnt[5:0] : 
                     (N4)? w_idx_i : 1'b0;
  assign N3 = N14;
  assign N4 = N13;
  assign w_data_li[49] = ~N15;
  assign w_data_li[48:0] = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N16)? { w_jmp_i, w_tag_i, w_tgt_i } : 1'b0;
  assign N5 = N15;
  assign N7 = ~N6;
  assign N9 = ~N8;
  assign N12 = N10 | N11;
  assign suppress_read = rw_same_addr & w_force_i;
  assign suppress_write = rw_same_addr & N38;
  assign N38 = ~w_force_i;
  assign w_v_li = N24 | N40;
  assign N40 = w_v_i & N39;
  assign N39 = ~suppress_write;
  assign N13 = ~N24;
  assign N14 = N24;
  assign N15 = N24 | N41;
  assign N41 = w_v_i & w_clr_i;
  assign N16 = ~N15;
  assign r_v_li = r_v_i & N42;
  assign N42 = ~suppress_read;
  assign r_idx_li[0] = r_addr_i[2] ^ r_addr_i[1];
  assign rw_same_addr = N43 & N17;
  assign N43 = r_v_i & w_v_i;
  assign w_yumi_o = init_done_o & w_v_li;
  assign r_tgt_v_o = N44 & N18;
  assign N44 = r_v_r & r_data_lo_v_;
  assign r_tgt_jmp_o = N45 & r_data_lo_jmp_;
  assign N45 = r_v_r & r_data_lo_v_;

  always @(posedge clk_i) begin
    if(reset_i) begin
      state_r_1_sv2v_reg <= 1'b0;
      state_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      state_r_1_sv2v_reg <= state_n[1];
      state_r_0_sv2v_reg <= state_n[0];
    end 
  end


endmodule



module bsg_counter_clear_up_max_val_p512_init_val_p0
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [9:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire [9:0] count_o;
  wire N0,N1,N4,N5,N6,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N2,N3,
  N7,N30,N23;
  reg count_o_9_sv2v_reg,count_o_8_sv2v_reg,count_o_7_sv2v_reg,count_o_6_sv2v_reg,
  count_o_5_sv2v_reg,count_o_4_sv2v_reg,count_o_3_sv2v_reg,count_o_2_sv2v_reg,
  count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[9] = count_o_9_sv2v_reg;
  assign count_o[8] = count_o_8_sv2v_reg;
  assign count_o[7] = count_o_7_sv2v_reg;
  assign count_o[6] = count_o_6_sv2v_reg;
  assign count_o[5] = count_o_5_sv2v_reg;
  assign count_o[4] = count_o_4_sv2v_reg;
  assign count_o[3] = count_o_3_sv2v_reg;
  assign count_o[2] = count_o_2_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign N23 = reset_i | clear_i;
  assign { N15, N14, N13, N12, N11, N10, N9, N8, N6, N5 } = count_o + 1'b1;
  assign N16 = (N0)? 1'b1 : 
               (N7)? 1'b1 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = clear_i;
  assign N18 = (N1)? 1'b1 : 
               (N30)? 1'b0 : 1'b0;
  assign N1 = up_i;
  assign N17 = (N0)? up_i : 
               (N7)? N5 : 1'b0;
  assign N4 = N22;
  assign N19 = ~reset_i;
  assign N20 = ~clear_i;
  assign N21 = N19 & N20;
  assign N22 = up_i & N21;
  assign N2 = up_i | clear_i;
  assign N3 = ~N2;
  assign N7 = up_i & N20;
  assign N30 = ~up_i;

  always @(posedge clk_i) begin
    if(N23) begin
      count_o_9_sv2v_reg <= 1'b0;
      count_o_8_sv2v_reg <= 1'b0;
      count_o_7_sv2v_reg <= 1'b0;
      count_o_6_sv2v_reg <= 1'b0;
      count_o_5_sv2v_reg <= 1'b0;
      count_o_4_sv2v_reg <= 1'b0;
      count_o_3_sv2v_reg <= 1'b0;
      count_o_2_sv2v_reg <= 1'b0;
      count_o_1_sv2v_reg <= 1'b0;
    end else if(N18) begin
      count_o_9_sv2v_reg <= N15;
      count_o_8_sv2v_reg <= N14;
      count_o_7_sv2v_reg <= N13;
      count_o_6_sv2v_reg <= N12;
      count_o_5_sv2v_reg <= N11;
      count_o_4_sv2v_reg <= N10;
      count_o_3_sv2v_reg <= N9;
      count_o_2_sv2v_reg <= N8;
      count_o_1_sv2v_reg <= N6;
    end 
    if(reset_i) begin
      count_o_0_sv2v_reg <= 1'b0;
    end else if(N16) begin
      count_o_0_sv2v_reg <= N17;
    end 
  end


endmodule



module bsg_mem_1r1w_sync_00000008_512_1
(
  clk_i,
  reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [8:0] w_addr_i;
  input [7:0] w_data_i;
  input [8:0] r_addr_i;
  output [7:0] r_data_o;
  input clk_i;
  input reset_i;
  input w_v_i;
  input r_v_i;
  wire [7:0] r_data_o;

  bsg_mem_1r1w_sync_synth
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_dff_en_00000009
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [8:0] data_i;
  output [8:0] data_o;
  input clk_i;
  input en_i;
  wire [8:0] data_o;
  reg data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,
  data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bp_fe_bht_00
(
  clk_i,
  reset_i,
  init_done_o,
  w_v_i,
  w_force_i,
  w_idx_i,
  w_offset_i,
  w_ghist_i,
  w_val_i,
  w_correct_i,
  w_yumi_o,
  r_v_i,
  r_addr_i,
  r_ghist_i,
  r_val_o,
  r_pred_o,
  r_idx_o,
  r_offset_o
);

  input [6:0] w_idx_i;
  input [1:0] w_offset_i;
  input [1:0] w_ghist_i;
  input [7:0] w_val_i;
  input [38:0] r_addr_i;
  input [1:0] r_ghist_i;
  output [7:0] r_val_o;
  output [6:0] r_idx_o;
  output [1:0] r_offset_o;
  input clk_i;
  input reset_i;
  input w_v_i;
  input w_force_i;
  input w_correct_i;
  input r_v_i;
  output init_done_o;
  output w_yumi_o;
  output r_pred_o;
  wire [7:0] r_val_o,w_data_li;
  wire [6:0] r_idx_o;
  wire [1:0] r_offset_o,state_r,state_n;
  wire init_done_o,w_yumi_o,r_pred_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,
  rw_same_addr,suppress_read,suppress_write,w_v_li,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,r_v_li,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97;
  wire [9:0] init_cnt;
  wire [8:0] w_addr_li;
  wire [3:0] w_mask_li;
  wire [0:0] r_idx_li;
  wire [2:0] pred_bit_lo;
  reg state_r_1_sv2v_reg,state_r_0_sv2v_reg;
  assign state_r[1] = state_r_1_sv2v_reg;
  assign state_r[0] = state_r_0_sv2v_reg;

  bsg_counter_clear_up_max_val_p512_init_val_p0
  init_counter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(1'b0),
    .up_i(N88),
    .count_o(init_cnt)
  );

  assign N5 = state_r[1] | N86;
  assign N7 = N64 | state_r[0];
  assign N9 = state_r[1] & state_r[0];
  assign N10 = N64 & N86;
  assign { N17, N16, N15, N14 } = { 1'b0, 1'b0, 1'b0, 1'b1 } << w_offset_i;
  assign N48 = { r_ghist_i, r_addr_i[8:3], r_idx_li[0:0] } == w_addr_li;

  bsg_mem_1r1w_sync_00000008_512_1
  bht_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(w_v_li),
    .w_addr_i(w_addr_li),
    .w_data_i(w_data_li),
    .r_v_i(r_v_li),
    .r_addr_i({ r_ghist_i, r_addr_i[8:3], r_idx_li[0:0] }),
    .r_data_o(r_val_o)
  );


  bsg_dff_en_00000009
  pred_idx_reg
  (
    .clk_i(clk_i),
    .data_i({ r_addr_i[10:3], r_idx_li[0:0] }),
    .en_i(r_v_i),
    .data_o({ r_offset_o, r_idx_o })
  );

  assign r_pred_o = (N56)? r_val_o[0] : 
                    (N58)? r_val_o[1] : 
                    (N60)? r_val_o[2] : 
                    (N62)? r_val_o[3] : 
                    (N57)? r_val_o[4] : 
                    (N59)? r_val_o[5] : 
                    (N61)? r_val_o[6] : 
                    (N63)? r_val_o[7] : 1'b0;
  assign N64 = ~state_r[1];
  assign N65 = state_r[0] | N64;
  assign init_done_o = ~N65;
  assign N67 = ~init_cnt[8];
  assign N68 = ~init_cnt[7];
  assign N69 = ~init_cnt[6];
  assign N70 = ~init_cnt[5];
  assign N71 = ~init_cnt[4];
  assign N72 = ~init_cnt[3];
  assign N73 = ~init_cnt[2];
  assign N74 = ~init_cnt[1];
  assign N75 = ~init_cnt[0];
  assign N76 = N67 | init_cnt[9];
  assign N77 = N68 | N76;
  assign N78 = N69 | N77;
  assign N79 = N70 | N78;
  assign N80 = N71 | N79;
  assign N81 = N72 | N80;
  assign N82 = N73 | N81;
  assign N83 = N74 | N82;
  assign N84 = N75 | N83;
  assign N85 = ~N84;
  assign N86 = ~state_r[0];
  assign N87 = N86 | state_r[1];
  assign N88 = ~N87;
  assign pred_bit_lo = { r_offset_o, 1'b0 } + 1'b1;
  assign state_n = (N0)? { N85, N84 } : 
                   (N1)? { 1'b1, 1'b0 } : 
                   (N2)? { 1'b0, 1'b1 } : 1'b0;
  assign N0 = N6;
  assign N1 = N8;
  assign N2 = N11;
  assign w_addr_li = (N3)? init_cnt[8:0] : 
                     (N4)? { w_ghist_i, w_idx_i } : 1'b0;
  assign N3 = N13;
  assign N4 = N12;
  assign w_mask_li = (N3)? { 1'b1, 1'b1, 1'b1, 1'b1 } : 
                     (N4)? { N17, N16, N15, N14 } : 1'b0;
  assign w_data_li[0] = (N3)? 1'b1 : 
                        (N22)? N20 : 
                        (N19)? w_val_i[0] : 1'b0;
  assign w_data_li[1] = (N3)? 1'b0 : 
                        (N26)? N25 : 
                        (N24)? w_val_i[1] : 1'b0;
  assign w_data_li[2] = (N3)? 1'b1 : 
                        (N29)? N20 : 
                        (N28)? w_val_i[2] : 1'b0;
  assign w_data_li[3] = (N3)? 1'b0 : 
                        (N33)? N32 : 
                        (N31)? w_val_i[3] : 1'b0;
  assign w_data_li[4] = (N3)? 1'b1 : 
                        (N36)? N20 : 
                        (N35)? w_val_i[4] : 1'b0;
  assign w_data_li[5] = (N3)? 1'b0 : 
                        (N40)? N39 : 
                        (N38)? w_val_i[5] : 1'b0;
  assign w_data_li[6] = (N3)? 1'b1 : 
                        (N43)? N20 : 
                        (N42)? w_val_i[6] : 1'b0;
  assign w_data_li[7] = (N3)? 1'b0 : 
                        (N47)? N46 : 
                        (N45)? w_val_i[7] : 1'b0;
  assign N6 = ~N5;
  assign N8 = ~N7;
  assign N11 = N9 | N10;
  assign suppress_read = rw_same_addr & w_force_i;
  assign suppress_write = rw_same_addr & N89;
  assign N89 = ~w_force_i;
  assign w_v_li = N88 | N91;
  assign N91 = w_v_i & N90;
  assign N90 = ~suppress_write;
  assign N12 = ~N88;
  assign N13 = N88;
  assign N18 = w_mask_li[0] | N13;
  assign N19 = ~N18;
  assign N20 = ~w_correct_i;
  assign N21 = ~N13;
  assign N22 = w_mask_li[0] & N21;
  assign N23 = w_mask_li[0] | N13;
  assign N24 = ~N23;
  assign N25 = w_val_i[1] ^ N92;
  assign N92 = N20 & w_val_i[0];
  assign N26 = w_mask_li[0] & N21;
  assign N27 = w_mask_li[1] | N13;
  assign N28 = ~N27;
  assign N29 = w_mask_li[1] & N21;
  assign N30 = w_mask_li[1] | N13;
  assign N31 = ~N30;
  assign N32 = w_val_i[3] ^ N93;
  assign N93 = N20 & w_val_i[2];
  assign N33 = w_mask_li[1] & N21;
  assign N34 = w_mask_li[2] | N13;
  assign N35 = ~N34;
  assign N36 = w_mask_li[2] & N21;
  assign N37 = w_mask_li[2] | N13;
  assign N38 = ~N37;
  assign N39 = w_val_i[5] ^ N94;
  assign N94 = N20 & w_val_i[4];
  assign N40 = w_mask_li[2] & N21;
  assign N41 = w_mask_li[3] | N13;
  assign N42 = ~N41;
  assign N43 = w_mask_li[3] & N21;
  assign N44 = w_mask_li[3] | N13;
  assign N45 = ~N44;
  assign N46 = w_val_i[7] ^ N95;
  assign N95 = N20 & w_val_i[6];
  assign N47 = w_mask_li[3] & N21;
  assign r_v_li = r_v_i & N96;
  assign N96 = ~suppress_read;
  assign r_idx_li[0] = r_addr_i[2] ^ r_addr_i[1];
  assign rw_same_addr = N97 & N48;
  assign N97 = r_v_i & w_v_i;
  assign w_yumi_o = init_done_o & w_v_li;
  assign N49 = ~pred_bit_lo[0];
  assign N50 = ~pred_bit_lo[1];
  assign N51 = N49 & N50;
  assign N52 = N49 & pred_bit_lo[1];
  assign N53 = pred_bit_lo[0] & N50;
  assign N54 = pred_bit_lo[0] & pred_bit_lo[1];
  assign N55 = ~pred_bit_lo[2];
  assign N56 = N51 & N55;
  assign N57 = N51 & pred_bit_lo[2];
  assign N58 = N53 & N55;
  assign N59 = N53 & pred_bit_lo[2];
  assign N60 = N52 & N55;
  assign N61 = N52 & pred_bit_lo[2];
  assign N62 = N54 & N55;
  assign N63 = N54 & pred_bit_lo[2];

  always @(posedge clk_i) begin
    if(reset_i) begin
      state_r_1_sv2v_reg <= 1'b0;
      state_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      state_r_1_sv2v_reg <= state_n[1];
      state_r_0_sv2v_reg <= state_n[0];
    end 
  end


endmodule



module bsg_dff_reset_en_0000005a
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [89:0] data_i;
  output [89:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [89:0] data_o;
  wire N0,N1,N2;
  reg data_o_89_sv2v_reg,data_o_88_sv2v_reg,data_o_87_sv2v_reg,data_o_86_sv2v_reg,
  data_o_85_sv2v_reg,data_o_84_sv2v_reg,data_o_83_sv2v_reg,data_o_82_sv2v_reg,
  data_o_81_sv2v_reg,data_o_80_sv2v_reg,data_o_79_sv2v_reg,data_o_78_sv2v_reg,
  data_o_77_sv2v_reg,data_o_76_sv2v_reg,data_o_75_sv2v_reg,data_o_74_sv2v_reg,
  data_o_73_sv2v_reg,data_o_72_sv2v_reg,data_o_71_sv2v_reg,data_o_70_sv2v_reg,data_o_69_sv2v_reg,
  data_o_68_sv2v_reg,data_o_67_sv2v_reg,data_o_66_sv2v_reg,data_o_65_sv2v_reg,
  data_o_64_sv2v_reg,data_o_63_sv2v_reg,data_o_62_sv2v_reg,data_o_61_sv2v_reg,
  data_o_60_sv2v_reg,data_o_59_sv2v_reg,data_o_58_sv2v_reg,data_o_57_sv2v_reg,
  data_o_56_sv2v_reg,data_o_55_sv2v_reg,data_o_54_sv2v_reg,data_o_53_sv2v_reg,
  data_o_52_sv2v_reg,data_o_51_sv2v_reg,data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,
  data_o_47_sv2v_reg,data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,
  data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,
  data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,
  data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,
  data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,
  data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,
  data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,
  data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,
  data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[89] = data_o_89_sv2v_reg;
  assign data_o[88] = data_o_88_sv2v_reg;
  assign data_o[87] = data_o_87_sv2v_reg;
  assign data_o[86] = data_o_86_sv2v_reg;
  assign data_o[85] = data_o_85_sv2v_reg;
  assign data_o[84] = data_o_84_sv2v_reg;
  assign data_o[83] = data_o_83_sv2v_reg;
  assign data_o[82] = data_o_82_sv2v_reg;
  assign data_o[81] = data_o_81_sv2v_reg;
  assign data_o[80] = data_o_80_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_89_sv2v_reg <= 1'b0;
      data_o_88_sv2v_reg <= 1'b0;
      data_o_87_sv2v_reg <= 1'b0;
      data_o_86_sv2v_reg <= 1'b0;
      data_o_85_sv2v_reg <= 1'b0;
      data_o_84_sv2v_reg <= 1'b0;
      data_o_83_sv2v_reg <= 1'b0;
      data_o_82_sv2v_reg <= 1'b0;
      data_o_81_sv2v_reg <= 1'b0;
      data_o_80_sv2v_reg <= 1'b0;
      data_o_79_sv2v_reg <= 1'b0;
      data_o_78_sv2v_reg <= 1'b0;
      data_o_77_sv2v_reg <= 1'b0;
      data_o_76_sv2v_reg <= 1'b0;
      data_o_75_sv2v_reg <= 1'b0;
      data_o_74_sv2v_reg <= 1'b0;
      data_o_73_sv2v_reg <= 1'b0;
      data_o_72_sv2v_reg <= 1'b0;
      data_o_71_sv2v_reg <= 1'b0;
      data_o_70_sv2v_reg <= 1'b0;
      data_o_69_sv2v_reg <= 1'b0;
      data_o_68_sv2v_reg <= 1'b0;
      data_o_67_sv2v_reg <= 1'b0;
      data_o_66_sv2v_reg <= 1'b0;
      data_o_65_sv2v_reg <= 1'b0;
      data_o_64_sv2v_reg <= 1'b0;
      data_o_63_sv2v_reg <= 1'b0;
      data_o_62_sv2v_reg <= 1'b0;
      data_o_61_sv2v_reg <= 1'b0;
      data_o_60_sv2v_reg <= 1'b0;
      data_o_59_sv2v_reg <= 1'b0;
      data_o_58_sv2v_reg <= 1'b0;
      data_o_57_sv2v_reg <= 1'b0;
      data_o_56_sv2v_reg <= 1'b0;
      data_o_55_sv2v_reg <= 1'b0;
      data_o_54_sv2v_reg <= 1'b0;
      data_o_53_sv2v_reg <= 1'b0;
      data_o_52_sv2v_reg <= 1'b0;
      data_o_51_sv2v_reg <= 1'b0;
      data_o_50_sv2v_reg <= 1'b0;
      data_o_49_sv2v_reg <= 1'b0;
      data_o_48_sv2v_reg <= 1'b0;
      data_o_47_sv2v_reg <= 1'b0;
      data_o_46_sv2v_reg <= 1'b0;
      data_o_45_sv2v_reg <= 1'b0;
      data_o_44_sv2v_reg <= 1'b0;
      data_o_43_sv2v_reg <= 1'b0;
      data_o_42_sv2v_reg <= 1'b0;
      data_o_41_sv2v_reg <= 1'b0;
      data_o_40_sv2v_reg <= 1'b0;
      data_o_39_sv2v_reg <= 1'b0;
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_89_sv2v_reg <= data_i[89];
      data_o_88_sv2v_reg <= data_i[88];
      data_o_87_sv2v_reg <= data_i[87];
      data_o_86_sv2v_reg <= data_i[86];
      data_o_85_sv2v_reg <= data_i[85];
      data_o_84_sv2v_reg <= data_i[84];
      data_o_83_sv2v_reg <= data_i[83];
      data_o_82_sv2v_reg <= data_i[82];
      data_o_81_sv2v_reg <= data_i[81];
      data_o_80_sv2v_reg <= data_i[80];
      data_o_79_sv2v_reg <= data_i[79];
      data_o_78_sv2v_reg <= data_i[78];
      data_o_77_sv2v_reg <= data_i[77];
      data_o_76_sv2v_reg <= data_i[76];
      data_o_75_sv2v_reg <= data_i[75];
      data_o_74_sv2v_reg <= data_i[74];
      data_o_73_sv2v_reg <= data_i[73];
      data_o_72_sv2v_reg <= data_i[72];
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_counter_clear_up_max_val_p16_init_val_p0
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [4:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire [4:0] count_o;
  wire N0,N1,N4,N5,N6,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N2,N3,N7,N30,N18;
  reg count_o_4_sv2v_reg,count_o_3_sv2v_reg,count_o_2_sv2v_reg,count_o_1_sv2v_reg,
  count_o_0_sv2v_reg;
  assign count_o[4] = count_o_4_sv2v_reg;
  assign count_o[3] = count_o_3_sv2v_reg;
  assign count_o[2] = count_o_2_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign N18 = reset_i | clear_i;
  assign { N10, N9, N8, N6, N5 } = count_o + 1'b1;
  assign N11 = (N0)? 1'b1 : 
               (N7)? 1'b1 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = clear_i;
  assign N13 = (N1)? 1'b1 : 
               (N30)? 1'b0 : 1'b0;
  assign N1 = up_i;
  assign N12 = (N0)? up_i : 
               (N7)? N5 : 1'b0;
  assign N4 = N17;
  assign N14 = ~reset_i;
  assign N15 = ~clear_i;
  assign N16 = N14 & N15;
  assign N17 = up_i & N16;
  assign N2 = up_i | clear_i;
  assign N3 = ~N2;
  assign N7 = up_i & N15;
  assign N30 = ~up_i;

  always @(posedge clk_i) begin
    if(N18) begin
      count_o_4_sv2v_reg <= 1'b0;
      count_o_3_sv2v_reg <= 1'b0;
      count_o_2_sv2v_reg <= 1'b0;
      count_o_1_sv2v_reg <= 1'b0;
    end else if(N13) begin
      count_o_4_sv2v_reg <= N10;
      count_o_3_sv2v_reg <= N9;
      count_o_2_sv2v_reg <= N8;
      count_o_1_sv2v_reg <= N6;
    end 
    if(reset_i) begin
      count_o_0_sv2v_reg <= 1'b0;
    end else if(N11) begin
      count_o_0_sv2v_reg <= N12;
    end 
  end


endmodule



module bsg_dff_reset_00000008
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [7:0] data_i;
  output [7:0] data_o;
  input clk_i;
  input reset_i;
  wire [7:0] data_o;
  reg data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_synth_0000002b_16_1
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [3:0] w_addr_i;
  input [42:0] w_data_i;
  input [3:0] r_addr_i;
  output [42:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [42:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82;
  wire [687:0] \nz.mem ;
  reg \nz.mem_687_sv2v_reg ,\nz.mem_686_sv2v_reg ,\nz.mem_685_sv2v_reg ,
  \nz.mem_684_sv2v_reg ,\nz.mem_683_sv2v_reg ,\nz.mem_682_sv2v_reg ,\nz.mem_681_sv2v_reg ,
  \nz.mem_680_sv2v_reg ,\nz.mem_679_sv2v_reg ,\nz.mem_678_sv2v_reg ,
  \nz.mem_677_sv2v_reg ,\nz.mem_676_sv2v_reg ,\nz.mem_675_sv2v_reg ,\nz.mem_674_sv2v_reg ,
  \nz.mem_673_sv2v_reg ,\nz.mem_672_sv2v_reg ,\nz.mem_671_sv2v_reg ,\nz.mem_670_sv2v_reg ,
  \nz.mem_669_sv2v_reg ,\nz.mem_668_sv2v_reg ,\nz.mem_667_sv2v_reg ,
  \nz.mem_666_sv2v_reg ,\nz.mem_665_sv2v_reg ,\nz.mem_664_sv2v_reg ,\nz.mem_663_sv2v_reg ,
  \nz.mem_662_sv2v_reg ,\nz.mem_661_sv2v_reg ,\nz.mem_660_sv2v_reg ,\nz.mem_659_sv2v_reg ,
  \nz.mem_658_sv2v_reg ,\nz.mem_657_sv2v_reg ,\nz.mem_656_sv2v_reg ,
  \nz.mem_655_sv2v_reg ,\nz.mem_654_sv2v_reg ,\nz.mem_653_sv2v_reg ,\nz.mem_652_sv2v_reg ,
  \nz.mem_651_sv2v_reg ,\nz.mem_650_sv2v_reg ,\nz.mem_649_sv2v_reg ,\nz.mem_648_sv2v_reg ,
  \nz.mem_647_sv2v_reg ,\nz.mem_646_sv2v_reg ,\nz.mem_645_sv2v_reg ,
  \nz.mem_644_sv2v_reg ,\nz.mem_643_sv2v_reg ,\nz.mem_642_sv2v_reg ,\nz.mem_641_sv2v_reg ,
  \nz.mem_640_sv2v_reg ,\nz.mem_639_sv2v_reg ,\nz.mem_638_sv2v_reg ,
  \nz.mem_637_sv2v_reg ,\nz.mem_636_sv2v_reg ,\nz.mem_635_sv2v_reg ,\nz.mem_634_sv2v_reg ,
  \nz.mem_633_sv2v_reg ,\nz.mem_632_sv2v_reg ,\nz.mem_631_sv2v_reg ,\nz.mem_630_sv2v_reg ,
  \nz.mem_629_sv2v_reg ,\nz.mem_628_sv2v_reg ,\nz.mem_627_sv2v_reg ,
  \nz.mem_626_sv2v_reg ,\nz.mem_625_sv2v_reg ,\nz.mem_624_sv2v_reg ,\nz.mem_623_sv2v_reg ,
  \nz.mem_622_sv2v_reg ,\nz.mem_621_sv2v_reg ,\nz.mem_620_sv2v_reg ,\nz.mem_619_sv2v_reg ,
  \nz.mem_618_sv2v_reg ,\nz.mem_617_sv2v_reg ,\nz.mem_616_sv2v_reg ,
  \nz.mem_615_sv2v_reg ,\nz.mem_614_sv2v_reg ,\nz.mem_613_sv2v_reg ,\nz.mem_612_sv2v_reg ,
  \nz.mem_611_sv2v_reg ,\nz.mem_610_sv2v_reg ,\nz.mem_609_sv2v_reg ,\nz.mem_608_sv2v_reg ,
  \nz.mem_607_sv2v_reg ,\nz.mem_606_sv2v_reg ,\nz.mem_605_sv2v_reg ,
  \nz.mem_604_sv2v_reg ,\nz.mem_603_sv2v_reg ,\nz.mem_602_sv2v_reg ,\nz.mem_601_sv2v_reg ,
  \nz.mem_600_sv2v_reg ,\nz.mem_599_sv2v_reg ,\nz.mem_598_sv2v_reg ,
  \nz.mem_597_sv2v_reg ,\nz.mem_596_sv2v_reg ,\nz.mem_595_sv2v_reg ,\nz.mem_594_sv2v_reg ,
  \nz.mem_593_sv2v_reg ,\nz.mem_592_sv2v_reg ,\nz.mem_591_sv2v_reg ,\nz.mem_590_sv2v_reg ,
  \nz.mem_589_sv2v_reg ,\nz.mem_588_sv2v_reg ,\nz.mem_587_sv2v_reg ,
  \nz.mem_586_sv2v_reg ,\nz.mem_585_sv2v_reg ,\nz.mem_584_sv2v_reg ,\nz.mem_583_sv2v_reg ,
  \nz.mem_582_sv2v_reg ,\nz.mem_581_sv2v_reg ,\nz.mem_580_sv2v_reg ,\nz.mem_579_sv2v_reg ,
  \nz.mem_578_sv2v_reg ,\nz.mem_577_sv2v_reg ,\nz.mem_576_sv2v_reg ,
  \nz.mem_575_sv2v_reg ,\nz.mem_574_sv2v_reg ,\nz.mem_573_sv2v_reg ,\nz.mem_572_sv2v_reg ,
  \nz.mem_571_sv2v_reg ,\nz.mem_570_sv2v_reg ,\nz.mem_569_sv2v_reg ,\nz.mem_568_sv2v_reg ,
  \nz.mem_567_sv2v_reg ,\nz.mem_566_sv2v_reg ,\nz.mem_565_sv2v_reg ,
  \nz.mem_564_sv2v_reg ,\nz.mem_563_sv2v_reg ,\nz.mem_562_sv2v_reg ,\nz.mem_561_sv2v_reg ,
  \nz.mem_560_sv2v_reg ,\nz.mem_559_sv2v_reg ,\nz.mem_558_sv2v_reg ,
  \nz.mem_557_sv2v_reg ,\nz.mem_556_sv2v_reg ,\nz.mem_555_sv2v_reg ,\nz.mem_554_sv2v_reg ,
  \nz.mem_553_sv2v_reg ,\nz.mem_552_sv2v_reg ,\nz.mem_551_sv2v_reg ,\nz.mem_550_sv2v_reg ,
  \nz.mem_549_sv2v_reg ,\nz.mem_548_sv2v_reg ,\nz.mem_547_sv2v_reg ,
  \nz.mem_546_sv2v_reg ,\nz.mem_545_sv2v_reg ,\nz.mem_544_sv2v_reg ,\nz.mem_543_sv2v_reg ,
  \nz.mem_542_sv2v_reg ,\nz.mem_541_sv2v_reg ,\nz.mem_540_sv2v_reg ,\nz.mem_539_sv2v_reg ,
  \nz.mem_538_sv2v_reg ,\nz.mem_537_sv2v_reg ,\nz.mem_536_sv2v_reg ,
  \nz.mem_535_sv2v_reg ,\nz.mem_534_sv2v_reg ,\nz.mem_533_sv2v_reg ,\nz.mem_532_sv2v_reg ,
  \nz.mem_531_sv2v_reg ,\nz.mem_530_sv2v_reg ,\nz.mem_529_sv2v_reg ,\nz.mem_528_sv2v_reg ,
  \nz.mem_527_sv2v_reg ,\nz.mem_526_sv2v_reg ,\nz.mem_525_sv2v_reg ,
  \nz.mem_524_sv2v_reg ,\nz.mem_523_sv2v_reg ,\nz.mem_522_sv2v_reg ,\nz.mem_521_sv2v_reg ,
  \nz.mem_520_sv2v_reg ,\nz.mem_519_sv2v_reg ,\nz.mem_518_sv2v_reg ,
  \nz.mem_517_sv2v_reg ,\nz.mem_516_sv2v_reg ,\nz.mem_515_sv2v_reg ,\nz.mem_514_sv2v_reg ,
  \nz.mem_513_sv2v_reg ,\nz.mem_512_sv2v_reg ,\nz.mem_511_sv2v_reg ,\nz.mem_510_sv2v_reg ,
  \nz.mem_509_sv2v_reg ,\nz.mem_508_sv2v_reg ,\nz.mem_507_sv2v_reg ,
  \nz.mem_506_sv2v_reg ,\nz.mem_505_sv2v_reg ,\nz.mem_504_sv2v_reg ,\nz.mem_503_sv2v_reg ,
  \nz.mem_502_sv2v_reg ,\nz.mem_501_sv2v_reg ,\nz.mem_500_sv2v_reg ,\nz.mem_499_sv2v_reg ,
  \nz.mem_498_sv2v_reg ,\nz.mem_497_sv2v_reg ,\nz.mem_496_sv2v_reg ,
  \nz.mem_495_sv2v_reg ,\nz.mem_494_sv2v_reg ,\nz.mem_493_sv2v_reg ,\nz.mem_492_sv2v_reg ,
  \nz.mem_491_sv2v_reg ,\nz.mem_490_sv2v_reg ,\nz.mem_489_sv2v_reg ,\nz.mem_488_sv2v_reg ,
  \nz.mem_487_sv2v_reg ,\nz.mem_486_sv2v_reg ,\nz.mem_485_sv2v_reg ,
  \nz.mem_484_sv2v_reg ,\nz.mem_483_sv2v_reg ,\nz.mem_482_sv2v_reg ,\nz.mem_481_sv2v_reg ,
  \nz.mem_480_sv2v_reg ,\nz.mem_479_sv2v_reg ,\nz.mem_478_sv2v_reg ,
  \nz.mem_477_sv2v_reg ,\nz.mem_476_sv2v_reg ,\nz.mem_475_sv2v_reg ,\nz.mem_474_sv2v_reg ,
  \nz.mem_473_sv2v_reg ,\nz.mem_472_sv2v_reg ,\nz.mem_471_sv2v_reg ,\nz.mem_470_sv2v_reg ,
  \nz.mem_469_sv2v_reg ,\nz.mem_468_sv2v_reg ,\nz.mem_467_sv2v_reg ,
  \nz.mem_466_sv2v_reg ,\nz.mem_465_sv2v_reg ,\nz.mem_464_sv2v_reg ,\nz.mem_463_sv2v_reg ,
  \nz.mem_462_sv2v_reg ,\nz.mem_461_sv2v_reg ,\nz.mem_460_sv2v_reg ,\nz.mem_459_sv2v_reg ,
  \nz.mem_458_sv2v_reg ,\nz.mem_457_sv2v_reg ,\nz.mem_456_sv2v_reg ,
  \nz.mem_455_sv2v_reg ,\nz.mem_454_sv2v_reg ,\nz.mem_453_sv2v_reg ,\nz.mem_452_sv2v_reg ,
  \nz.mem_451_sv2v_reg ,\nz.mem_450_sv2v_reg ,\nz.mem_449_sv2v_reg ,\nz.mem_448_sv2v_reg ,
  \nz.mem_447_sv2v_reg ,\nz.mem_446_sv2v_reg ,\nz.mem_445_sv2v_reg ,
  \nz.mem_444_sv2v_reg ,\nz.mem_443_sv2v_reg ,\nz.mem_442_sv2v_reg ,\nz.mem_441_sv2v_reg ,
  \nz.mem_440_sv2v_reg ,\nz.mem_439_sv2v_reg ,\nz.mem_438_sv2v_reg ,
  \nz.mem_437_sv2v_reg ,\nz.mem_436_sv2v_reg ,\nz.mem_435_sv2v_reg ,\nz.mem_434_sv2v_reg ,
  \nz.mem_433_sv2v_reg ,\nz.mem_432_sv2v_reg ,\nz.mem_431_sv2v_reg ,\nz.mem_430_sv2v_reg ,
  \nz.mem_429_sv2v_reg ,\nz.mem_428_sv2v_reg ,\nz.mem_427_sv2v_reg ,
  \nz.mem_426_sv2v_reg ,\nz.mem_425_sv2v_reg ,\nz.mem_424_sv2v_reg ,\nz.mem_423_sv2v_reg ,
  \nz.mem_422_sv2v_reg ,\nz.mem_421_sv2v_reg ,\nz.mem_420_sv2v_reg ,\nz.mem_419_sv2v_reg ,
  \nz.mem_418_sv2v_reg ,\nz.mem_417_sv2v_reg ,\nz.mem_416_sv2v_reg ,
  \nz.mem_415_sv2v_reg ,\nz.mem_414_sv2v_reg ,\nz.mem_413_sv2v_reg ,\nz.mem_412_sv2v_reg ,
  \nz.mem_411_sv2v_reg ,\nz.mem_410_sv2v_reg ,\nz.mem_409_sv2v_reg ,\nz.mem_408_sv2v_reg ,
  \nz.mem_407_sv2v_reg ,\nz.mem_406_sv2v_reg ,\nz.mem_405_sv2v_reg ,
  \nz.mem_404_sv2v_reg ,\nz.mem_403_sv2v_reg ,\nz.mem_402_sv2v_reg ,\nz.mem_401_sv2v_reg ,
  \nz.mem_400_sv2v_reg ,\nz.mem_399_sv2v_reg ,\nz.mem_398_sv2v_reg ,
  \nz.mem_397_sv2v_reg ,\nz.mem_396_sv2v_reg ,\nz.mem_395_sv2v_reg ,\nz.mem_394_sv2v_reg ,
  \nz.mem_393_sv2v_reg ,\nz.mem_392_sv2v_reg ,\nz.mem_391_sv2v_reg ,\nz.mem_390_sv2v_reg ,
  \nz.mem_389_sv2v_reg ,\nz.mem_388_sv2v_reg ,\nz.mem_387_sv2v_reg ,
  \nz.mem_386_sv2v_reg ,\nz.mem_385_sv2v_reg ,\nz.mem_384_sv2v_reg ,\nz.mem_383_sv2v_reg ,
  \nz.mem_382_sv2v_reg ,\nz.mem_381_sv2v_reg ,\nz.mem_380_sv2v_reg ,\nz.mem_379_sv2v_reg ,
  \nz.mem_378_sv2v_reg ,\nz.mem_377_sv2v_reg ,\nz.mem_376_sv2v_reg ,
  \nz.mem_375_sv2v_reg ,\nz.mem_374_sv2v_reg ,\nz.mem_373_sv2v_reg ,\nz.mem_372_sv2v_reg ,
  \nz.mem_371_sv2v_reg ,\nz.mem_370_sv2v_reg ,\nz.mem_369_sv2v_reg ,\nz.mem_368_sv2v_reg ,
  \nz.mem_367_sv2v_reg ,\nz.mem_366_sv2v_reg ,\nz.mem_365_sv2v_reg ,
  \nz.mem_364_sv2v_reg ,\nz.mem_363_sv2v_reg ,\nz.mem_362_sv2v_reg ,\nz.mem_361_sv2v_reg ,
  \nz.mem_360_sv2v_reg ,\nz.mem_359_sv2v_reg ,\nz.mem_358_sv2v_reg ,
  \nz.mem_357_sv2v_reg ,\nz.mem_356_sv2v_reg ,\nz.mem_355_sv2v_reg ,\nz.mem_354_sv2v_reg ,
  \nz.mem_353_sv2v_reg ,\nz.mem_352_sv2v_reg ,\nz.mem_351_sv2v_reg ,\nz.mem_350_sv2v_reg ,
  \nz.mem_349_sv2v_reg ,\nz.mem_348_sv2v_reg ,\nz.mem_347_sv2v_reg ,
  \nz.mem_346_sv2v_reg ,\nz.mem_345_sv2v_reg ,\nz.mem_344_sv2v_reg ,\nz.mem_343_sv2v_reg ,
  \nz.mem_342_sv2v_reg ,\nz.mem_341_sv2v_reg ,\nz.mem_340_sv2v_reg ,\nz.mem_339_sv2v_reg ,
  \nz.mem_338_sv2v_reg ,\nz.mem_337_sv2v_reg ,\nz.mem_336_sv2v_reg ,
  \nz.mem_335_sv2v_reg ,\nz.mem_334_sv2v_reg ,\nz.mem_333_sv2v_reg ,\nz.mem_332_sv2v_reg ,
  \nz.mem_331_sv2v_reg ,\nz.mem_330_sv2v_reg ,\nz.mem_329_sv2v_reg ,\nz.mem_328_sv2v_reg ,
  \nz.mem_327_sv2v_reg ,\nz.mem_326_sv2v_reg ,\nz.mem_325_sv2v_reg ,
  \nz.mem_324_sv2v_reg ,\nz.mem_323_sv2v_reg ,\nz.mem_322_sv2v_reg ,\nz.mem_321_sv2v_reg ,
  \nz.mem_320_sv2v_reg ,\nz.mem_319_sv2v_reg ,\nz.mem_318_sv2v_reg ,
  \nz.mem_317_sv2v_reg ,\nz.mem_316_sv2v_reg ,\nz.mem_315_sv2v_reg ,\nz.mem_314_sv2v_reg ,
  \nz.mem_313_sv2v_reg ,\nz.mem_312_sv2v_reg ,\nz.mem_311_sv2v_reg ,\nz.mem_310_sv2v_reg ,
  \nz.mem_309_sv2v_reg ,\nz.mem_308_sv2v_reg ,\nz.mem_307_sv2v_reg ,
  \nz.mem_306_sv2v_reg ,\nz.mem_305_sv2v_reg ,\nz.mem_304_sv2v_reg ,\nz.mem_303_sv2v_reg ,
  \nz.mem_302_sv2v_reg ,\nz.mem_301_sv2v_reg ,\nz.mem_300_sv2v_reg ,\nz.mem_299_sv2v_reg ,
  \nz.mem_298_sv2v_reg ,\nz.mem_297_sv2v_reg ,\nz.mem_296_sv2v_reg ,
  \nz.mem_295_sv2v_reg ,\nz.mem_294_sv2v_reg ,\nz.mem_293_sv2v_reg ,\nz.mem_292_sv2v_reg ,
  \nz.mem_291_sv2v_reg ,\nz.mem_290_sv2v_reg ,\nz.mem_289_sv2v_reg ,\nz.mem_288_sv2v_reg ,
  \nz.mem_287_sv2v_reg ,\nz.mem_286_sv2v_reg ,\nz.mem_285_sv2v_reg ,
  \nz.mem_284_sv2v_reg ,\nz.mem_283_sv2v_reg ,\nz.mem_282_sv2v_reg ,\nz.mem_281_sv2v_reg ,
  \nz.mem_280_sv2v_reg ,\nz.mem_279_sv2v_reg ,\nz.mem_278_sv2v_reg ,
  \nz.mem_277_sv2v_reg ,\nz.mem_276_sv2v_reg ,\nz.mem_275_sv2v_reg ,\nz.mem_274_sv2v_reg ,
  \nz.mem_273_sv2v_reg ,\nz.mem_272_sv2v_reg ,\nz.mem_271_sv2v_reg ,\nz.mem_270_sv2v_reg ,
  \nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,\nz.mem_267_sv2v_reg ,
  \nz.mem_266_sv2v_reg ,\nz.mem_265_sv2v_reg ,\nz.mem_264_sv2v_reg ,\nz.mem_263_sv2v_reg ,
  \nz.mem_262_sv2v_reg ,\nz.mem_261_sv2v_reg ,\nz.mem_260_sv2v_reg ,\nz.mem_259_sv2v_reg ,
  \nz.mem_258_sv2v_reg ,\nz.mem_257_sv2v_reg ,\nz.mem_256_sv2v_reg ,
  \nz.mem_255_sv2v_reg ,\nz.mem_254_sv2v_reg ,\nz.mem_253_sv2v_reg ,\nz.mem_252_sv2v_reg ,
  \nz.mem_251_sv2v_reg ,\nz.mem_250_sv2v_reg ,\nz.mem_249_sv2v_reg ,\nz.mem_248_sv2v_reg ,
  \nz.mem_247_sv2v_reg ,\nz.mem_246_sv2v_reg ,\nz.mem_245_sv2v_reg ,
  \nz.mem_244_sv2v_reg ,\nz.mem_243_sv2v_reg ,\nz.mem_242_sv2v_reg ,\nz.mem_241_sv2v_reg ,
  \nz.mem_240_sv2v_reg ,\nz.mem_239_sv2v_reg ,\nz.mem_238_sv2v_reg ,
  \nz.mem_237_sv2v_reg ,\nz.mem_236_sv2v_reg ,\nz.mem_235_sv2v_reg ,\nz.mem_234_sv2v_reg ,
  \nz.mem_233_sv2v_reg ,\nz.mem_232_sv2v_reg ,\nz.mem_231_sv2v_reg ,\nz.mem_230_sv2v_reg ,
  \nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,\nz.mem_227_sv2v_reg ,
  \nz.mem_226_sv2v_reg ,\nz.mem_225_sv2v_reg ,\nz.mem_224_sv2v_reg ,\nz.mem_223_sv2v_reg ,
  \nz.mem_222_sv2v_reg ,\nz.mem_221_sv2v_reg ,\nz.mem_220_sv2v_reg ,\nz.mem_219_sv2v_reg ,
  \nz.mem_218_sv2v_reg ,\nz.mem_217_sv2v_reg ,\nz.mem_216_sv2v_reg ,
  \nz.mem_215_sv2v_reg ,\nz.mem_214_sv2v_reg ,\nz.mem_213_sv2v_reg ,\nz.mem_212_sv2v_reg ,
  \nz.mem_211_sv2v_reg ,\nz.mem_210_sv2v_reg ,\nz.mem_209_sv2v_reg ,\nz.mem_208_sv2v_reg ,
  \nz.mem_207_sv2v_reg ,\nz.mem_206_sv2v_reg ,\nz.mem_205_sv2v_reg ,
  \nz.mem_204_sv2v_reg ,\nz.mem_203_sv2v_reg ,\nz.mem_202_sv2v_reg ,\nz.mem_201_sv2v_reg ,
  \nz.mem_200_sv2v_reg ,\nz.mem_199_sv2v_reg ,\nz.mem_198_sv2v_reg ,
  \nz.mem_197_sv2v_reg ,\nz.mem_196_sv2v_reg ,\nz.mem_195_sv2v_reg ,\nz.mem_194_sv2v_reg ,
  \nz.mem_193_sv2v_reg ,\nz.mem_192_sv2v_reg ,\nz.mem_191_sv2v_reg ,\nz.mem_190_sv2v_reg ,
  \nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,\nz.mem_187_sv2v_reg ,
  \nz.mem_186_sv2v_reg ,\nz.mem_185_sv2v_reg ,\nz.mem_184_sv2v_reg ,\nz.mem_183_sv2v_reg ,
  \nz.mem_182_sv2v_reg ,\nz.mem_181_sv2v_reg ,\nz.mem_180_sv2v_reg ,\nz.mem_179_sv2v_reg ,
  \nz.mem_178_sv2v_reg ,\nz.mem_177_sv2v_reg ,\nz.mem_176_sv2v_reg ,
  \nz.mem_175_sv2v_reg ,\nz.mem_174_sv2v_reg ,\nz.mem_173_sv2v_reg ,\nz.mem_172_sv2v_reg ,
  \nz.mem_171_sv2v_reg ,\nz.mem_170_sv2v_reg ,\nz.mem_169_sv2v_reg ,\nz.mem_168_sv2v_reg ,
  \nz.mem_167_sv2v_reg ,\nz.mem_166_sv2v_reg ,\nz.mem_165_sv2v_reg ,
  \nz.mem_164_sv2v_reg ,\nz.mem_163_sv2v_reg ,\nz.mem_162_sv2v_reg ,\nz.mem_161_sv2v_reg ,
  \nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,\nz.mem_158_sv2v_reg ,
  \nz.mem_157_sv2v_reg ,\nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,\nz.mem_154_sv2v_reg ,
  \nz.mem_153_sv2v_reg ,\nz.mem_152_sv2v_reg ,\nz.mem_151_sv2v_reg ,\nz.mem_150_sv2v_reg ,
  \nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,\nz.mem_147_sv2v_reg ,
  \nz.mem_146_sv2v_reg ,\nz.mem_145_sv2v_reg ,\nz.mem_144_sv2v_reg ,\nz.mem_143_sv2v_reg ,
  \nz.mem_142_sv2v_reg ,\nz.mem_141_sv2v_reg ,\nz.mem_140_sv2v_reg ,\nz.mem_139_sv2v_reg ,
  \nz.mem_138_sv2v_reg ,\nz.mem_137_sv2v_reg ,\nz.mem_136_sv2v_reg ,
  \nz.mem_135_sv2v_reg ,\nz.mem_134_sv2v_reg ,\nz.mem_133_sv2v_reg ,\nz.mem_132_sv2v_reg ,
  \nz.mem_131_sv2v_reg ,\nz.mem_130_sv2v_reg ,\nz.mem_129_sv2v_reg ,\nz.mem_128_sv2v_reg ,
  \nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,\nz.mem_125_sv2v_reg ,
  \nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,\nz.mem_122_sv2v_reg ,\nz.mem_121_sv2v_reg ,
  \nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,\nz.mem_118_sv2v_reg ,
  \nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,\nz.mem_114_sv2v_reg ,
  \nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,\nz.mem_111_sv2v_reg ,\nz.mem_110_sv2v_reg ,
  \nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,\nz.mem_107_sv2v_reg ,
  \nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,\nz.mem_103_sv2v_reg ,
  \nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,\nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,
  \nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,\nz.mem_96_sv2v_reg ,
  \nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,\nz.mem_92_sv2v_reg ,
  \nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,\nz.mem_88_sv2v_reg ,
  \nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,
  \nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,\nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,
  \nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,\nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,
  \nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,\nz.mem_73_sv2v_reg ,
  \nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,\nz.mem_69_sv2v_reg ,
  \nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,
  \nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,
  \nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,
  \nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,
  \nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,
  \nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,
  \nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,
  \nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,
  \nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,
  \nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,
  \nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,
  \nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,
  \nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,
  \nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,
  \nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,
  \nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,
  \nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,
  \nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.mem [687] = \nz.mem_687_sv2v_reg ;
  assign \nz.mem [686] = \nz.mem_686_sv2v_reg ;
  assign \nz.mem [685] = \nz.mem_685_sv2v_reg ;
  assign \nz.mem [684] = \nz.mem_684_sv2v_reg ;
  assign \nz.mem [683] = \nz.mem_683_sv2v_reg ;
  assign \nz.mem [682] = \nz.mem_682_sv2v_reg ;
  assign \nz.mem [681] = \nz.mem_681_sv2v_reg ;
  assign \nz.mem [680] = \nz.mem_680_sv2v_reg ;
  assign \nz.mem [679] = \nz.mem_679_sv2v_reg ;
  assign \nz.mem [678] = \nz.mem_678_sv2v_reg ;
  assign \nz.mem [677] = \nz.mem_677_sv2v_reg ;
  assign \nz.mem [676] = \nz.mem_676_sv2v_reg ;
  assign \nz.mem [675] = \nz.mem_675_sv2v_reg ;
  assign \nz.mem [674] = \nz.mem_674_sv2v_reg ;
  assign \nz.mem [673] = \nz.mem_673_sv2v_reg ;
  assign \nz.mem [672] = \nz.mem_672_sv2v_reg ;
  assign \nz.mem [671] = \nz.mem_671_sv2v_reg ;
  assign \nz.mem [670] = \nz.mem_670_sv2v_reg ;
  assign \nz.mem [669] = \nz.mem_669_sv2v_reg ;
  assign \nz.mem [668] = \nz.mem_668_sv2v_reg ;
  assign \nz.mem [667] = \nz.mem_667_sv2v_reg ;
  assign \nz.mem [666] = \nz.mem_666_sv2v_reg ;
  assign \nz.mem [665] = \nz.mem_665_sv2v_reg ;
  assign \nz.mem [664] = \nz.mem_664_sv2v_reg ;
  assign \nz.mem [663] = \nz.mem_663_sv2v_reg ;
  assign \nz.mem [662] = \nz.mem_662_sv2v_reg ;
  assign \nz.mem [661] = \nz.mem_661_sv2v_reg ;
  assign \nz.mem [660] = \nz.mem_660_sv2v_reg ;
  assign \nz.mem [659] = \nz.mem_659_sv2v_reg ;
  assign \nz.mem [658] = \nz.mem_658_sv2v_reg ;
  assign \nz.mem [657] = \nz.mem_657_sv2v_reg ;
  assign \nz.mem [656] = \nz.mem_656_sv2v_reg ;
  assign \nz.mem [655] = \nz.mem_655_sv2v_reg ;
  assign \nz.mem [654] = \nz.mem_654_sv2v_reg ;
  assign \nz.mem [653] = \nz.mem_653_sv2v_reg ;
  assign \nz.mem [652] = \nz.mem_652_sv2v_reg ;
  assign \nz.mem [651] = \nz.mem_651_sv2v_reg ;
  assign \nz.mem [650] = \nz.mem_650_sv2v_reg ;
  assign \nz.mem [649] = \nz.mem_649_sv2v_reg ;
  assign \nz.mem [648] = \nz.mem_648_sv2v_reg ;
  assign \nz.mem [647] = \nz.mem_647_sv2v_reg ;
  assign \nz.mem [646] = \nz.mem_646_sv2v_reg ;
  assign \nz.mem [645] = \nz.mem_645_sv2v_reg ;
  assign \nz.mem [644] = \nz.mem_644_sv2v_reg ;
  assign \nz.mem [643] = \nz.mem_643_sv2v_reg ;
  assign \nz.mem [642] = \nz.mem_642_sv2v_reg ;
  assign \nz.mem [641] = \nz.mem_641_sv2v_reg ;
  assign \nz.mem [640] = \nz.mem_640_sv2v_reg ;
  assign \nz.mem [639] = \nz.mem_639_sv2v_reg ;
  assign \nz.mem [638] = \nz.mem_638_sv2v_reg ;
  assign \nz.mem [637] = \nz.mem_637_sv2v_reg ;
  assign \nz.mem [636] = \nz.mem_636_sv2v_reg ;
  assign \nz.mem [635] = \nz.mem_635_sv2v_reg ;
  assign \nz.mem [634] = \nz.mem_634_sv2v_reg ;
  assign \nz.mem [633] = \nz.mem_633_sv2v_reg ;
  assign \nz.mem [632] = \nz.mem_632_sv2v_reg ;
  assign \nz.mem [631] = \nz.mem_631_sv2v_reg ;
  assign \nz.mem [630] = \nz.mem_630_sv2v_reg ;
  assign \nz.mem [629] = \nz.mem_629_sv2v_reg ;
  assign \nz.mem [628] = \nz.mem_628_sv2v_reg ;
  assign \nz.mem [627] = \nz.mem_627_sv2v_reg ;
  assign \nz.mem [626] = \nz.mem_626_sv2v_reg ;
  assign \nz.mem [625] = \nz.mem_625_sv2v_reg ;
  assign \nz.mem [624] = \nz.mem_624_sv2v_reg ;
  assign \nz.mem [623] = \nz.mem_623_sv2v_reg ;
  assign \nz.mem [622] = \nz.mem_622_sv2v_reg ;
  assign \nz.mem [621] = \nz.mem_621_sv2v_reg ;
  assign \nz.mem [620] = \nz.mem_620_sv2v_reg ;
  assign \nz.mem [619] = \nz.mem_619_sv2v_reg ;
  assign \nz.mem [618] = \nz.mem_618_sv2v_reg ;
  assign \nz.mem [617] = \nz.mem_617_sv2v_reg ;
  assign \nz.mem [616] = \nz.mem_616_sv2v_reg ;
  assign \nz.mem [615] = \nz.mem_615_sv2v_reg ;
  assign \nz.mem [614] = \nz.mem_614_sv2v_reg ;
  assign \nz.mem [613] = \nz.mem_613_sv2v_reg ;
  assign \nz.mem [612] = \nz.mem_612_sv2v_reg ;
  assign \nz.mem [611] = \nz.mem_611_sv2v_reg ;
  assign \nz.mem [610] = \nz.mem_610_sv2v_reg ;
  assign \nz.mem [609] = \nz.mem_609_sv2v_reg ;
  assign \nz.mem [608] = \nz.mem_608_sv2v_reg ;
  assign \nz.mem [607] = \nz.mem_607_sv2v_reg ;
  assign \nz.mem [606] = \nz.mem_606_sv2v_reg ;
  assign \nz.mem [605] = \nz.mem_605_sv2v_reg ;
  assign \nz.mem [604] = \nz.mem_604_sv2v_reg ;
  assign \nz.mem [603] = \nz.mem_603_sv2v_reg ;
  assign \nz.mem [602] = \nz.mem_602_sv2v_reg ;
  assign \nz.mem [601] = \nz.mem_601_sv2v_reg ;
  assign \nz.mem [600] = \nz.mem_600_sv2v_reg ;
  assign \nz.mem [599] = \nz.mem_599_sv2v_reg ;
  assign \nz.mem [598] = \nz.mem_598_sv2v_reg ;
  assign \nz.mem [597] = \nz.mem_597_sv2v_reg ;
  assign \nz.mem [596] = \nz.mem_596_sv2v_reg ;
  assign \nz.mem [595] = \nz.mem_595_sv2v_reg ;
  assign \nz.mem [594] = \nz.mem_594_sv2v_reg ;
  assign \nz.mem [593] = \nz.mem_593_sv2v_reg ;
  assign \nz.mem [592] = \nz.mem_592_sv2v_reg ;
  assign \nz.mem [591] = \nz.mem_591_sv2v_reg ;
  assign \nz.mem [590] = \nz.mem_590_sv2v_reg ;
  assign \nz.mem [589] = \nz.mem_589_sv2v_reg ;
  assign \nz.mem [588] = \nz.mem_588_sv2v_reg ;
  assign \nz.mem [587] = \nz.mem_587_sv2v_reg ;
  assign \nz.mem [586] = \nz.mem_586_sv2v_reg ;
  assign \nz.mem [585] = \nz.mem_585_sv2v_reg ;
  assign \nz.mem [584] = \nz.mem_584_sv2v_reg ;
  assign \nz.mem [583] = \nz.mem_583_sv2v_reg ;
  assign \nz.mem [582] = \nz.mem_582_sv2v_reg ;
  assign \nz.mem [581] = \nz.mem_581_sv2v_reg ;
  assign \nz.mem [580] = \nz.mem_580_sv2v_reg ;
  assign \nz.mem [579] = \nz.mem_579_sv2v_reg ;
  assign \nz.mem [578] = \nz.mem_578_sv2v_reg ;
  assign \nz.mem [577] = \nz.mem_577_sv2v_reg ;
  assign \nz.mem [576] = \nz.mem_576_sv2v_reg ;
  assign \nz.mem [575] = \nz.mem_575_sv2v_reg ;
  assign \nz.mem [574] = \nz.mem_574_sv2v_reg ;
  assign \nz.mem [573] = \nz.mem_573_sv2v_reg ;
  assign \nz.mem [572] = \nz.mem_572_sv2v_reg ;
  assign \nz.mem [571] = \nz.mem_571_sv2v_reg ;
  assign \nz.mem [570] = \nz.mem_570_sv2v_reg ;
  assign \nz.mem [569] = \nz.mem_569_sv2v_reg ;
  assign \nz.mem [568] = \nz.mem_568_sv2v_reg ;
  assign \nz.mem [567] = \nz.mem_567_sv2v_reg ;
  assign \nz.mem [566] = \nz.mem_566_sv2v_reg ;
  assign \nz.mem [565] = \nz.mem_565_sv2v_reg ;
  assign \nz.mem [564] = \nz.mem_564_sv2v_reg ;
  assign \nz.mem [563] = \nz.mem_563_sv2v_reg ;
  assign \nz.mem [562] = \nz.mem_562_sv2v_reg ;
  assign \nz.mem [561] = \nz.mem_561_sv2v_reg ;
  assign \nz.mem [560] = \nz.mem_560_sv2v_reg ;
  assign \nz.mem [559] = \nz.mem_559_sv2v_reg ;
  assign \nz.mem [558] = \nz.mem_558_sv2v_reg ;
  assign \nz.mem [557] = \nz.mem_557_sv2v_reg ;
  assign \nz.mem [556] = \nz.mem_556_sv2v_reg ;
  assign \nz.mem [555] = \nz.mem_555_sv2v_reg ;
  assign \nz.mem [554] = \nz.mem_554_sv2v_reg ;
  assign \nz.mem [553] = \nz.mem_553_sv2v_reg ;
  assign \nz.mem [552] = \nz.mem_552_sv2v_reg ;
  assign \nz.mem [551] = \nz.mem_551_sv2v_reg ;
  assign \nz.mem [550] = \nz.mem_550_sv2v_reg ;
  assign \nz.mem [549] = \nz.mem_549_sv2v_reg ;
  assign \nz.mem [548] = \nz.mem_548_sv2v_reg ;
  assign \nz.mem [547] = \nz.mem_547_sv2v_reg ;
  assign \nz.mem [546] = \nz.mem_546_sv2v_reg ;
  assign \nz.mem [545] = \nz.mem_545_sv2v_reg ;
  assign \nz.mem [544] = \nz.mem_544_sv2v_reg ;
  assign \nz.mem [543] = \nz.mem_543_sv2v_reg ;
  assign \nz.mem [542] = \nz.mem_542_sv2v_reg ;
  assign \nz.mem [541] = \nz.mem_541_sv2v_reg ;
  assign \nz.mem [540] = \nz.mem_540_sv2v_reg ;
  assign \nz.mem [539] = \nz.mem_539_sv2v_reg ;
  assign \nz.mem [538] = \nz.mem_538_sv2v_reg ;
  assign \nz.mem [537] = \nz.mem_537_sv2v_reg ;
  assign \nz.mem [536] = \nz.mem_536_sv2v_reg ;
  assign \nz.mem [535] = \nz.mem_535_sv2v_reg ;
  assign \nz.mem [534] = \nz.mem_534_sv2v_reg ;
  assign \nz.mem [533] = \nz.mem_533_sv2v_reg ;
  assign \nz.mem [532] = \nz.mem_532_sv2v_reg ;
  assign \nz.mem [531] = \nz.mem_531_sv2v_reg ;
  assign \nz.mem [530] = \nz.mem_530_sv2v_reg ;
  assign \nz.mem [529] = \nz.mem_529_sv2v_reg ;
  assign \nz.mem [528] = \nz.mem_528_sv2v_reg ;
  assign \nz.mem [527] = \nz.mem_527_sv2v_reg ;
  assign \nz.mem [526] = \nz.mem_526_sv2v_reg ;
  assign \nz.mem [525] = \nz.mem_525_sv2v_reg ;
  assign \nz.mem [524] = \nz.mem_524_sv2v_reg ;
  assign \nz.mem [523] = \nz.mem_523_sv2v_reg ;
  assign \nz.mem [522] = \nz.mem_522_sv2v_reg ;
  assign \nz.mem [521] = \nz.mem_521_sv2v_reg ;
  assign \nz.mem [520] = \nz.mem_520_sv2v_reg ;
  assign \nz.mem [519] = \nz.mem_519_sv2v_reg ;
  assign \nz.mem [518] = \nz.mem_518_sv2v_reg ;
  assign \nz.mem [517] = \nz.mem_517_sv2v_reg ;
  assign \nz.mem [516] = \nz.mem_516_sv2v_reg ;
  assign \nz.mem [515] = \nz.mem_515_sv2v_reg ;
  assign \nz.mem [514] = \nz.mem_514_sv2v_reg ;
  assign \nz.mem [513] = \nz.mem_513_sv2v_reg ;
  assign \nz.mem [512] = \nz.mem_512_sv2v_reg ;
  assign \nz.mem [511] = \nz.mem_511_sv2v_reg ;
  assign \nz.mem [510] = \nz.mem_510_sv2v_reg ;
  assign \nz.mem [509] = \nz.mem_509_sv2v_reg ;
  assign \nz.mem [508] = \nz.mem_508_sv2v_reg ;
  assign \nz.mem [507] = \nz.mem_507_sv2v_reg ;
  assign \nz.mem [506] = \nz.mem_506_sv2v_reg ;
  assign \nz.mem [505] = \nz.mem_505_sv2v_reg ;
  assign \nz.mem [504] = \nz.mem_504_sv2v_reg ;
  assign \nz.mem [503] = \nz.mem_503_sv2v_reg ;
  assign \nz.mem [502] = \nz.mem_502_sv2v_reg ;
  assign \nz.mem [501] = \nz.mem_501_sv2v_reg ;
  assign \nz.mem [500] = \nz.mem_500_sv2v_reg ;
  assign \nz.mem [499] = \nz.mem_499_sv2v_reg ;
  assign \nz.mem [498] = \nz.mem_498_sv2v_reg ;
  assign \nz.mem [497] = \nz.mem_497_sv2v_reg ;
  assign \nz.mem [496] = \nz.mem_496_sv2v_reg ;
  assign \nz.mem [495] = \nz.mem_495_sv2v_reg ;
  assign \nz.mem [494] = \nz.mem_494_sv2v_reg ;
  assign \nz.mem [493] = \nz.mem_493_sv2v_reg ;
  assign \nz.mem [492] = \nz.mem_492_sv2v_reg ;
  assign \nz.mem [491] = \nz.mem_491_sv2v_reg ;
  assign \nz.mem [490] = \nz.mem_490_sv2v_reg ;
  assign \nz.mem [489] = \nz.mem_489_sv2v_reg ;
  assign \nz.mem [488] = \nz.mem_488_sv2v_reg ;
  assign \nz.mem [487] = \nz.mem_487_sv2v_reg ;
  assign \nz.mem [486] = \nz.mem_486_sv2v_reg ;
  assign \nz.mem [485] = \nz.mem_485_sv2v_reg ;
  assign \nz.mem [484] = \nz.mem_484_sv2v_reg ;
  assign \nz.mem [483] = \nz.mem_483_sv2v_reg ;
  assign \nz.mem [482] = \nz.mem_482_sv2v_reg ;
  assign \nz.mem [481] = \nz.mem_481_sv2v_reg ;
  assign \nz.mem [480] = \nz.mem_480_sv2v_reg ;
  assign \nz.mem [479] = \nz.mem_479_sv2v_reg ;
  assign \nz.mem [478] = \nz.mem_478_sv2v_reg ;
  assign \nz.mem [477] = \nz.mem_477_sv2v_reg ;
  assign \nz.mem [476] = \nz.mem_476_sv2v_reg ;
  assign \nz.mem [475] = \nz.mem_475_sv2v_reg ;
  assign \nz.mem [474] = \nz.mem_474_sv2v_reg ;
  assign \nz.mem [473] = \nz.mem_473_sv2v_reg ;
  assign \nz.mem [472] = \nz.mem_472_sv2v_reg ;
  assign \nz.mem [471] = \nz.mem_471_sv2v_reg ;
  assign \nz.mem [470] = \nz.mem_470_sv2v_reg ;
  assign \nz.mem [469] = \nz.mem_469_sv2v_reg ;
  assign \nz.mem [468] = \nz.mem_468_sv2v_reg ;
  assign \nz.mem [467] = \nz.mem_467_sv2v_reg ;
  assign \nz.mem [466] = \nz.mem_466_sv2v_reg ;
  assign \nz.mem [465] = \nz.mem_465_sv2v_reg ;
  assign \nz.mem [464] = \nz.mem_464_sv2v_reg ;
  assign \nz.mem [463] = \nz.mem_463_sv2v_reg ;
  assign \nz.mem [462] = \nz.mem_462_sv2v_reg ;
  assign \nz.mem [461] = \nz.mem_461_sv2v_reg ;
  assign \nz.mem [460] = \nz.mem_460_sv2v_reg ;
  assign \nz.mem [459] = \nz.mem_459_sv2v_reg ;
  assign \nz.mem [458] = \nz.mem_458_sv2v_reg ;
  assign \nz.mem [457] = \nz.mem_457_sv2v_reg ;
  assign \nz.mem [456] = \nz.mem_456_sv2v_reg ;
  assign \nz.mem [455] = \nz.mem_455_sv2v_reg ;
  assign \nz.mem [454] = \nz.mem_454_sv2v_reg ;
  assign \nz.mem [453] = \nz.mem_453_sv2v_reg ;
  assign \nz.mem [452] = \nz.mem_452_sv2v_reg ;
  assign \nz.mem [451] = \nz.mem_451_sv2v_reg ;
  assign \nz.mem [450] = \nz.mem_450_sv2v_reg ;
  assign \nz.mem [449] = \nz.mem_449_sv2v_reg ;
  assign \nz.mem [448] = \nz.mem_448_sv2v_reg ;
  assign \nz.mem [447] = \nz.mem_447_sv2v_reg ;
  assign \nz.mem [446] = \nz.mem_446_sv2v_reg ;
  assign \nz.mem [445] = \nz.mem_445_sv2v_reg ;
  assign \nz.mem [444] = \nz.mem_444_sv2v_reg ;
  assign \nz.mem [443] = \nz.mem_443_sv2v_reg ;
  assign \nz.mem [442] = \nz.mem_442_sv2v_reg ;
  assign \nz.mem [441] = \nz.mem_441_sv2v_reg ;
  assign \nz.mem [440] = \nz.mem_440_sv2v_reg ;
  assign \nz.mem [439] = \nz.mem_439_sv2v_reg ;
  assign \nz.mem [438] = \nz.mem_438_sv2v_reg ;
  assign \nz.mem [437] = \nz.mem_437_sv2v_reg ;
  assign \nz.mem [436] = \nz.mem_436_sv2v_reg ;
  assign \nz.mem [435] = \nz.mem_435_sv2v_reg ;
  assign \nz.mem [434] = \nz.mem_434_sv2v_reg ;
  assign \nz.mem [433] = \nz.mem_433_sv2v_reg ;
  assign \nz.mem [432] = \nz.mem_432_sv2v_reg ;
  assign \nz.mem [431] = \nz.mem_431_sv2v_reg ;
  assign \nz.mem [430] = \nz.mem_430_sv2v_reg ;
  assign \nz.mem [429] = \nz.mem_429_sv2v_reg ;
  assign \nz.mem [428] = \nz.mem_428_sv2v_reg ;
  assign \nz.mem [427] = \nz.mem_427_sv2v_reg ;
  assign \nz.mem [426] = \nz.mem_426_sv2v_reg ;
  assign \nz.mem [425] = \nz.mem_425_sv2v_reg ;
  assign \nz.mem [424] = \nz.mem_424_sv2v_reg ;
  assign \nz.mem [423] = \nz.mem_423_sv2v_reg ;
  assign \nz.mem [422] = \nz.mem_422_sv2v_reg ;
  assign \nz.mem [421] = \nz.mem_421_sv2v_reg ;
  assign \nz.mem [420] = \nz.mem_420_sv2v_reg ;
  assign \nz.mem [419] = \nz.mem_419_sv2v_reg ;
  assign \nz.mem [418] = \nz.mem_418_sv2v_reg ;
  assign \nz.mem [417] = \nz.mem_417_sv2v_reg ;
  assign \nz.mem [416] = \nz.mem_416_sv2v_reg ;
  assign \nz.mem [415] = \nz.mem_415_sv2v_reg ;
  assign \nz.mem [414] = \nz.mem_414_sv2v_reg ;
  assign \nz.mem [413] = \nz.mem_413_sv2v_reg ;
  assign \nz.mem [412] = \nz.mem_412_sv2v_reg ;
  assign \nz.mem [411] = \nz.mem_411_sv2v_reg ;
  assign \nz.mem [410] = \nz.mem_410_sv2v_reg ;
  assign \nz.mem [409] = \nz.mem_409_sv2v_reg ;
  assign \nz.mem [408] = \nz.mem_408_sv2v_reg ;
  assign \nz.mem [407] = \nz.mem_407_sv2v_reg ;
  assign \nz.mem [406] = \nz.mem_406_sv2v_reg ;
  assign \nz.mem [405] = \nz.mem_405_sv2v_reg ;
  assign \nz.mem [404] = \nz.mem_404_sv2v_reg ;
  assign \nz.mem [403] = \nz.mem_403_sv2v_reg ;
  assign \nz.mem [402] = \nz.mem_402_sv2v_reg ;
  assign \nz.mem [401] = \nz.mem_401_sv2v_reg ;
  assign \nz.mem [400] = \nz.mem_400_sv2v_reg ;
  assign \nz.mem [399] = \nz.mem_399_sv2v_reg ;
  assign \nz.mem [398] = \nz.mem_398_sv2v_reg ;
  assign \nz.mem [397] = \nz.mem_397_sv2v_reg ;
  assign \nz.mem [396] = \nz.mem_396_sv2v_reg ;
  assign \nz.mem [395] = \nz.mem_395_sv2v_reg ;
  assign \nz.mem [394] = \nz.mem_394_sv2v_reg ;
  assign \nz.mem [393] = \nz.mem_393_sv2v_reg ;
  assign \nz.mem [392] = \nz.mem_392_sv2v_reg ;
  assign \nz.mem [391] = \nz.mem_391_sv2v_reg ;
  assign \nz.mem [390] = \nz.mem_390_sv2v_reg ;
  assign \nz.mem [389] = \nz.mem_389_sv2v_reg ;
  assign \nz.mem [388] = \nz.mem_388_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[42] = (N26)? \nz.mem [42] : 
                        (N28)? \nz.mem [85] : 
                        (N30)? \nz.mem [128] : 
                        (N32)? \nz.mem [171] : 
                        (N34)? \nz.mem [214] : 
                        (N36)? \nz.mem [257] : 
                        (N38)? \nz.mem [300] : 
                        (N40)? \nz.mem [343] : 
                        (N27)? \nz.mem [386] : 
                        (N29)? \nz.mem [429] : 
                        (N31)? \nz.mem [472] : 
                        (N33)? \nz.mem [515] : 
                        (N35)? \nz.mem [558] : 
                        (N37)? \nz.mem [601] : 
                        (N39)? \nz.mem [644] : 
                        (N41)? \nz.mem [687] : 1'b0;
  assign r_data_o[41] = (N26)? \nz.mem [41] : 
                        (N28)? \nz.mem [84] : 
                        (N30)? \nz.mem [127] : 
                        (N32)? \nz.mem [170] : 
                        (N34)? \nz.mem [213] : 
                        (N36)? \nz.mem [256] : 
                        (N38)? \nz.mem [299] : 
                        (N40)? \nz.mem [342] : 
                        (N27)? \nz.mem [385] : 
                        (N29)? \nz.mem [428] : 
                        (N31)? \nz.mem [471] : 
                        (N33)? \nz.mem [514] : 
                        (N35)? \nz.mem [557] : 
                        (N37)? \nz.mem [600] : 
                        (N39)? \nz.mem [643] : 
                        (N41)? \nz.mem [686] : 1'b0;
  assign r_data_o[40] = (N26)? \nz.mem [40] : 
                        (N28)? \nz.mem [83] : 
                        (N30)? \nz.mem [126] : 
                        (N32)? \nz.mem [169] : 
                        (N34)? \nz.mem [212] : 
                        (N36)? \nz.mem [255] : 
                        (N38)? \nz.mem [298] : 
                        (N40)? \nz.mem [341] : 
                        (N27)? \nz.mem [384] : 
                        (N29)? \nz.mem [427] : 
                        (N31)? \nz.mem [470] : 
                        (N33)? \nz.mem [513] : 
                        (N35)? \nz.mem [556] : 
                        (N37)? \nz.mem [599] : 
                        (N39)? \nz.mem [642] : 
                        (N41)? \nz.mem [685] : 1'b0;
  assign r_data_o[39] = (N26)? \nz.mem [39] : 
                        (N28)? \nz.mem [82] : 
                        (N30)? \nz.mem [125] : 
                        (N32)? \nz.mem [168] : 
                        (N34)? \nz.mem [211] : 
                        (N36)? \nz.mem [254] : 
                        (N38)? \nz.mem [297] : 
                        (N40)? \nz.mem [340] : 
                        (N27)? \nz.mem [383] : 
                        (N29)? \nz.mem [426] : 
                        (N31)? \nz.mem [469] : 
                        (N33)? \nz.mem [512] : 
                        (N35)? \nz.mem [555] : 
                        (N37)? \nz.mem [598] : 
                        (N39)? \nz.mem [641] : 
                        (N41)? \nz.mem [684] : 1'b0;
  assign r_data_o[38] = (N26)? \nz.mem [38] : 
                        (N28)? \nz.mem [81] : 
                        (N30)? \nz.mem [124] : 
                        (N32)? \nz.mem [167] : 
                        (N34)? \nz.mem [210] : 
                        (N36)? \nz.mem [253] : 
                        (N38)? \nz.mem [296] : 
                        (N40)? \nz.mem [339] : 
                        (N27)? \nz.mem [382] : 
                        (N29)? \nz.mem [425] : 
                        (N31)? \nz.mem [468] : 
                        (N33)? \nz.mem [511] : 
                        (N35)? \nz.mem [554] : 
                        (N37)? \nz.mem [597] : 
                        (N39)? \nz.mem [640] : 
                        (N41)? \nz.mem [683] : 1'b0;
  assign r_data_o[37] = (N26)? \nz.mem [37] : 
                        (N28)? \nz.mem [80] : 
                        (N30)? \nz.mem [123] : 
                        (N32)? \nz.mem [166] : 
                        (N34)? \nz.mem [209] : 
                        (N36)? \nz.mem [252] : 
                        (N38)? \nz.mem [295] : 
                        (N40)? \nz.mem [338] : 
                        (N27)? \nz.mem [381] : 
                        (N29)? \nz.mem [424] : 
                        (N31)? \nz.mem [467] : 
                        (N33)? \nz.mem [510] : 
                        (N35)? \nz.mem [553] : 
                        (N37)? \nz.mem [596] : 
                        (N39)? \nz.mem [639] : 
                        (N41)? \nz.mem [682] : 1'b0;
  assign r_data_o[36] = (N26)? \nz.mem [36] : 
                        (N28)? \nz.mem [79] : 
                        (N30)? \nz.mem [122] : 
                        (N32)? \nz.mem [165] : 
                        (N34)? \nz.mem [208] : 
                        (N36)? \nz.mem [251] : 
                        (N38)? \nz.mem [294] : 
                        (N40)? \nz.mem [337] : 
                        (N27)? \nz.mem [380] : 
                        (N29)? \nz.mem [423] : 
                        (N31)? \nz.mem [466] : 
                        (N33)? \nz.mem [509] : 
                        (N35)? \nz.mem [552] : 
                        (N37)? \nz.mem [595] : 
                        (N39)? \nz.mem [638] : 
                        (N41)? \nz.mem [681] : 1'b0;
  assign r_data_o[35] = (N26)? \nz.mem [35] : 
                        (N28)? \nz.mem [78] : 
                        (N30)? \nz.mem [121] : 
                        (N32)? \nz.mem [164] : 
                        (N34)? \nz.mem [207] : 
                        (N36)? \nz.mem [250] : 
                        (N38)? \nz.mem [293] : 
                        (N40)? \nz.mem [336] : 
                        (N27)? \nz.mem [379] : 
                        (N29)? \nz.mem [422] : 
                        (N31)? \nz.mem [465] : 
                        (N33)? \nz.mem [508] : 
                        (N35)? \nz.mem [551] : 
                        (N37)? \nz.mem [594] : 
                        (N39)? \nz.mem [637] : 
                        (N41)? \nz.mem [680] : 1'b0;
  assign r_data_o[34] = (N26)? \nz.mem [34] : 
                        (N28)? \nz.mem [77] : 
                        (N30)? \nz.mem [120] : 
                        (N32)? \nz.mem [163] : 
                        (N34)? \nz.mem [206] : 
                        (N36)? \nz.mem [249] : 
                        (N38)? \nz.mem [292] : 
                        (N40)? \nz.mem [335] : 
                        (N27)? \nz.mem [378] : 
                        (N29)? \nz.mem [421] : 
                        (N31)? \nz.mem [464] : 
                        (N33)? \nz.mem [507] : 
                        (N35)? \nz.mem [550] : 
                        (N37)? \nz.mem [593] : 
                        (N39)? \nz.mem [636] : 
                        (N41)? \nz.mem [679] : 1'b0;
  assign r_data_o[33] = (N26)? \nz.mem [33] : 
                        (N28)? \nz.mem [76] : 
                        (N30)? \nz.mem [119] : 
                        (N32)? \nz.mem [162] : 
                        (N34)? \nz.mem [205] : 
                        (N36)? \nz.mem [248] : 
                        (N38)? \nz.mem [291] : 
                        (N40)? \nz.mem [334] : 
                        (N27)? \nz.mem [377] : 
                        (N29)? \nz.mem [420] : 
                        (N31)? \nz.mem [463] : 
                        (N33)? \nz.mem [506] : 
                        (N35)? \nz.mem [549] : 
                        (N37)? \nz.mem [592] : 
                        (N39)? \nz.mem [635] : 
                        (N41)? \nz.mem [678] : 1'b0;
  assign r_data_o[32] = (N26)? \nz.mem [32] : 
                        (N28)? \nz.mem [75] : 
                        (N30)? \nz.mem [118] : 
                        (N32)? \nz.mem [161] : 
                        (N34)? \nz.mem [204] : 
                        (N36)? \nz.mem [247] : 
                        (N38)? \nz.mem [290] : 
                        (N40)? \nz.mem [333] : 
                        (N27)? \nz.mem [376] : 
                        (N29)? \nz.mem [419] : 
                        (N31)? \nz.mem [462] : 
                        (N33)? \nz.mem [505] : 
                        (N35)? \nz.mem [548] : 
                        (N37)? \nz.mem [591] : 
                        (N39)? \nz.mem [634] : 
                        (N41)? \nz.mem [677] : 1'b0;
  assign r_data_o[31] = (N26)? \nz.mem [31] : 
                        (N28)? \nz.mem [74] : 
                        (N30)? \nz.mem [117] : 
                        (N32)? \nz.mem [160] : 
                        (N34)? \nz.mem [203] : 
                        (N36)? \nz.mem [246] : 
                        (N38)? \nz.mem [289] : 
                        (N40)? \nz.mem [332] : 
                        (N27)? \nz.mem [375] : 
                        (N29)? \nz.mem [418] : 
                        (N31)? \nz.mem [461] : 
                        (N33)? \nz.mem [504] : 
                        (N35)? \nz.mem [547] : 
                        (N37)? \nz.mem [590] : 
                        (N39)? \nz.mem [633] : 
                        (N41)? \nz.mem [676] : 1'b0;
  assign r_data_o[30] = (N26)? \nz.mem [30] : 
                        (N28)? \nz.mem [73] : 
                        (N30)? \nz.mem [116] : 
                        (N32)? \nz.mem [159] : 
                        (N34)? \nz.mem [202] : 
                        (N36)? \nz.mem [245] : 
                        (N38)? \nz.mem [288] : 
                        (N40)? \nz.mem [331] : 
                        (N27)? \nz.mem [374] : 
                        (N29)? \nz.mem [417] : 
                        (N31)? \nz.mem [460] : 
                        (N33)? \nz.mem [503] : 
                        (N35)? \nz.mem [546] : 
                        (N37)? \nz.mem [589] : 
                        (N39)? \nz.mem [632] : 
                        (N41)? \nz.mem [675] : 1'b0;
  assign r_data_o[29] = (N26)? \nz.mem [29] : 
                        (N28)? \nz.mem [72] : 
                        (N30)? \nz.mem [115] : 
                        (N32)? \nz.mem [158] : 
                        (N34)? \nz.mem [201] : 
                        (N36)? \nz.mem [244] : 
                        (N38)? \nz.mem [287] : 
                        (N40)? \nz.mem [330] : 
                        (N27)? \nz.mem [373] : 
                        (N29)? \nz.mem [416] : 
                        (N31)? \nz.mem [459] : 
                        (N33)? \nz.mem [502] : 
                        (N35)? \nz.mem [545] : 
                        (N37)? \nz.mem [588] : 
                        (N39)? \nz.mem [631] : 
                        (N41)? \nz.mem [674] : 1'b0;
  assign r_data_o[28] = (N26)? \nz.mem [28] : 
                        (N28)? \nz.mem [71] : 
                        (N30)? \nz.mem [114] : 
                        (N32)? \nz.mem [157] : 
                        (N34)? \nz.mem [200] : 
                        (N36)? \nz.mem [243] : 
                        (N38)? \nz.mem [286] : 
                        (N40)? \nz.mem [329] : 
                        (N27)? \nz.mem [372] : 
                        (N29)? \nz.mem [415] : 
                        (N31)? \nz.mem [458] : 
                        (N33)? \nz.mem [501] : 
                        (N35)? \nz.mem [544] : 
                        (N37)? \nz.mem [587] : 
                        (N39)? \nz.mem [630] : 
                        (N41)? \nz.mem [673] : 1'b0;
  assign r_data_o[27] = (N26)? \nz.mem [27] : 
                        (N28)? \nz.mem [70] : 
                        (N30)? \nz.mem [113] : 
                        (N32)? \nz.mem [156] : 
                        (N34)? \nz.mem [199] : 
                        (N36)? \nz.mem [242] : 
                        (N38)? \nz.mem [285] : 
                        (N40)? \nz.mem [328] : 
                        (N27)? \nz.mem [371] : 
                        (N29)? \nz.mem [414] : 
                        (N31)? \nz.mem [457] : 
                        (N33)? \nz.mem [500] : 
                        (N35)? \nz.mem [543] : 
                        (N37)? \nz.mem [586] : 
                        (N39)? \nz.mem [629] : 
                        (N41)? \nz.mem [672] : 1'b0;
  assign r_data_o[26] = (N26)? \nz.mem [26] : 
                        (N28)? \nz.mem [69] : 
                        (N30)? \nz.mem [112] : 
                        (N32)? \nz.mem [155] : 
                        (N34)? \nz.mem [198] : 
                        (N36)? \nz.mem [241] : 
                        (N38)? \nz.mem [284] : 
                        (N40)? \nz.mem [327] : 
                        (N27)? \nz.mem [370] : 
                        (N29)? \nz.mem [413] : 
                        (N31)? \nz.mem [456] : 
                        (N33)? \nz.mem [499] : 
                        (N35)? \nz.mem [542] : 
                        (N37)? \nz.mem [585] : 
                        (N39)? \nz.mem [628] : 
                        (N41)? \nz.mem [671] : 1'b0;
  assign r_data_o[25] = (N26)? \nz.mem [25] : 
                        (N28)? \nz.mem [68] : 
                        (N30)? \nz.mem [111] : 
                        (N32)? \nz.mem [154] : 
                        (N34)? \nz.mem [197] : 
                        (N36)? \nz.mem [240] : 
                        (N38)? \nz.mem [283] : 
                        (N40)? \nz.mem [326] : 
                        (N27)? \nz.mem [369] : 
                        (N29)? \nz.mem [412] : 
                        (N31)? \nz.mem [455] : 
                        (N33)? \nz.mem [498] : 
                        (N35)? \nz.mem [541] : 
                        (N37)? \nz.mem [584] : 
                        (N39)? \nz.mem [627] : 
                        (N41)? \nz.mem [670] : 1'b0;
  assign r_data_o[24] = (N26)? \nz.mem [24] : 
                        (N28)? \nz.mem [67] : 
                        (N30)? \nz.mem [110] : 
                        (N32)? \nz.mem [153] : 
                        (N34)? \nz.mem [196] : 
                        (N36)? \nz.mem [239] : 
                        (N38)? \nz.mem [282] : 
                        (N40)? \nz.mem [325] : 
                        (N27)? \nz.mem [368] : 
                        (N29)? \nz.mem [411] : 
                        (N31)? \nz.mem [454] : 
                        (N33)? \nz.mem [497] : 
                        (N35)? \nz.mem [540] : 
                        (N37)? \nz.mem [583] : 
                        (N39)? \nz.mem [626] : 
                        (N41)? \nz.mem [669] : 1'b0;
  assign r_data_o[23] = (N26)? \nz.mem [23] : 
                        (N28)? \nz.mem [66] : 
                        (N30)? \nz.mem [109] : 
                        (N32)? \nz.mem [152] : 
                        (N34)? \nz.mem [195] : 
                        (N36)? \nz.mem [238] : 
                        (N38)? \nz.mem [281] : 
                        (N40)? \nz.mem [324] : 
                        (N27)? \nz.mem [367] : 
                        (N29)? \nz.mem [410] : 
                        (N31)? \nz.mem [453] : 
                        (N33)? \nz.mem [496] : 
                        (N35)? \nz.mem [539] : 
                        (N37)? \nz.mem [582] : 
                        (N39)? \nz.mem [625] : 
                        (N41)? \nz.mem [668] : 1'b0;
  assign r_data_o[22] = (N26)? \nz.mem [22] : 
                        (N28)? \nz.mem [65] : 
                        (N30)? \nz.mem [108] : 
                        (N32)? \nz.mem [151] : 
                        (N34)? \nz.mem [194] : 
                        (N36)? \nz.mem [237] : 
                        (N38)? \nz.mem [280] : 
                        (N40)? \nz.mem [323] : 
                        (N27)? \nz.mem [366] : 
                        (N29)? \nz.mem [409] : 
                        (N31)? \nz.mem [452] : 
                        (N33)? \nz.mem [495] : 
                        (N35)? \nz.mem [538] : 
                        (N37)? \nz.mem [581] : 
                        (N39)? \nz.mem [624] : 
                        (N41)? \nz.mem [667] : 1'b0;
  assign r_data_o[21] = (N26)? \nz.mem [21] : 
                        (N28)? \nz.mem [64] : 
                        (N30)? \nz.mem [107] : 
                        (N32)? \nz.mem [150] : 
                        (N34)? \nz.mem [193] : 
                        (N36)? \nz.mem [236] : 
                        (N38)? \nz.mem [279] : 
                        (N40)? \nz.mem [322] : 
                        (N27)? \nz.mem [365] : 
                        (N29)? \nz.mem [408] : 
                        (N31)? \nz.mem [451] : 
                        (N33)? \nz.mem [494] : 
                        (N35)? \nz.mem [537] : 
                        (N37)? \nz.mem [580] : 
                        (N39)? \nz.mem [623] : 
                        (N41)? \nz.mem [666] : 1'b0;
  assign r_data_o[20] = (N26)? \nz.mem [20] : 
                        (N28)? \nz.mem [63] : 
                        (N30)? \nz.mem [106] : 
                        (N32)? \nz.mem [149] : 
                        (N34)? \nz.mem [192] : 
                        (N36)? \nz.mem [235] : 
                        (N38)? \nz.mem [278] : 
                        (N40)? \nz.mem [321] : 
                        (N27)? \nz.mem [364] : 
                        (N29)? \nz.mem [407] : 
                        (N31)? \nz.mem [450] : 
                        (N33)? \nz.mem [493] : 
                        (N35)? \nz.mem [536] : 
                        (N37)? \nz.mem [579] : 
                        (N39)? \nz.mem [622] : 
                        (N41)? \nz.mem [665] : 1'b0;
  assign r_data_o[19] = (N26)? \nz.mem [19] : 
                        (N28)? \nz.mem [62] : 
                        (N30)? \nz.mem [105] : 
                        (N32)? \nz.mem [148] : 
                        (N34)? \nz.mem [191] : 
                        (N36)? \nz.mem [234] : 
                        (N38)? \nz.mem [277] : 
                        (N40)? \nz.mem [320] : 
                        (N27)? \nz.mem [363] : 
                        (N29)? \nz.mem [406] : 
                        (N31)? \nz.mem [449] : 
                        (N33)? \nz.mem [492] : 
                        (N35)? \nz.mem [535] : 
                        (N37)? \nz.mem [578] : 
                        (N39)? \nz.mem [621] : 
                        (N41)? \nz.mem [664] : 1'b0;
  assign r_data_o[18] = (N26)? \nz.mem [18] : 
                        (N28)? \nz.mem [61] : 
                        (N30)? \nz.mem [104] : 
                        (N32)? \nz.mem [147] : 
                        (N34)? \nz.mem [190] : 
                        (N36)? \nz.mem [233] : 
                        (N38)? \nz.mem [276] : 
                        (N40)? \nz.mem [319] : 
                        (N27)? \nz.mem [362] : 
                        (N29)? \nz.mem [405] : 
                        (N31)? \nz.mem [448] : 
                        (N33)? \nz.mem [491] : 
                        (N35)? \nz.mem [534] : 
                        (N37)? \nz.mem [577] : 
                        (N39)? \nz.mem [620] : 
                        (N41)? \nz.mem [663] : 1'b0;
  assign r_data_o[17] = (N26)? \nz.mem [17] : 
                        (N28)? \nz.mem [60] : 
                        (N30)? \nz.mem [103] : 
                        (N32)? \nz.mem [146] : 
                        (N34)? \nz.mem [189] : 
                        (N36)? \nz.mem [232] : 
                        (N38)? \nz.mem [275] : 
                        (N40)? \nz.mem [318] : 
                        (N27)? \nz.mem [361] : 
                        (N29)? \nz.mem [404] : 
                        (N31)? \nz.mem [447] : 
                        (N33)? \nz.mem [490] : 
                        (N35)? \nz.mem [533] : 
                        (N37)? \nz.mem [576] : 
                        (N39)? \nz.mem [619] : 
                        (N41)? \nz.mem [662] : 1'b0;
  assign r_data_o[16] = (N26)? \nz.mem [16] : 
                        (N28)? \nz.mem [59] : 
                        (N30)? \nz.mem [102] : 
                        (N32)? \nz.mem [145] : 
                        (N34)? \nz.mem [188] : 
                        (N36)? \nz.mem [231] : 
                        (N38)? \nz.mem [274] : 
                        (N40)? \nz.mem [317] : 
                        (N27)? \nz.mem [360] : 
                        (N29)? \nz.mem [403] : 
                        (N31)? \nz.mem [446] : 
                        (N33)? \nz.mem [489] : 
                        (N35)? \nz.mem [532] : 
                        (N37)? \nz.mem [575] : 
                        (N39)? \nz.mem [618] : 
                        (N41)? \nz.mem [661] : 1'b0;
  assign r_data_o[15] = (N26)? \nz.mem [15] : 
                        (N28)? \nz.mem [58] : 
                        (N30)? \nz.mem [101] : 
                        (N32)? \nz.mem [144] : 
                        (N34)? \nz.mem [187] : 
                        (N36)? \nz.mem [230] : 
                        (N38)? \nz.mem [273] : 
                        (N40)? \nz.mem [316] : 
                        (N27)? \nz.mem [359] : 
                        (N29)? \nz.mem [402] : 
                        (N31)? \nz.mem [445] : 
                        (N33)? \nz.mem [488] : 
                        (N35)? \nz.mem [531] : 
                        (N37)? \nz.mem [574] : 
                        (N39)? \nz.mem [617] : 
                        (N41)? \nz.mem [660] : 1'b0;
  assign r_data_o[14] = (N26)? \nz.mem [14] : 
                        (N28)? \nz.mem [57] : 
                        (N30)? \nz.mem [100] : 
                        (N32)? \nz.mem [143] : 
                        (N34)? \nz.mem [186] : 
                        (N36)? \nz.mem [229] : 
                        (N38)? \nz.mem [272] : 
                        (N40)? \nz.mem [315] : 
                        (N27)? \nz.mem [358] : 
                        (N29)? \nz.mem [401] : 
                        (N31)? \nz.mem [444] : 
                        (N33)? \nz.mem [487] : 
                        (N35)? \nz.mem [530] : 
                        (N37)? \nz.mem [573] : 
                        (N39)? \nz.mem [616] : 
                        (N41)? \nz.mem [659] : 1'b0;
  assign r_data_o[13] = (N26)? \nz.mem [13] : 
                        (N28)? \nz.mem [56] : 
                        (N30)? \nz.mem [99] : 
                        (N32)? \nz.mem [142] : 
                        (N34)? \nz.mem [185] : 
                        (N36)? \nz.mem [228] : 
                        (N38)? \nz.mem [271] : 
                        (N40)? \nz.mem [314] : 
                        (N27)? \nz.mem [357] : 
                        (N29)? \nz.mem [400] : 
                        (N31)? \nz.mem [443] : 
                        (N33)? \nz.mem [486] : 
                        (N35)? \nz.mem [529] : 
                        (N37)? \nz.mem [572] : 
                        (N39)? \nz.mem [615] : 
                        (N41)? \nz.mem [658] : 1'b0;
  assign r_data_o[12] = (N26)? \nz.mem [12] : 
                        (N28)? \nz.mem [55] : 
                        (N30)? \nz.mem [98] : 
                        (N32)? \nz.mem [141] : 
                        (N34)? \nz.mem [184] : 
                        (N36)? \nz.mem [227] : 
                        (N38)? \nz.mem [270] : 
                        (N40)? \nz.mem [313] : 
                        (N27)? \nz.mem [356] : 
                        (N29)? \nz.mem [399] : 
                        (N31)? \nz.mem [442] : 
                        (N33)? \nz.mem [485] : 
                        (N35)? \nz.mem [528] : 
                        (N37)? \nz.mem [571] : 
                        (N39)? \nz.mem [614] : 
                        (N41)? \nz.mem [657] : 1'b0;
  assign r_data_o[11] = (N26)? \nz.mem [11] : 
                        (N28)? \nz.mem [54] : 
                        (N30)? \nz.mem [97] : 
                        (N32)? \nz.mem [140] : 
                        (N34)? \nz.mem [183] : 
                        (N36)? \nz.mem [226] : 
                        (N38)? \nz.mem [269] : 
                        (N40)? \nz.mem [312] : 
                        (N27)? \nz.mem [355] : 
                        (N29)? \nz.mem [398] : 
                        (N31)? \nz.mem [441] : 
                        (N33)? \nz.mem [484] : 
                        (N35)? \nz.mem [527] : 
                        (N37)? \nz.mem [570] : 
                        (N39)? \nz.mem [613] : 
                        (N41)? \nz.mem [656] : 1'b0;
  assign r_data_o[10] = (N26)? \nz.mem [10] : 
                        (N28)? \nz.mem [53] : 
                        (N30)? \nz.mem [96] : 
                        (N32)? \nz.mem [139] : 
                        (N34)? \nz.mem [182] : 
                        (N36)? \nz.mem [225] : 
                        (N38)? \nz.mem [268] : 
                        (N40)? \nz.mem [311] : 
                        (N27)? \nz.mem [354] : 
                        (N29)? \nz.mem [397] : 
                        (N31)? \nz.mem [440] : 
                        (N33)? \nz.mem [483] : 
                        (N35)? \nz.mem [526] : 
                        (N37)? \nz.mem [569] : 
                        (N39)? \nz.mem [612] : 
                        (N41)? \nz.mem [655] : 1'b0;
  assign r_data_o[9] = (N26)? \nz.mem [9] : 
                       (N28)? \nz.mem [52] : 
                       (N30)? \nz.mem [95] : 
                       (N32)? \nz.mem [138] : 
                       (N34)? \nz.mem [181] : 
                       (N36)? \nz.mem [224] : 
                       (N38)? \nz.mem [267] : 
                       (N40)? \nz.mem [310] : 
                       (N27)? \nz.mem [353] : 
                       (N29)? \nz.mem [396] : 
                       (N31)? \nz.mem [439] : 
                       (N33)? \nz.mem [482] : 
                       (N35)? \nz.mem [525] : 
                       (N37)? \nz.mem [568] : 
                       (N39)? \nz.mem [611] : 
                       (N41)? \nz.mem [654] : 1'b0;
  assign r_data_o[8] = (N26)? \nz.mem [8] : 
                       (N28)? \nz.mem [51] : 
                       (N30)? \nz.mem [94] : 
                       (N32)? \nz.mem [137] : 
                       (N34)? \nz.mem [180] : 
                       (N36)? \nz.mem [223] : 
                       (N38)? \nz.mem [266] : 
                       (N40)? \nz.mem [309] : 
                       (N27)? \nz.mem [352] : 
                       (N29)? \nz.mem [395] : 
                       (N31)? \nz.mem [438] : 
                       (N33)? \nz.mem [481] : 
                       (N35)? \nz.mem [524] : 
                       (N37)? \nz.mem [567] : 
                       (N39)? \nz.mem [610] : 
                       (N41)? \nz.mem [653] : 1'b0;
  assign r_data_o[7] = (N26)? \nz.mem [7] : 
                       (N28)? \nz.mem [50] : 
                       (N30)? \nz.mem [93] : 
                       (N32)? \nz.mem [136] : 
                       (N34)? \nz.mem [179] : 
                       (N36)? \nz.mem [222] : 
                       (N38)? \nz.mem [265] : 
                       (N40)? \nz.mem [308] : 
                       (N27)? \nz.mem [351] : 
                       (N29)? \nz.mem [394] : 
                       (N31)? \nz.mem [437] : 
                       (N33)? \nz.mem [480] : 
                       (N35)? \nz.mem [523] : 
                       (N37)? \nz.mem [566] : 
                       (N39)? \nz.mem [609] : 
                       (N41)? \nz.mem [652] : 1'b0;
  assign r_data_o[6] = (N26)? \nz.mem [6] : 
                       (N28)? \nz.mem [49] : 
                       (N30)? \nz.mem [92] : 
                       (N32)? \nz.mem [135] : 
                       (N34)? \nz.mem [178] : 
                       (N36)? \nz.mem [221] : 
                       (N38)? \nz.mem [264] : 
                       (N40)? \nz.mem [307] : 
                       (N27)? \nz.mem [350] : 
                       (N29)? \nz.mem [393] : 
                       (N31)? \nz.mem [436] : 
                       (N33)? \nz.mem [479] : 
                       (N35)? \nz.mem [522] : 
                       (N37)? \nz.mem [565] : 
                       (N39)? \nz.mem [608] : 
                       (N41)? \nz.mem [651] : 1'b0;
  assign r_data_o[5] = (N26)? \nz.mem [5] : 
                       (N28)? \nz.mem [48] : 
                       (N30)? \nz.mem [91] : 
                       (N32)? \nz.mem [134] : 
                       (N34)? \nz.mem [177] : 
                       (N36)? \nz.mem [220] : 
                       (N38)? \nz.mem [263] : 
                       (N40)? \nz.mem [306] : 
                       (N27)? \nz.mem [349] : 
                       (N29)? \nz.mem [392] : 
                       (N31)? \nz.mem [435] : 
                       (N33)? \nz.mem [478] : 
                       (N35)? \nz.mem [521] : 
                       (N37)? \nz.mem [564] : 
                       (N39)? \nz.mem [607] : 
                       (N41)? \nz.mem [650] : 1'b0;
  assign r_data_o[4] = (N26)? \nz.mem [4] : 
                       (N28)? \nz.mem [47] : 
                       (N30)? \nz.mem [90] : 
                       (N32)? \nz.mem [133] : 
                       (N34)? \nz.mem [176] : 
                       (N36)? \nz.mem [219] : 
                       (N38)? \nz.mem [262] : 
                       (N40)? \nz.mem [305] : 
                       (N27)? \nz.mem [348] : 
                       (N29)? \nz.mem [391] : 
                       (N31)? \nz.mem [434] : 
                       (N33)? \nz.mem [477] : 
                       (N35)? \nz.mem [520] : 
                       (N37)? \nz.mem [563] : 
                       (N39)? \nz.mem [606] : 
                       (N41)? \nz.mem [649] : 1'b0;
  assign r_data_o[3] = (N26)? \nz.mem [3] : 
                       (N28)? \nz.mem [46] : 
                       (N30)? \nz.mem [89] : 
                       (N32)? \nz.mem [132] : 
                       (N34)? \nz.mem [175] : 
                       (N36)? \nz.mem [218] : 
                       (N38)? \nz.mem [261] : 
                       (N40)? \nz.mem [304] : 
                       (N27)? \nz.mem [347] : 
                       (N29)? \nz.mem [390] : 
                       (N31)? \nz.mem [433] : 
                       (N33)? \nz.mem [476] : 
                       (N35)? \nz.mem [519] : 
                       (N37)? \nz.mem [562] : 
                       (N39)? \nz.mem [605] : 
                       (N41)? \nz.mem [648] : 1'b0;
  assign r_data_o[2] = (N26)? \nz.mem [2] : 
                       (N28)? \nz.mem [45] : 
                       (N30)? \nz.mem [88] : 
                       (N32)? \nz.mem [131] : 
                       (N34)? \nz.mem [174] : 
                       (N36)? \nz.mem [217] : 
                       (N38)? \nz.mem [260] : 
                       (N40)? \nz.mem [303] : 
                       (N27)? \nz.mem [346] : 
                       (N29)? \nz.mem [389] : 
                       (N31)? \nz.mem [432] : 
                       (N33)? \nz.mem [475] : 
                       (N35)? \nz.mem [518] : 
                       (N37)? \nz.mem [561] : 
                       (N39)? \nz.mem [604] : 
                       (N41)? \nz.mem [647] : 1'b0;
  assign r_data_o[1] = (N26)? \nz.mem [1] : 
                       (N28)? \nz.mem [44] : 
                       (N30)? \nz.mem [87] : 
                       (N32)? \nz.mem [130] : 
                       (N34)? \nz.mem [173] : 
                       (N36)? \nz.mem [216] : 
                       (N38)? \nz.mem [259] : 
                       (N40)? \nz.mem [302] : 
                       (N27)? \nz.mem [345] : 
                       (N29)? \nz.mem [388] : 
                       (N31)? \nz.mem [431] : 
                       (N33)? \nz.mem [474] : 
                       (N35)? \nz.mem [517] : 
                       (N37)? \nz.mem [560] : 
                       (N39)? \nz.mem [603] : 
                       (N41)? \nz.mem [646] : 1'b0;
  assign r_data_o[0] = (N26)? \nz.mem [0] : 
                       (N28)? \nz.mem [43] : 
                       (N30)? \nz.mem [86] : 
                       (N32)? \nz.mem [129] : 
                       (N34)? \nz.mem [172] : 
                       (N36)? \nz.mem [215] : 
                       (N38)? \nz.mem [258] : 
                       (N40)? \nz.mem [301] : 
                       (N27)? \nz.mem [344] : 
                       (N29)? \nz.mem [387] : 
                       (N31)? \nz.mem [430] : 
                       (N33)? \nz.mem [473] : 
                       (N35)? \nz.mem [516] : 
                       (N37)? \nz.mem [559] : 
                       (N39)? \nz.mem [602] : 
                       (N41)? \nz.mem [645] : 1'b0;
  assign N75 = w_addr_i[2] & w_addr_i[3];
  assign N76 = N0 & w_addr_i[3];
  assign N0 = ~w_addr_i[2];
  assign N77 = w_addr_i[2] & N1;
  assign N1 = ~w_addr_i[3];
  assign N78 = N2 & N3;
  assign N2 = ~w_addr_i[2];
  assign N3 = ~w_addr_i[3];
  assign N79 = w_addr_i[0] & w_addr_i[1];
  assign N80 = N4 & w_addr_i[1];
  assign N4 = ~w_addr_i[0];
  assign N81 = w_addr_i[0] & N5;
  assign N5 = ~w_addr_i[1];
  assign N82 = N6 & N7;
  assign N6 = ~w_addr_i[0];
  assign N7 = ~w_addr_i[1];
  assign N58 = N75 & N79;
  assign N57 = N75 & N80;
  assign N56 = N75 & N81;
  assign N55 = N75 & N82;
  assign N54 = N76 & N79;
  assign N53 = N76 & N80;
  assign N52 = N76 & N81;
  assign N51 = N76 & N82;
  assign N50 = N77 & N79;
  assign N49 = N77 & N80;
  assign N48 = N77 & N81;
  assign N47 = N77 & N82;
  assign N46 = N78 & N79;
  assign N45 = N78 & N80;
  assign N44 = N78 & N81;
  assign N43 = N78 & N82;
  assign { N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59 } = (N8)? { N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43 } : 
                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N42;
  assign N10 = ~r_addr_i[0];
  assign N11 = ~r_addr_i[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r_addr_i[1];
  assign N14 = r_addr_i[0] & N11;
  assign N15 = r_addr_i[0] & r_addr_i[1];
  assign N16 = ~r_addr_i[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r_addr_i[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r_addr_i[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r_addr_i[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r_addr_i[2];
  assign N25 = ~r_addr_i[3];
  assign N26 = N17 & N25;
  assign N27 = N17 & r_addr_i[3];
  assign N28 = N19 & N25;
  assign N29 = N19 & r_addr_i[3];
  assign N30 = N21 & N25;
  assign N31 = N21 & r_addr_i[3];
  assign N32 = N23 & N25;
  assign N33 = N23 & r_addr_i[3];
  assign N34 = N18 & N25;
  assign N35 = N18 & r_addr_i[3];
  assign N36 = N20 & N25;
  assign N37 = N20 & r_addr_i[3];
  assign N38 = N22 & N25;
  assign N39 = N22 & r_addr_i[3];
  assign N40 = N24 & N25;
  assign N41 = N24 & r_addr_i[3];
  assign N42 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N74) begin
      \nz.mem_687_sv2v_reg  <= w_data_i[42];
      \nz.mem_686_sv2v_reg  <= w_data_i[41];
      \nz.mem_685_sv2v_reg  <= w_data_i[40];
      \nz.mem_684_sv2v_reg  <= w_data_i[39];
      \nz.mem_683_sv2v_reg  <= w_data_i[38];
      \nz.mem_682_sv2v_reg  <= w_data_i[37];
      \nz.mem_681_sv2v_reg  <= w_data_i[36];
      \nz.mem_680_sv2v_reg  <= w_data_i[35];
      \nz.mem_679_sv2v_reg  <= w_data_i[34];
      \nz.mem_678_sv2v_reg  <= w_data_i[33];
      \nz.mem_677_sv2v_reg  <= w_data_i[32];
      \nz.mem_676_sv2v_reg  <= w_data_i[31];
      \nz.mem_675_sv2v_reg  <= w_data_i[30];
      \nz.mem_674_sv2v_reg  <= w_data_i[29];
      \nz.mem_673_sv2v_reg  <= w_data_i[28];
      \nz.mem_672_sv2v_reg  <= w_data_i[27];
      \nz.mem_671_sv2v_reg  <= w_data_i[26];
      \nz.mem_670_sv2v_reg  <= w_data_i[25];
      \nz.mem_669_sv2v_reg  <= w_data_i[24];
      \nz.mem_668_sv2v_reg  <= w_data_i[23];
      \nz.mem_667_sv2v_reg  <= w_data_i[22];
      \nz.mem_666_sv2v_reg  <= w_data_i[21];
      \nz.mem_665_sv2v_reg  <= w_data_i[20];
      \nz.mem_664_sv2v_reg  <= w_data_i[19];
      \nz.mem_663_sv2v_reg  <= w_data_i[18];
      \nz.mem_662_sv2v_reg  <= w_data_i[17];
      \nz.mem_661_sv2v_reg  <= w_data_i[16];
      \nz.mem_660_sv2v_reg  <= w_data_i[15];
      \nz.mem_659_sv2v_reg  <= w_data_i[14];
      \nz.mem_658_sv2v_reg  <= w_data_i[13];
      \nz.mem_657_sv2v_reg  <= w_data_i[12];
      \nz.mem_656_sv2v_reg  <= w_data_i[11];
      \nz.mem_655_sv2v_reg  <= w_data_i[10];
      \nz.mem_654_sv2v_reg  <= w_data_i[9];
      \nz.mem_653_sv2v_reg  <= w_data_i[8];
      \nz.mem_652_sv2v_reg  <= w_data_i[7];
      \nz.mem_651_sv2v_reg  <= w_data_i[6];
      \nz.mem_650_sv2v_reg  <= w_data_i[5];
      \nz.mem_649_sv2v_reg  <= w_data_i[4];
      \nz.mem_648_sv2v_reg  <= w_data_i[3];
      \nz.mem_647_sv2v_reg  <= w_data_i[2];
      \nz.mem_646_sv2v_reg  <= w_data_i[1];
      \nz.mem_645_sv2v_reg  <= w_data_i[0];
    end 
    if(N73) begin
      \nz.mem_644_sv2v_reg  <= w_data_i[42];
      \nz.mem_643_sv2v_reg  <= w_data_i[41];
      \nz.mem_642_sv2v_reg  <= w_data_i[40];
      \nz.mem_641_sv2v_reg  <= w_data_i[39];
      \nz.mem_640_sv2v_reg  <= w_data_i[38];
      \nz.mem_639_sv2v_reg  <= w_data_i[37];
      \nz.mem_638_sv2v_reg  <= w_data_i[36];
      \nz.mem_637_sv2v_reg  <= w_data_i[35];
      \nz.mem_636_sv2v_reg  <= w_data_i[34];
      \nz.mem_635_sv2v_reg  <= w_data_i[33];
      \nz.mem_634_sv2v_reg  <= w_data_i[32];
      \nz.mem_633_sv2v_reg  <= w_data_i[31];
      \nz.mem_632_sv2v_reg  <= w_data_i[30];
      \nz.mem_631_sv2v_reg  <= w_data_i[29];
      \nz.mem_630_sv2v_reg  <= w_data_i[28];
      \nz.mem_629_sv2v_reg  <= w_data_i[27];
      \nz.mem_628_sv2v_reg  <= w_data_i[26];
      \nz.mem_627_sv2v_reg  <= w_data_i[25];
      \nz.mem_626_sv2v_reg  <= w_data_i[24];
      \nz.mem_625_sv2v_reg  <= w_data_i[23];
      \nz.mem_624_sv2v_reg  <= w_data_i[22];
      \nz.mem_623_sv2v_reg  <= w_data_i[21];
      \nz.mem_622_sv2v_reg  <= w_data_i[20];
      \nz.mem_621_sv2v_reg  <= w_data_i[19];
      \nz.mem_620_sv2v_reg  <= w_data_i[18];
      \nz.mem_619_sv2v_reg  <= w_data_i[17];
      \nz.mem_618_sv2v_reg  <= w_data_i[16];
      \nz.mem_617_sv2v_reg  <= w_data_i[15];
      \nz.mem_616_sv2v_reg  <= w_data_i[14];
      \nz.mem_615_sv2v_reg  <= w_data_i[13];
      \nz.mem_614_sv2v_reg  <= w_data_i[12];
      \nz.mem_613_sv2v_reg  <= w_data_i[11];
      \nz.mem_612_sv2v_reg  <= w_data_i[10];
      \nz.mem_611_sv2v_reg  <= w_data_i[9];
      \nz.mem_610_sv2v_reg  <= w_data_i[8];
      \nz.mem_609_sv2v_reg  <= w_data_i[7];
      \nz.mem_608_sv2v_reg  <= w_data_i[6];
      \nz.mem_607_sv2v_reg  <= w_data_i[5];
      \nz.mem_606_sv2v_reg  <= w_data_i[4];
      \nz.mem_605_sv2v_reg  <= w_data_i[3];
      \nz.mem_604_sv2v_reg  <= w_data_i[2];
      \nz.mem_603_sv2v_reg  <= w_data_i[1];
      \nz.mem_602_sv2v_reg  <= w_data_i[0];
    end 
    if(N72) begin
      \nz.mem_601_sv2v_reg  <= w_data_i[42];
      \nz.mem_600_sv2v_reg  <= w_data_i[41];
      \nz.mem_599_sv2v_reg  <= w_data_i[40];
      \nz.mem_598_sv2v_reg  <= w_data_i[39];
      \nz.mem_597_sv2v_reg  <= w_data_i[38];
      \nz.mem_596_sv2v_reg  <= w_data_i[37];
      \nz.mem_595_sv2v_reg  <= w_data_i[36];
      \nz.mem_594_sv2v_reg  <= w_data_i[35];
      \nz.mem_593_sv2v_reg  <= w_data_i[34];
      \nz.mem_592_sv2v_reg  <= w_data_i[33];
      \nz.mem_591_sv2v_reg  <= w_data_i[32];
      \nz.mem_590_sv2v_reg  <= w_data_i[31];
      \nz.mem_589_sv2v_reg  <= w_data_i[30];
      \nz.mem_588_sv2v_reg  <= w_data_i[29];
      \nz.mem_587_sv2v_reg  <= w_data_i[28];
      \nz.mem_586_sv2v_reg  <= w_data_i[27];
      \nz.mem_585_sv2v_reg  <= w_data_i[26];
      \nz.mem_584_sv2v_reg  <= w_data_i[25];
      \nz.mem_583_sv2v_reg  <= w_data_i[24];
      \nz.mem_582_sv2v_reg  <= w_data_i[23];
      \nz.mem_581_sv2v_reg  <= w_data_i[22];
      \nz.mem_580_sv2v_reg  <= w_data_i[21];
      \nz.mem_579_sv2v_reg  <= w_data_i[20];
      \nz.mem_578_sv2v_reg  <= w_data_i[19];
      \nz.mem_577_sv2v_reg  <= w_data_i[18];
      \nz.mem_576_sv2v_reg  <= w_data_i[17];
      \nz.mem_575_sv2v_reg  <= w_data_i[16];
      \nz.mem_574_sv2v_reg  <= w_data_i[15];
      \nz.mem_573_sv2v_reg  <= w_data_i[14];
      \nz.mem_572_sv2v_reg  <= w_data_i[13];
      \nz.mem_571_sv2v_reg  <= w_data_i[12];
      \nz.mem_570_sv2v_reg  <= w_data_i[11];
      \nz.mem_569_sv2v_reg  <= w_data_i[10];
      \nz.mem_568_sv2v_reg  <= w_data_i[9];
      \nz.mem_567_sv2v_reg  <= w_data_i[8];
      \nz.mem_566_sv2v_reg  <= w_data_i[7];
      \nz.mem_565_sv2v_reg  <= w_data_i[6];
      \nz.mem_564_sv2v_reg  <= w_data_i[5];
      \nz.mem_563_sv2v_reg  <= w_data_i[4];
      \nz.mem_562_sv2v_reg  <= w_data_i[3];
      \nz.mem_561_sv2v_reg  <= w_data_i[2];
      \nz.mem_560_sv2v_reg  <= w_data_i[1];
      \nz.mem_559_sv2v_reg  <= w_data_i[0];
    end 
    if(N71) begin
      \nz.mem_558_sv2v_reg  <= w_data_i[42];
      \nz.mem_557_sv2v_reg  <= w_data_i[41];
      \nz.mem_556_sv2v_reg  <= w_data_i[40];
      \nz.mem_555_sv2v_reg  <= w_data_i[39];
      \nz.mem_554_sv2v_reg  <= w_data_i[38];
      \nz.mem_553_sv2v_reg  <= w_data_i[37];
      \nz.mem_552_sv2v_reg  <= w_data_i[36];
      \nz.mem_551_sv2v_reg  <= w_data_i[35];
      \nz.mem_550_sv2v_reg  <= w_data_i[34];
      \nz.mem_549_sv2v_reg  <= w_data_i[33];
      \nz.mem_548_sv2v_reg  <= w_data_i[32];
      \nz.mem_547_sv2v_reg  <= w_data_i[31];
      \nz.mem_546_sv2v_reg  <= w_data_i[30];
      \nz.mem_545_sv2v_reg  <= w_data_i[29];
      \nz.mem_544_sv2v_reg  <= w_data_i[28];
      \nz.mem_543_sv2v_reg  <= w_data_i[27];
      \nz.mem_542_sv2v_reg  <= w_data_i[26];
      \nz.mem_541_sv2v_reg  <= w_data_i[25];
      \nz.mem_540_sv2v_reg  <= w_data_i[24];
      \nz.mem_539_sv2v_reg  <= w_data_i[23];
      \nz.mem_538_sv2v_reg  <= w_data_i[22];
      \nz.mem_537_sv2v_reg  <= w_data_i[21];
      \nz.mem_536_sv2v_reg  <= w_data_i[20];
      \nz.mem_535_sv2v_reg  <= w_data_i[19];
      \nz.mem_534_sv2v_reg  <= w_data_i[18];
      \nz.mem_533_sv2v_reg  <= w_data_i[17];
      \nz.mem_532_sv2v_reg  <= w_data_i[16];
      \nz.mem_531_sv2v_reg  <= w_data_i[15];
      \nz.mem_530_sv2v_reg  <= w_data_i[14];
      \nz.mem_529_sv2v_reg  <= w_data_i[13];
      \nz.mem_528_sv2v_reg  <= w_data_i[12];
      \nz.mem_527_sv2v_reg  <= w_data_i[11];
      \nz.mem_526_sv2v_reg  <= w_data_i[10];
      \nz.mem_525_sv2v_reg  <= w_data_i[9];
      \nz.mem_524_sv2v_reg  <= w_data_i[8];
      \nz.mem_523_sv2v_reg  <= w_data_i[7];
      \nz.mem_522_sv2v_reg  <= w_data_i[6];
      \nz.mem_521_sv2v_reg  <= w_data_i[5];
      \nz.mem_520_sv2v_reg  <= w_data_i[4];
      \nz.mem_519_sv2v_reg  <= w_data_i[3];
      \nz.mem_518_sv2v_reg  <= w_data_i[2];
      \nz.mem_517_sv2v_reg  <= w_data_i[1];
      \nz.mem_516_sv2v_reg  <= w_data_i[0];
    end 
    if(N70) begin
      \nz.mem_515_sv2v_reg  <= w_data_i[42];
      \nz.mem_514_sv2v_reg  <= w_data_i[41];
      \nz.mem_513_sv2v_reg  <= w_data_i[40];
      \nz.mem_512_sv2v_reg  <= w_data_i[39];
      \nz.mem_511_sv2v_reg  <= w_data_i[38];
      \nz.mem_510_sv2v_reg  <= w_data_i[37];
      \nz.mem_509_sv2v_reg  <= w_data_i[36];
      \nz.mem_508_sv2v_reg  <= w_data_i[35];
      \nz.mem_507_sv2v_reg  <= w_data_i[34];
      \nz.mem_506_sv2v_reg  <= w_data_i[33];
      \nz.mem_505_sv2v_reg  <= w_data_i[32];
      \nz.mem_504_sv2v_reg  <= w_data_i[31];
      \nz.mem_503_sv2v_reg  <= w_data_i[30];
      \nz.mem_502_sv2v_reg  <= w_data_i[29];
      \nz.mem_501_sv2v_reg  <= w_data_i[28];
      \nz.mem_500_sv2v_reg  <= w_data_i[27];
      \nz.mem_499_sv2v_reg  <= w_data_i[26];
      \nz.mem_498_sv2v_reg  <= w_data_i[25];
      \nz.mem_497_sv2v_reg  <= w_data_i[24];
      \nz.mem_496_sv2v_reg  <= w_data_i[23];
      \nz.mem_495_sv2v_reg  <= w_data_i[22];
      \nz.mem_494_sv2v_reg  <= w_data_i[21];
      \nz.mem_493_sv2v_reg  <= w_data_i[20];
      \nz.mem_492_sv2v_reg  <= w_data_i[19];
      \nz.mem_491_sv2v_reg  <= w_data_i[18];
      \nz.mem_490_sv2v_reg  <= w_data_i[17];
      \nz.mem_489_sv2v_reg  <= w_data_i[16];
      \nz.mem_488_sv2v_reg  <= w_data_i[15];
      \nz.mem_487_sv2v_reg  <= w_data_i[14];
      \nz.mem_486_sv2v_reg  <= w_data_i[13];
      \nz.mem_485_sv2v_reg  <= w_data_i[12];
      \nz.mem_484_sv2v_reg  <= w_data_i[11];
      \nz.mem_483_sv2v_reg  <= w_data_i[10];
      \nz.mem_482_sv2v_reg  <= w_data_i[9];
      \nz.mem_481_sv2v_reg  <= w_data_i[8];
      \nz.mem_480_sv2v_reg  <= w_data_i[7];
      \nz.mem_479_sv2v_reg  <= w_data_i[6];
      \nz.mem_478_sv2v_reg  <= w_data_i[5];
      \nz.mem_477_sv2v_reg  <= w_data_i[4];
      \nz.mem_476_sv2v_reg  <= w_data_i[3];
      \nz.mem_475_sv2v_reg  <= w_data_i[2];
      \nz.mem_474_sv2v_reg  <= w_data_i[1];
      \nz.mem_473_sv2v_reg  <= w_data_i[0];
    end 
    if(N69) begin
      \nz.mem_472_sv2v_reg  <= w_data_i[42];
      \nz.mem_471_sv2v_reg  <= w_data_i[41];
      \nz.mem_470_sv2v_reg  <= w_data_i[40];
      \nz.mem_469_sv2v_reg  <= w_data_i[39];
      \nz.mem_468_sv2v_reg  <= w_data_i[38];
      \nz.mem_467_sv2v_reg  <= w_data_i[37];
      \nz.mem_466_sv2v_reg  <= w_data_i[36];
      \nz.mem_465_sv2v_reg  <= w_data_i[35];
      \nz.mem_464_sv2v_reg  <= w_data_i[34];
      \nz.mem_463_sv2v_reg  <= w_data_i[33];
      \nz.mem_462_sv2v_reg  <= w_data_i[32];
      \nz.mem_461_sv2v_reg  <= w_data_i[31];
      \nz.mem_460_sv2v_reg  <= w_data_i[30];
      \nz.mem_459_sv2v_reg  <= w_data_i[29];
      \nz.mem_458_sv2v_reg  <= w_data_i[28];
      \nz.mem_457_sv2v_reg  <= w_data_i[27];
      \nz.mem_456_sv2v_reg  <= w_data_i[26];
      \nz.mem_455_sv2v_reg  <= w_data_i[25];
      \nz.mem_454_sv2v_reg  <= w_data_i[24];
      \nz.mem_453_sv2v_reg  <= w_data_i[23];
      \nz.mem_452_sv2v_reg  <= w_data_i[22];
      \nz.mem_451_sv2v_reg  <= w_data_i[21];
      \nz.mem_450_sv2v_reg  <= w_data_i[20];
      \nz.mem_449_sv2v_reg  <= w_data_i[19];
      \nz.mem_448_sv2v_reg  <= w_data_i[18];
      \nz.mem_447_sv2v_reg  <= w_data_i[17];
      \nz.mem_446_sv2v_reg  <= w_data_i[16];
      \nz.mem_445_sv2v_reg  <= w_data_i[15];
      \nz.mem_444_sv2v_reg  <= w_data_i[14];
      \nz.mem_443_sv2v_reg  <= w_data_i[13];
      \nz.mem_442_sv2v_reg  <= w_data_i[12];
      \nz.mem_441_sv2v_reg  <= w_data_i[11];
      \nz.mem_440_sv2v_reg  <= w_data_i[10];
      \nz.mem_439_sv2v_reg  <= w_data_i[9];
      \nz.mem_438_sv2v_reg  <= w_data_i[8];
      \nz.mem_437_sv2v_reg  <= w_data_i[7];
      \nz.mem_436_sv2v_reg  <= w_data_i[6];
      \nz.mem_435_sv2v_reg  <= w_data_i[5];
      \nz.mem_434_sv2v_reg  <= w_data_i[4];
      \nz.mem_433_sv2v_reg  <= w_data_i[3];
      \nz.mem_432_sv2v_reg  <= w_data_i[2];
      \nz.mem_431_sv2v_reg  <= w_data_i[1];
      \nz.mem_430_sv2v_reg  <= w_data_i[0];
    end 
    if(N68) begin
      \nz.mem_429_sv2v_reg  <= w_data_i[42];
      \nz.mem_428_sv2v_reg  <= w_data_i[41];
      \nz.mem_427_sv2v_reg  <= w_data_i[40];
      \nz.mem_426_sv2v_reg  <= w_data_i[39];
      \nz.mem_425_sv2v_reg  <= w_data_i[38];
      \nz.mem_424_sv2v_reg  <= w_data_i[37];
      \nz.mem_423_sv2v_reg  <= w_data_i[36];
      \nz.mem_422_sv2v_reg  <= w_data_i[35];
      \nz.mem_421_sv2v_reg  <= w_data_i[34];
      \nz.mem_420_sv2v_reg  <= w_data_i[33];
      \nz.mem_419_sv2v_reg  <= w_data_i[32];
      \nz.mem_418_sv2v_reg  <= w_data_i[31];
      \nz.mem_417_sv2v_reg  <= w_data_i[30];
      \nz.mem_416_sv2v_reg  <= w_data_i[29];
      \nz.mem_415_sv2v_reg  <= w_data_i[28];
      \nz.mem_414_sv2v_reg  <= w_data_i[27];
      \nz.mem_413_sv2v_reg  <= w_data_i[26];
      \nz.mem_412_sv2v_reg  <= w_data_i[25];
      \nz.mem_411_sv2v_reg  <= w_data_i[24];
      \nz.mem_410_sv2v_reg  <= w_data_i[23];
      \nz.mem_409_sv2v_reg  <= w_data_i[22];
      \nz.mem_408_sv2v_reg  <= w_data_i[21];
      \nz.mem_407_sv2v_reg  <= w_data_i[20];
      \nz.mem_406_sv2v_reg  <= w_data_i[19];
      \nz.mem_405_sv2v_reg  <= w_data_i[18];
      \nz.mem_404_sv2v_reg  <= w_data_i[17];
      \nz.mem_403_sv2v_reg  <= w_data_i[16];
      \nz.mem_402_sv2v_reg  <= w_data_i[15];
      \nz.mem_401_sv2v_reg  <= w_data_i[14];
      \nz.mem_400_sv2v_reg  <= w_data_i[13];
      \nz.mem_399_sv2v_reg  <= w_data_i[12];
      \nz.mem_398_sv2v_reg  <= w_data_i[11];
      \nz.mem_397_sv2v_reg  <= w_data_i[10];
      \nz.mem_396_sv2v_reg  <= w_data_i[9];
      \nz.mem_395_sv2v_reg  <= w_data_i[8];
      \nz.mem_394_sv2v_reg  <= w_data_i[7];
      \nz.mem_393_sv2v_reg  <= w_data_i[6];
      \nz.mem_392_sv2v_reg  <= w_data_i[5];
      \nz.mem_391_sv2v_reg  <= w_data_i[4];
      \nz.mem_390_sv2v_reg  <= w_data_i[3];
      \nz.mem_389_sv2v_reg  <= w_data_i[2];
      \nz.mem_388_sv2v_reg  <= w_data_i[1];
      \nz.mem_387_sv2v_reg  <= w_data_i[0];
    end 
    if(N67) begin
      \nz.mem_386_sv2v_reg  <= w_data_i[42];
      \nz.mem_385_sv2v_reg  <= w_data_i[41];
      \nz.mem_384_sv2v_reg  <= w_data_i[40];
      \nz.mem_383_sv2v_reg  <= w_data_i[39];
      \nz.mem_382_sv2v_reg  <= w_data_i[38];
      \nz.mem_381_sv2v_reg  <= w_data_i[37];
      \nz.mem_380_sv2v_reg  <= w_data_i[36];
      \nz.mem_379_sv2v_reg  <= w_data_i[35];
      \nz.mem_378_sv2v_reg  <= w_data_i[34];
      \nz.mem_377_sv2v_reg  <= w_data_i[33];
      \nz.mem_376_sv2v_reg  <= w_data_i[32];
      \nz.mem_375_sv2v_reg  <= w_data_i[31];
      \nz.mem_374_sv2v_reg  <= w_data_i[30];
      \nz.mem_373_sv2v_reg  <= w_data_i[29];
      \nz.mem_372_sv2v_reg  <= w_data_i[28];
      \nz.mem_371_sv2v_reg  <= w_data_i[27];
      \nz.mem_370_sv2v_reg  <= w_data_i[26];
      \nz.mem_369_sv2v_reg  <= w_data_i[25];
      \nz.mem_368_sv2v_reg  <= w_data_i[24];
      \nz.mem_367_sv2v_reg  <= w_data_i[23];
      \nz.mem_366_sv2v_reg  <= w_data_i[22];
      \nz.mem_365_sv2v_reg  <= w_data_i[21];
      \nz.mem_364_sv2v_reg  <= w_data_i[20];
      \nz.mem_363_sv2v_reg  <= w_data_i[19];
      \nz.mem_362_sv2v_reg  <= w_data_i[18];
      \nz.mem_361_sv2v_reg  <= w_data_i[17];
      \nz.mem_360_sv2v_reg  <= w_data_i[16];
      \nz.mem_359_sv2v_reg  <= w_data_i[15];
      \nz.mem_358_sv2v_reg  <= w_data_i[14];
      \nz.mem_357_sv2v_reg  <= w_data_i[13];
      \nz.mem_356_sv2v_reg  <= w_data_i[12];
      \nz.mem_355_sv2v_reg  <= w_data_i[11];
      \nz.mem_354_sv2v_reg  <= w_data_i[10];
      \nz.mem_353_sv2v_reg  <= w_data_i[9];
      \nz.mem_352_sv2v_reg  <= w_data_i[8];
      \nz.mem_351_sv2v_reg  <= w_data_i[7];
      \nz.mem_350_sv2v_reg  <= w_data_i[6];
      \nz.mem_349_sv2v_reg  <= w_data_i[5];
      \nz.mem_348_sv2v_reg  <= w_data_i[4];
      \nz.mem_347_sv2v_reg  <= w_data_i[3];
      \nz.mem_346_sv2v_reg  <= w_data_i[2];
      \nz.mem_345_sv2v_reg  <= w_data_i[1];
      \nz.mem_344_sv2v_reg  <= w_data_i[0];
    end 
    if(N66) begin
      \nz.mem_343_sv2v_reg  <= w_data_i[42];
      \nz.mem_342_sv2v_reg  <= w_data_i[41];
      \nz.mem_341_sv2v_reg  <= w_data_i[40];
      \nz.mem_340_sv2v_reg  <= w_data_i[39];
      \nz.mem_339_sv2v_reg  <= w_data_i[38];
      \nz.mem_338_sv2v_reg  <= w_data_i[37];
      \nz.mem_337_sv2v_reg  <= w_data_i[36];
      \nz.mem_336_sv2v_reg  <= w_data_i[35];
      \nz.mem_335_sv2v_reg  <= w_data_i[34];
      \nz.mem_334_sv2v_reg  <= w_data_i[33];
      \nz.mem_333_sv2v_reg  <= w_data_i[32];
      \nz.mem_332_sv2v_reg  <= w_data_i[31];
      \nz.mem_331_sv2v_reg  <= w_data_i[30];
      \nz.mem_330_sv2v_reg  <= w_data_i[29];
      \nz.mem_329_sv2v_reg  <= w_data_i[28];
      \nz.mem_328_sv2v_reg  <= w_data_i[27];
      \nz.mem_327_sv2v_reg  <= w_data_i[26];
      \nz.mem_326_sv2v_reg  <= w_data_i[25];
      \nz.mem_325_sv2v_reg  <= w_data_i[24];
      \nz.mem_324_sv2v_reg  <= w_data_i[23];
      \nz.mem_323_sv2v_reg  <= w_data_i[22];
      \nz.mem_322_sv2v_reg  <= w_data_i[21];
      \nz.mem_321_sv2v_reg  <= w_data_i[20];
      \nz.mem_320_sv2v_reg  <= w_data_i[19];
      \nz.mem_319_sv2v_reg  <= w_data_i[18];
      \nz.mem_318_sv2v_reg  <= w_data_i[17];
      \nz.mem_317_sv2v_reg  <= w_data_i[16];
      \nz.mem_316_sv2v_reg  <= w_data_i[15];
      \nz.mem_315_sv2v_reg  <= w_data_i[14];
      \nz.mem_314_sv2v_reg  <= w_data_i[13];
      \nz.mem_313_sv2v_reg  <= w_data_i[12];
      \nz.mem_312_sv2v_reg  <= w_data_i[11];
      \nz.mem_311_sv2v_reg  <= w_data_i[10];
      \nz.mem_310_sv2v_reg  <= w_data_i[9];
      \nz.mem_309_sv2v_reg  <= w_data_i[8];
      \nz.mem_308_sv2v_reg  <= w_data_i[7];
      \nz.mem_307_sv2v_reg  <= w_data_i[6];
      \nz.mem_306_sv2v_reg  <= w_data_i[5];
      \nz.mem_305_sv2v_reg  <= w_data_i[4];
      \nz.mem_304_sv2v_reg  <= w_data_i[3];
      \nz.mem_303_sv2v_reg  <= w_data_i[2];
      \nz.mem_302_sv2v_reg  <= w_data_i[1];
      \nz.mem_301_sv2v_reg  <= w_data_i[0];
    end 
    if(N65) begin
      \nz.mem_300_sv2v_reg  <= w_data_i[42];
      \nz.mem_299_sv2v_reg  <= w_data_i[41];
      \nz.mem_298_sv2v_reg  <= w_data_i[40];
      \nz.mem_297_sv2v_reg  <= w_data_i[39];
      \nz.mem_296_sv2v_reg  <= w_data_i[38];
      \nz.mem_295_sv2v_reg  <= w_data_i[37];
      \nz.mem_294_sv2v_reg  <= w_data_i[36];
      \nz.mem_293_sv2v_reg  <= w_data_i[35];
      \nz.mem_292_sv2v_reg  <= w_data_i[34];
      \nz.mem_291_sv2v_reg  <= w_data_i[33];
      \nz.mem_290_sv2v_reg  <= w_data_i[32];
      \nz.mem_289_sv2v_reg  <= w_data_i[31];
      \nz.mem_288_sv2v_reg  <= w_data_i[30];
      \nz.mem_287_sv2v_reg  <= w_data_i[29];
      \nz.mem_286_sv2v_reg  <= w_data_i[28];
      \nz.mem_285_sv2v_reg  <= w_data_i[27];
      \nz.mem_284_sv2v_reg  <= w_data_i[26];
      \nz.mem_283_sv2v_reg  <= w_data_i[25];
      \nz.mem_282_sv2v_reg  <= w_data_i[24];
      \nz.mem_281_sv2v_reg  <= w_data_i[23];
      \nz.mem_280_sv2v_reg  <= w_data_i[22];
      \nz.mem_279_sv2v_reg  <= w_data_i[21];
      \nz.mem_278_sv2v_reg  <= w_data_i[20];
      \nz.mem_277_sv2v_reg  <= w_data_i[19];
      \nz.mem_276_sv2v_reg  <= w_data_i[18];
      \nz.mem_275_sv2v_reg  <= w_data_i[17];
      \nz.mem_274_sv2v_reg  <= w_data_i[16];
      \nz.mem_273_sv2v_reg  <= w_data_i[15];
      \nz.mem_272_sv2v_reg  <= w_data_i[14];
      \nz.mem_271_sv2v_reg  <= w_data_i[13];
      \nz.mem_270_sv2v_reg  <= w_data_i[12];
      \nz.mem_269_sv2v_reg  <= w_data_i[11];
      \nz.mem_268_sv2v_reg  <= w_data_i[10];
      \nz.mem_267_sv2v_reg  <= w_data_i[9];
      \nz.mem_266_sv2v_reg  <= w_data_i[8];
      \nz.mem_265_sv2v_reg  <= w_data_i[7];
      \nz.mem_264_sv2v_reg  <= w_data_i[6];
      \nz.mem_263_sv2v_reg  <= w_data_i[5];
      \nz.mem_262_sv2v_reg  <= w_data_i[4];
      \nz.mem_261_sv2v_reg  <= w_data_i[3];
      \nz.mem_260_sv2v_reg  <= w_data_i[2];
      \nz.mem_259_sv2v_reg  <= w_data_i[1];
      \nz.mem_258_sv2v_reg  <= w_data_i[0];
    end 
    if(N64) begin
      \nz.mem_257_sv2v_reg  <= w_data_i[42];
      \nz.mem_256_sv2v_reg  <= w_data_i[41];
      \nz.mem_255_sv2v_reg  <= w_data_i[40];
      \nz.mem_254_sv2v_reg  <= w_data_i[39];
      \nz.mem_253_sv2v_reg  <= w_data_i[38];
      \nz.mem_252_sv2v_reg  <= w_data_i[37];
      \nz.mem_251_sv2v_reg  <= w_data_i[36];
      \nz.mem_250_sv2v_reg  <= w_data_i[35];
      \nz.mem_249_sv2v_reg  <= w_data_i[34];
      \nz.mem_248_sv2v_reg  <= w_data_i[33];
      \nz.mem_247_sv2v_reg  <= w_data_i[32];
      \nz.mem_246_sv2v_reg  <= w_data_i[31];
      \nz.mem_245_sv2v_reg  <= w_data_i[30];
      \nz.mem_244_sv2v_reg  <= w_data_i[29];
      \nz.mem_243_sv2v_reg  <= w_data_i[28];
      \nz.mem_242_sv2v_reg  <= w_data_i[27];
      \nz.mem_241_sv2v_reg  <= w_data_i[26];
      \nz.mem_240_sv2v_reg  <= w_data_i[25];
      \nz.mem_239_sv2v_reg  <= w_data_i[24];
      \nz.mem_238_sv2v_reg  <= w_data_i[23];
      \nz.mem_237_sv2v_reg  <= w_data_i[22];
      \nz.mem_236_sv2v_reg  <= w_data_i[21];
      \nz.mem_235_sv2v_reg  <= w_data_i[20];
      \nz.mem_234_sv2v_reg  <= w_data_i[19];
      \nz.mem_233_sv2v_reg  <= w_data_i[18];
      \nz.mem_232_sv2v_reg  <= w_data_i[17];
      \nz.mem_231_sv2v_reg  <= w_data_i[16];
      \nz.mem_230_sv2v_reg  <= w_data_i[15];
      \nz.mem_229_sv2v_reg  <= w_data_i[14];
      \nz.mem_228_sv2v_reg  <= w_data_i[13];
      \nz.mem_227_sv2v_reg  <= w_data_i[12];
      \nz.mem_226_sv2v_reg  <= w_data_i[11];
      \nz.mem_225_sv2v_reg  <= w_data_i[10];
      \nz.mem_224_sv2v_reg  <= w_data_i[9];
      \nz.mem_223_sv2v_reg  <= w_data_i[8];
      \nz.mem_222_sv2v_reg  <= w_data_i[7];
      \nz.mem_221_sv2v_reg  <= w_data_i[6];
      \nz.mem_220_sv2v_reg  <= w_data_i[5];
      \nz.mem_219_sv2v_reg  <= w_data_i[4];
      \nz.mem_218_sv2v_reg  <= w_data_i[3];
      \nz.mem_217_sv2v_reg  <= w_data_i[2];
      \nz.mem_216_sv2v_reg  <= w_data_i[1];
      \nz.mem_215_sv2v_reg  <= w_data_i[0];
    end 
    if(N63) begin
      \nz.mem_214_sv2v_reg  <= w_data_i[42];
      \nz.mem_213_sv2v_reg  <= w_data_i[41];
      \nz.mem_212_sv2v_reg  <= w_data_i[40];
      \nz.mem_211_sv2v_reg  <= w_data_i[39];
      \nz.mem_210_sv2v_reg  <= w_data_i[38];
      \nz.mem_209_sv2v_reg  <= w_data_i[37];
      \nz.mem_208_sv2v_reg  <= w_data_i[36];
      \nz.mem_207_sv2v_reg  <= w_data_i[35];
      \nz.mem_206_sv2v_reg  <= w_data_i[34];
      \nz.mem_205_sv2v_reg  <= w_data_i[33];
      \nz.mem_204_sv2v_reg  <= w_data_i[32];
      \nz.mem_203_sv2v_reg  <= w_data_i[31];
      \nz.mem_202_sv2v_reg  <= w_data_i[30];
      \nz.mem_201_sv2v_reg  <= w_data_i[29];
      \nz.mem_200_sv2v_reg  <= w_data_i[28];
      \nz.mem_199_sv2v_reg  <= w_data_i[27];
      \nz.mem_198_sv2v_reg  <= w_data_i[26];
      \nz.mem_197_sv2v_reg  <= w_data_i[25];
      \nz.mem_196_sv2v_reg  <= w_data_i[24];
      \nz.mem_195_sv2v_reg  <= w_data_i[23];
      \nz.mem_194_sv2v_reg  <= w_data_i[22];
      \nz.mem_193_sv2v_reg  <= w_data_i[21];
      \nz.mem_192_sv2v_reg  <= w_data_i[20];
      \nz.mem_191_sv2v_reg  <= w_data_i[19];
      \nz.mem_190_sv2v_reg  <= w_data_i[18];
      \nz.mem_189_sv2v_reg  <= w_data_i[17];
      \nz.mem_188_sv2v_reg  <= w_data_i[16];
      \nz.mem_187_sv2v_reg  <= w_data_i[15];
      \nz.mem_186_sv2v_reg  <= w_data_i[14];
      \nz.mem_185_sv2v_reg  <= w_data_i[13];
      \nz.mem_184_sv2v_reg  <= w_data_i[12];
      \nz.mem_183_sv2v_reg  <= w_data_i[11];
      \nz.mem_182_sv2v_reg  <= w_data_i[10];
      \nz.mem_181_sv2v_reg  <= w_data_i[9];
      \nz.mem_180_sv2v_reg  <= w_data_i[8];
      \nz.mem_179_sv2v_reg  <= w_data_i[7];
      \nz.mem_178_sv2v_reg  <= w_data_i[6];
      \nz.mem_177_sv2v_reg  <= w_data_i[5];
      \nz.mem_176_sv2v_reg  <= w_data_i[4];
      \nz.mem_175_sv2v_reg  <= w_data_i[3];
      \nz.mem_174_sv2v_reg  <= w_data_i[2];
      \nz.mem_173_sv2v_reg  <= w_data_i[1];
      \nz.mem_172_sv2v_reg  <= w_data_i[0];
    end 
    if(N62) begin
      \nz.mem_171_sv2v_reg  <= w_data_i[42];
      \nz.mem_170_sv2v_reg  <= w_data_i[41];
      \nz.mem_169_sv2v_reg  <= w_data_i[40];
      \nz.mem_168_sv2v_reg  <= w_data_i[39];
      \nz.mem_167_sv2v_reg  <= w_data_i[38];
      \nz.mem_166_sv2v_reg  <= w_data_i[37];
      \nz.mem_165_sv2v_reg  <= w_data_i[36];
      \nz.mem_164_sv2v_reg  <= w_data_i[35];
      \nz.mem_163_sv2v_reg  <= w_data_i[34];
      \nz.mem_162_sv2v_reg  <= w_data_i[33];
      \nz.mem_161_sv2v_reg  <= w_data_i[32];
      \nz.mem_160_sv2v_reg  <= w_data_i[31];
      \nz.mem_159_sv2v_reg  <= w_data_i[30];
      \nz.mem_158_sv2v_reg  <= w_data_i[29];
      \nz.mem_157_sv2v_reg  <= w_data_i[28];
      \nz.mem_156_sv2v_reg  <= w_data_i[27];
      \nz.mem_155_sv2v_reg  <= w_data_i[26];
      \nz.mem_154_sv2v_reg  <= w_data_i[25];
      \nz.mem_153_sv2v_reg  <= w_data_i[24];
      \nz.mem_152_sv2v_reg  <= w_data_i[23];
      \nz.mem_151_sv2v_reg  <= w_data_i[22];
      \nz.mem_150_sv2v_reg  <= w_data_i[21];
      \nz.mem_149_sv2v_reg  <= w_data_i[20];
      \nz.mem_148_sv2v_reg  <= w_data_i[19];
      \nz.mem_147_sv2v_reg  <= w_data_i[18];
      \nz.mem_146_sv2v_reg  <= w_data_i[17];
      \nz.mem_145_sv2v_reg  <= w_data_i[16];
      \nz.mem_144_sv2v_reg  <= w_data_i[15];
      \nz.mem_143_sv2v_reg  <= w_data_i[14];
      \nz.mem_142_sv2v_reg  <= w_data_i[13];
      \nz.mem_141_sv2v_reg  <= w_data_i[12];
      \nz.mem_140_sv2v_reg  <= w_data_i[11];
      \nz.mem_139_sv2v_reg  <= w_data_i[10];
      \nz.mem_138_sv2v_reg  <= w_data_i[9];
      \nz.mem_137_sv2v_reg  <= w_data_i[8];
      \nz.mem_136_sv2v_reg  <= w_data_i[7];
      \nz.mem_135_sv2v_reg  <= w_data_i[6];
      \nz.mem_134_sv2v_reg  <= w_data_i[5];
      \nz.mem_133_sv2v_reg  <= w_data_i[4];
      \nz.mem_132_sv2v_reg  <= w_data_i[3];
      \nz.mem_131_sv2v_reg  <= w_data_i[2];
      \nz.mem_130_sv2v_reg  <= w_data_i[1];
      \nz.mem_129_sv2v_reg  <= w_data_i[0];
    end 
    if(N61) begin
      \nz.mem_128_sv2v_reg  <= w_data_i[42];
      \nz.mem_127_sv2v_reg  <= w_data_i[41];
      \nz.mem_126_sv2v_reg  <= w_data_i[40];
      \nz.mem_125_sv2v_reg  <= w_data_i[39];
      \nz.mem_124_sv2v_reg  <= w_data_i[38];
      \nz.mem_123_sv2v_reg  <= w_data_i[37];
      \nz.mem_122_sv2v_reg  <= w_data_i[36];
      \nz.mem_121_sv2v_reg  <= w_data_i[35];
      \nz.mem_120_sv2v_reg  <= w_data_i[34];
      \nz.mem_119_sv2v_reg  <= w_data_i[33];
      \nz.mem_118_sv2v_reg  <= w_data_i[32];
      \nz.mem_117_sv2v_reg  <= w_data_i[31];
      \nz.mem_116_sv2v_reg  <= w_data_i[30];
      \nz.mem_115_sv2v_reg  <= w_data_i[29];
      \nz.mem_114_sv2v_reg  <= w_data_i[28];
      \nz.mem_113_sv2v_reg  <= w_data_i[27];
      \nz.mem_112_sv2v_reg  <= w_data_i[26];
      \nz.mem_111_sv2v_reg  <= w_data_i[25];
      \nz.mem_110_sv2v_reg  <= w_data_i[24];
      \nz.mem_109_sv2v_reg  <= w_data_i[23];
      \nz.mem_108_sv2v_reg  <= w_data_i[22];
      \nz.mem_107_sv2v_reg  <= w_data_i[21];
      \nz.mem_106_sv2v_reg  <= w_data_i[20];
      \nz.mem_105_sv2v_reg  <= w_data_i[19];
      \nz.mem_104_sv2v_reg  <= w_data_i[18];
      \nz.mem_103_sv2v_reg  <= w_data_i[17];
      \nz.mem_102_sv2v_reg  <= w_data_i[16];
      \nz.mem_101_sv2v_reg  <= w_data_i[15];
      \nz.mem_100_sv2v_reg  <= w_data_i[14];
      \nz.mem_99_sv2v_reg  <= w_data_i[13];
      \nz.mem_98_sv2v_reg  <= w_data_i[12];
      \nz.mem_97_sv2v_reg  <= w_data_i[11];
      \nz.mem_96_sv2v_reg  <= w_data_i[10];
      \nz.mem_95_sv2v_reg  <= w_data_i[9];
      \nz.mem_94_sv2v_reg  <= w_data_i[8];
      \nz.mem_93_sv2v_reg  <= w_data_i[7];
      \nz.mem_92_sv2v_reg  <= w_data_i[6];
      \nz.mem_91_sv2v_reg  <= w_data_i[5];
      \nz.mem_90_sv2v_reg  <= w_data_i[4];
      \nz.mem_89_sv2v_reg  <= w_data_i[3];
      \nz.mem_88_sv2v_reg  <= w_data_i[2];
      \nz.mem_87_sv2v_reg  <= w_data_i[1];
      \nz.mem_86_sv2v_reg  <= w_data_i[0];
    end 
    if(N60) begin
      \nz.mem_85_sv2v_reg  <= w_data_i[42];
      \nz.mem_84_sv2v_reg  <= w_data_i[41];
      \nz.mem_83_sv2v_reg  <= w_data_i[40];
      \nz.mem_82_sv2v_reg  <= w_data_i[39];
      \nz.mem_81_sv2v_reg  <= w_data_i[38];
      \nz.mem_80_sv2v_reg  <= w_data_i[37];
      \nz.mem_79_sv2v_reg  <= w_data_i[36];
      \nz.mem_78_sv2v_reg  <= w_data_i[35];
      \nz.mem_77_sv2v_reg  <= w_data_i[34];
      \nz.mem_76_sv2v_reg  <= w_data_i[33];
      \nz.mem_75_sv2v_reg  <= w_data_i[32];
      \nz.mem_74_sv2v_reg  <= w_data_i[31];
      \nz.mem_73_sv2v_reg  <= w_data_i[30];
      \nz.mem_72_sv2v_reg  <= w_data_i[29];
      \nz.mem_71_sv2v_reg  <= w_data_i[28];
      \nz.mem_70_sv2v_reg  <= w_data_i[27];
      \nz.mem_69_sv2v_reg  <= w_data_i[26];
      \nz.mem_68_sv2v_reg  <= w_data_i[25];
      \nz.mem_67_sv2v_reg  <= w_data_i[24];
      \nz.mem_66_sv2v_reg  <= w_data_i[23];
      \nz.mem_65_sv2v_reg  <= w_data_i[22];
      \nz.mem_64_sv2v_reg  <= w_data_i[21];
      \nz.mem_63_sv2v_reg  <= w_data_i[20];
      \nz.mem_62_sv2v_reg  <= w_data_i[19];
      \nz.mem_61_sv2v_reg  <= w_data_i[18];
      \nz.mem_60_sv2v_reg  <= w_data_i[17];
      \nz.mem_59_sv2v_reg  <= w_data_i[16];
      \nz.mem_58_sv2v_reg  <= w_data_i[15];
      \nz.mem_57_sv2v_reg  <= w_data_i[14];
      \nz.mem_56_sv2v_reg  <= w_data_i[13];
      \nz.mem_55_sv2v_reg  <= w_data_i[12];
      \nz.mem_54_sv2v_reg  <= w_data_i[11];
      \nz.mem_53_sv2v_reg  <= w_data_i[10];
      \nz.mem_52_sv2v_reg  <= w_data_i[9];
      \nz.mem_51_sv2v_reg  <= w_data_i[8];
      \nz.mem_50_sv2v_reg  <= w_data_i[7];
      \nz.mem_49_sv2v_reg  <= w_data_i[6];
      \nz.mem_48_sv2v_reg  <= w_data_i[5];
      \nz.mem_47_sv2v_reg  <= w_data_i[4];
      \nz.mem_46_sv2v_reg  <= w_data_i[3];
      \nz.mem_45_sv2v_reg  <= w_data_i[2];
      \nz.mem_44_sv2v_reg  <= w_data_i[1];
      \nz.mem_43_sv2v_reg  <= w_data_i[0];
    end 
    if(N59) begin
      \nz.mem_42_sv2v_reg  <= w_data_i[42];
      \nz.mem_41_sv2v_reg  <= w_data_i[41];
      \nz.mem_40_sv2v_reg  <= w_data_i[40];
      \nz.mem_39_sv2v_reg  <= w_data_i[39];
      \nz.mem_38_sv2v_reg  <= w_data_i[38];
      \nz.mem_37_sv2v_reg  <= w_data_i[37];
      \nz.mem_36_sv2v_reg  <= w_data_i[36];
      \nz.mem_35_sv2v_reg  <= w_data_i[35];
      \nz.mem_34_sv2v_reg  <= w_data_i[34];
      \nz.mem_33_sv2v_reg  <= w_data_i[33];
      \nz.mem_32_sv2v_reg  <= w_data_i[32];
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_0000002b_16_1
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [3:0] w_addr_i;
  input [42:0] w_data_i;
  input [3:0] r_addr_i;
  output [42:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [42:0] r_data_o;

  bsg_mem_1r1w_synth_0000002b_16_1
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bp_fe_ras_00
(
  clk_i,
  reset_i,
  init_done_o,
  restore_i,
  w_next_i,
  w_tos_i,
  call_i,
  addr_i,
  v_o,
  tgt_o,
  next_o,
  tos_o,
  return_i
);

  input [3:0] w_next_i;
  input [3:0] w_tos_i;
  input [38:0] addr_i;
  output [38:0] tgt_o;
  output [3:0] next_o;
  output [3:0] tos_o;
  input clk_i;
  input reset_i;
  input restore_i;
  input call_i;
  input return_i;
  output init_done_o;
  output v_o;
  wire [38:0] tgt_o;
  wire [3:0] next_o,tos_o,next_n,tos_n,nos_lo,w_addr_li;
  wire init_done_o,v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,
  N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,w_v_li,N30,N31,N32,N33,N34,N36,
  N37,N38,N39,N40,N41,N42,N43,N44;
  wire [1:0] state_r,state_n;
  wire [4:0] init_cnt;
  wire [42:0] w_data_li;
  reg state_r_1_sv2v_reg,state_r_0_sv2v_reg;
  assign state_r[1] = state_r_1_sv2v_reg;
  assign state_r[0] = state_r_0_sv2v_reg;
  assign v_o = 1'b1;

  bsg_counter_clear_up_max_val_p16_init_val_p0
  init_counter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(1'b0),
    .up_i(N32),
    .count_o(init_cnt)
  );

  assign N6 = state_r[1] | N30;
  assign N8 = N33 | state_r[0];
  assign N10 = state_r[1] & state_r[0];
  assign N11 = N33 & N30;

  bsg_dff_reset_00000008
  ptr_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ next_n, tos_n }),
    .data_o({ next_o, tos_o })
  );


  bsg_mem_1r1w_0000002b_16_1
  mem
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(w_v_li),
    .w_addr_i(w_addr_li),
    .w_data_i(w_data_li),
    .r_v_i(return_i),
    .r_addr_i(tos_o),
    .r_data_o({ nos_lo, tgt_o })
  );

  assign N30 = ~state_r[0];
  assign N31 = N30 | state_r[1];
  assign N32 = ~N31;
  assign N33 = ~state_r[1];
  assign N34 = state_r[0] | N33;
  assign init_done_o = ~N34;
  assign N36 = ~init_cnt[3];
  assign N37 = ~init_cnt[2];
  assign N38 = ~init_cnt[1];
  assign N39 = ~init_cnt[0];
  assign N40 = N36 | init_cnt[4];
  assign N41 = N37 | N40;
  assign N42 = N38 | N41;
  assign N43 = N39 | N42;
  assign N44 = ~N43;
  assign { N19, N18, N17, N16 } = next_o + 1'b1;
  assign state_n = (N0)? { N44, N43 } : 
                   (N1)? { 1'b1, 1'b0 } : 
                   (N2)? { 1'b0, 1'b1 } : 1'b0;
  assign N0 = N7;
  assign N1 = N9;
  assign N2 = N12;
  assign next_n = (N3)? w_next_i : 
                  (N21)? { N19, N18, N17, N16 } : 
                  (N14)? next_o : 1'b0;
  assign N3 = restore_i;
  assign tos_n = (N3)? w_tos_i : 
                 (N26)? next_o : 
                 (N29)? nos_lo : 
                 (N25)? tos_o : 1'b0;
  assign w_v_li = (N4)? call_i : 
                  (N5)? 1'b1 : 1'b0;
  assign N4 = init_done_o;
  assign N5 = N34;
  assign w_addr_li = (N4)? next_o : 
                     (N5)? init_cnt[3:0] : 1'b0;
  assign w_data_li = (N4)? { tos_o, addr_i } : 
                     (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N7 = ~N6;
  assign N9 = ~N8;
  assign N12 = N10 | N11;
  assign N13 = call_i | restore_i;
  assign N14 = ~N13;
  assign N15 = N21;
  assign N20 = ~restore_i;
  assign N21 = call_i & N20;
  assign N22 = return_i;
  assign N23 = call_i | restore_i;
  assign N24 = N22 | N23;
  assign N25 = ~N24;
  assign N26 = call_i & N20;
  assign N27 = ~call_i;
  assign N28 = N20 & N27;
  assign N29 = N22 & N28;

  always @(posedge clk_i) begin
    if(reset_i) begin
      state_r_1_sv2v_reg <= 1'b0;
      state_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      state_r_1_sv2v_reg <= state_n[1];
      state_r_0_sv2v_reg <= state_n[0];
    end 
  end


endmodule



module bsg_dff_reset_en_00000002
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [1:0] data_i;
  output [1:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [1:0] data_o;
  wire N0,N1,N2;
  reg data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bp_fe_pc_gen_00
(
  clk_i,
  reset_i,
  init_done_o,
  attaboy_v_i,
  attaboy_force_i,
  attaboy_pc_i,
  attaboy_br_metadata_fwd_i,
  attaboy_taken_i,
  attaboy_ntaken_i,
  attaboy_yumi_o,
  redirect_v_i,
  redirect_pc_i,
  redirect_npc_i,
  redirect_br_v_i,
  redirect_br_metadata_fwd_i,
  redirect_br_taken_i,
  redirect_br_ntaken_i,
  redirect_br_nonbr_i,
  next_pc_o,
  icache_yumi_i,
  ovr_o,
  icache_tv_we_i,
  icache_hit_v_i,
  icache_miss_v_i,
  icache_hit_yumi_o,
  icache_data_i,
  if2_hit_v_o,
  if2_miss_v_o,
  if2_pc_o,
  if2_data_o,
  if2_br_metadata_fwd_o,
  if2_yumi_i,
  fetch_yumi_i,
  fetch_scan_i,
  fetch_pc_i,
  fetch_count_i,
  fetch_startup_i,
  fetch_catchup_i,
  fetch_rebase_i,
  fetch_linear_i,
  fetch_taken_o
);

  input [38:0] attaboy_pc_i;
  input [48:0] attaboy_br_metadata_fwd_i;
  input [38:0] redirect_pc_i;
  input [38:0] redirect_npc_i;
  input [48:0] redirect_br_metadata_fwd_i;
  output [38:0] next_pc_o;
  input [63:0] icache_data_i;
  output [38:0] if2_pc_o;
  output [63:0] if2_data_o;
  output [48:0] if2_br_metadata_fwd_o;
  input [124:0] fetch_scan_i;
  input [38:0] fetch_pc_i;
  input [2:0] fetch_count_i;
  input clk_i;
  input reset_i;
  input attaboy_v_i;
  input attaboy_force_i;
  input attaboy_taken_i;
  input attaboy_ntaken_i;
  input redirect_v_i;
  input redirect_br_v_i;
  input redirect_br_taken_i;
  input redirect_br_ntaken_i;
  input redirect_br_nonbr_i;
  input icache_yumi_i;
  input icache_tv_we_i;
  input icache_hit_v_i;
  input icache_miss_v_i;
  input if2_yumi_i;
  input fetch_yumi_i;
  input fetch_startup_i;
  input fetch_catchup_i;
  input fetch_rebase_i;
  input fetch_linear_i;
  output init_done_o;
  output attaboy_yumi_o;
  output ovr_o;
  output icache_hit_yumi_o;
  output if2_hit_v_o;
  output if2_miss_v_o;
  output fetch_taken_o;
  wire [38:0] next_pc_o,if2_pc_o,ras_tgt_lo,taken_tgt_lo,ntaken_tgt_lo,linear_tgt_lo,
  btb_br_tgt_lo,pc_plus,btb_tgt_li,pc_if1;
  wire [63:0] if2_data_o;
  wire [48:0] if2_br_metadata_fwd_o,next_metadata,metadata_if1,metadata_if2_n;
  wire init_done_o,attaboy_yumi_o,ovr_o,icache_hit_yumi_o,if2_hit_v_o,if2_miss_v_o,
  fetch_taken_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,next_pred,next_taken,ovr_btaken,ovr_ret,
  ovr_jmp,N29,N30,ovr_rebase,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,
  N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,
  N65,N66,N67,N68,N69,N70,N71,N72,bht_pred_lo,btb_taken,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,
  btb_br_tgt_v_lo,N113,N114,N115,N116,N117,N118,N119,btb_w_v_li,btb_w_force_li,btb_clr_li,N120,
  N121,N122,btb_jmp_li,N123,N124,N125,N126,N127,N128,N129,btb_br_tgt_jmp_lo,
  btb_w_yumi_lo,btb_init_done_lo,bht_w_v_li,bht_w_force_li,N130,N131,N132,N133,N134,N135,
  N136,N137,bht_w_yumi_lo,bht_init_done_lo,metadata_if1_r_site_br_,
  metadata_if1_r_site_jal_,metadata_if1_r_site_jalr_,metadata_if1_r_site_call_,
  metadata_if1_r_site_return_,pred_if1_r,N138,N139,N140,_2_net_,metadata_if2_r_ras_next__3_,
  metadata_if2_r_ras_next__2_,metadata_if2_r_ras_next__1_,metadata_if2_r_ras_next__0_,
  metadata_if2_r_ras_tos__3_,metadata_if2_r_ras_tos__2_,metadata_if2_r_ras_tos__1_,
  metadata_if2_r_ras_tos__0_,pred_if2_r,taken_if2_r,ras_init_done_lo,ras_call_li,
  ras_valid_lo,ras_return_li,btb_miss_ras,btb_miss_br,rebase_miss,linear_miss,
  ovr_linear,N141,N142,N143,N144,N145,N146,ghistory_w_v,N147,N148,N149,N150,N151,N152,
  N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,
  N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,
  N185,N186,N187,N188,N189;
  wire [7:0] bht_row_lo,bht_row_li;
  wire [1:0] ghistory_r,bht_offset,bht_r_ghist_li,bht_w_offset_li,bht_w_ghist_li;
  wire [8:0] btb_tag,btb_tag_li;
  wire [5:0] btb_idx,btb_idx_li;
  wire [6:0] bht_idx,bht_w_idx_li;
  wire [2:0] pc_if1_r;
  wire [38:3] pc_if1_aligned;
  assign if2_hit_v_o = icache_hit_v_i;
  assign if2_miss_v_o = icache_miss_v_i;
  assign if2_data_o[63] = icache_data_i[63];
  assign if2_data_o[62] = icache_data_i[62];
  assign if2_data_o[61] = icache_data_i[61];
  assign if2_data_o[60] = icache_data_i[60];
  assign if2_data_o[59] = icache_data_i[59];
  assign if2_data_o[58] = icache_data_i[58];
  assign if2_data_o[57] = icache_data_i[57];
  assign if2_data_o[56] = icache_data_i[56];
  assign if2_data_o[55] = icache_data_i[55];
  assign if2_data_o[54] = icache_data_i[54];
  assign if2_data_o[53] = icache_data_i[53];
  assign if2_data_o[52] = icache_data_i[52];
  assign if2_data_o[51] = icache_data_i[51];
  assign if2_data_o[50] = icache_data_i[50];
  assign if2_data_o[49] = icache_data_i[49];
  assign if2_data_o[48] = icache_data_i[48];
  assign if2_data_o[47] = icache_data_i[47];
  assign if2_data_o[46] = icache_data_i[46];
  assign if2_data_o[45] = icache_data_i[45];
  assign if2_data_o[44] = icache_data_i[44];
  assign if2_data_o[43] = icache_data_i[43];
  assign if2_data_o[42] = icache_data_i[42];
  assign if2_data_o[41] = icache_data_i[41];
  assign if2_data_o[40] = icache_data_i[40];
  assign if2_data_o[39] = icache_data_i[39];
  assign if2_data_o[38] = icache_data_i[38];
  assign if2_data_o[37] = icache_data_i[37];
  assign if2_data_o[36] = icache_data_i[36];
  assign if2_data_o[35] = icache_data_i[35];
  assign if2_data_o[34] = icache_data_i[34];
  assign if2_data_o[33] = icache_data_i[33];
  assign if2_data_o[32] = icache_data_i[32];
  assign if2_data_o[31] = icache_data_i[31];
  assign if2_data_o[30] = icache_data_i[30];
  assign if2_data_o[29] = icache_data_i[29];
  assign if2_data_o[28] = icache_data_i[28];
  assign if2_data_o[27] = icache_data_i[27];
  assign if2_data_o[26] = icache_data_i[26];
  assign if2_data_o[25] = icache_data_i[25];
  assign if2_data_o[24] = icache_data_i[24];
  assign if2_data_o[23] = icache_data_i[23];
  assign if2_data_o[22] = icache_data_i[22];
  assign if2_data_o[21] = icache_data_i[21];
  assign if2_data_o[20] = icache_data_i[20];
  assign if2_data_o[19] = icache_data_i[19];
  assign if2_data_o[18] = icache_data_i[18];
  assign if2_data_o[17] = icache_data_i[17];
  assign if2_data_o[16] = icache_data_i[16];
  assign if2_data_o[15] = icache_data_i[15];
  assign if2_data_o[14] = icache_data_i[14];
  assign if2_data_o[13] = icache_data_i[13];
  assign if2_data_o[12] = icache_data_i[12];
  assign if2_data_o[11] = icache_data_i[11];
  assign if2_data_o[10] = icache_data_i[10];
  assign if2_data_o[9] = icache_data_i[9];
  assign if2_data_o[8] = icache_data_i[8];
  assign if2_data_o[7] = icache_data_i[7];
  assign if2_data_o[6] = icache_data_i[6];
  assign if2_data_o[5] = icache_data_i[5];
  assign if2_data_o[4] = icache_data_i[4];
  assign if2_data_o[3] = icache_data_i[3];
  assign if2_data_o[2] = icache_data_i[2];
  assign if2_data_o[1] = icache_data_i[1];
  assign if2_data_o[0] = icache_data_i[0];

  bp_fe_btb_00
  btb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .init_done_o(btb_init_done_lo),
    .r_addr_i(next_pc_o),
    .r_v_i(icache_yumi_i),
    .r_tag_o(btb_tag),
    .r_idx_o(btb_idx),
    .r_tgt_o(btb_br_tgt_lo),
    .r_tgt_v_o(btb_br_tgt_v_lo),
    .r_tgt_jmp_o(btb_br_tgt_jmp_lo),
    .w_v_i(btb_w_v_li),
    .w_force_i(btb_w_force_li),
    .w_clr_i(btb_clr_li),
    .w_jmp_i(btb_jmp_li),
    .w_tag_i(btb_tag_li),
    .w_idx_i(btb_idx_li),
    .w_tgt_i(btb_tgt_li),
    .w_yumi_o(btb_w_yumi_lo)
  );


  bp_fe_bht_00
  bht
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .init_done_o(bht_init_done_lo),
    .w_v_i(bht_w_v_li),
    .w_force_i(bht_w_force_li),
    .w_idx_i(bht_w_idx_li),
    .w_offset_i(bht_w_offset_li),
    .w_ghist_i(bht_w_ghist_li),
    .w_val_i(bht_row_li),
    .w_correct_i(attaboy_yumi_o),
    .w_yumi_o(bht_w_yumi_lo),
    .r_v_i(icache_yumi_i),
    .r_addr_i(next_pc_o),
    .r_ghist_i(bht_r_ghist_li),
    .r_val_o(bht_row_lo),
    .r_pred_o(bht_pred_lo),
    .r_idx_o(bht_idx),
    .r_offset_o(bht_offset)
  );


  bsg_dff_reset_en_0000005a
  if1_stage_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(icache_yumi_i),
    .data_i({ next_pred, next_taken, next_metadata, next_pc_o }),
    .data_o({ pred_if1_r, linear_miss, metadata_if1_r_site_br_, metadata_if1_r_site_jal_, metadata_if1_r_site_jalr_, metadata_if1_r_site_call_, metadata_if1_r_site_return_, metadata_if1[43:0], pc_if1_aligned, pc_if1_r })
  );


  bsg_dff_reset_en_0000005a
  if2_stage_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(_2_net_),
    .data_i({ pred_if1_r, linear_miss, pc_if1, metadata_if2_n }),
    .data_o({ pred_if2_r, taken_if2_r, if2_pc_o, if2_br_metadata_fwd_o[48:42], metadata_if2_r_ras_next__3_, metadata_if2_r_ras_next__2_, metadata_if2_r_ras_next__1_, metadata_if2_r_ras_next__0_, metadata_if2_r_ras_tos__3_, metadata_if2_r_ras_tos__2_, metadata_if2_r_ras_tos__1_, metadata_if2_r_ras_tos__0_, if2_br_metadata_fwd_o[33:0] })
  );


  bp_fe_ras_00
  ras
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .init_done_o(ras_init_done_lo),
    .restore_i(redirect_br_v_i),
    .w_next_i(redirect_br_metadata_fwd_i[41:38]),
    .w_tos_i(redirect_br_metadata_fwd_i[37:34]),
    .call_i(ras_call_li),
    .addr_i(ntaken_tgt_lo),
    .v_o(ras_valid_lo),
    .tgt_o(ras_tgt_lo),
    .next_o(if2_br_metadata_fwd_o[41:38]),
    .tos_o(if2_br_metadata_fwd_o[37:34]),
    .return_i(ras_return_li)
  );

  assign btb_miss_ras = { pc_if1_aligned, pc_if1_r } != ras_tgt_lo;
  assign btb_miss_br = { pc_if1_aligned, pc_if1_r } != taken_tgt_lo;

  bsg_dff_reset_en_00000002
  ghist_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(ghistory_w_v),
    .data_i(bht_r_ghist_li),
    .data_o(ghistory_r)
  );

  assign ntaken_tgt_lo = fetch_pc_i + fetch_scan_i[77:39];
  assign linear_tgt_lo = fetch_pc_i + fetch_scan_i[116:78];
  assign taken_tgt_lo = fetch_pc_i + fetch_scan_i[38:0];
  assign pc_plus = { pc_if1_aligned, 1'b0, 1'b0, 1'b0 } + { 1'b1, 1'b0, 1'b0, 1'b0 };
  assign { N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34 } = (N0)? ras_tgt_lo : 
                                                                                                                                                                                                                 (N116)? taken_tgt_lo : 
                                                                                                                                                                                                                 (N119)? ntaken_tgt_lo : 
                                                                                                                                                                                                                 (N33)? linear_tgt_lo : 1'b0;
  assign N0 = ovr_ret;
  assign { N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74 } = (N1)? btb_br_tgt_lo : 
                                                                                                                                                                                                                              (N2)? pc_plus : 1'b0;
  assign N1 = btb_taken;
  assign N2 = N73;
  assign next_pred = (N3)? 1'b0 : 
                     (N114)? ovr_btaken : 
                     (N28)? bht_pred_lo : 1'b0;
  assign N3 = redirect_v_i;
  assign next_taken = (N3)? redirect_br_taken_i : 
                      (N114)? N29 : 
                      (N28)? btb_taken : 1'b0;
  assign next_pc_o = (N3)? redirect_npc_i : 
                     (N114)? { N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34 } : 
                     (N28)? { N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74 } : 1'b0;
  assign next_metadata = (N3)? redirect_br_metadata_fwd_i : 
                         (N114)? { metadata_if1[48:44], ovr_ret, metadata_if1[42:0] } : 
                         (N28)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, btb_br_tgt_v_lo, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, btb_tag, btb_idx, bht_idx, bht_row_lo, bht_offset, ghistory_r } : 1'b0;
  assign btb_jmp_li = (N4)? N122 : 
                      (N5)? N123 : 1'b0;
  assign N4 = N121;
  assign N5 = N120;
  assign btb_tag_li = (N6)? redirect_br_metadata_fwd_i[33:25] : 
                      (N7)? attaboy_br_metadata_fwd_i[33:25] : 1'b0;
  assign N6 = N125;
  assign N7 = N124;
  assign btb_idx_li = (N8)? redirect_br_metadata_fwd_i[24:19] : 
                      (N9)? attaboy_br_metadata_fwd_i[24:19] : 1'b0;
  assign N8 = N127;
  assign N9 = N126;
  assign btb_tgt_li = (N10)? redirect_pc_i : 
                      (N11)? attaboy_pc_i : 1'b0;
  assign N10 = N129;
  assign N11 = N128;
  assign bht_w_idx_li = (N12)? redirect_br_metadata_fwd_i[18:12] : 
                        (N13)? attaboy_br_metadata_fwd_i[18:12] : 1'b0;
  assign N12 = N131;
  assign N13 = N130;
  assign bht_w_offset_li = (N14)? redirect_br_metadata_fwd_i[3:2] : 
                           (N15)? attaboy_br_metadata_fwd_i[3:2] : 1'b0;
  assign N14 = N133;
  assign N15 = N132;
  assign bht_w_ghist_li = (N16)? redirect_br_metadata_fwd_i[1:0] : 
                          (N17)? attaboy_br_metadata_fwd_i[1:0] : 1'b0;
  assign N16 = N135;
  assign N17 = N134;
  assign bht_row_li = (N18)? redirect_br_metadata_fwd_i[11:4] : 
                      (N19)? attaboy_br_metadata_fwd_i[11:4] : 1'b0;
  assign N18 = N137;
  assign N19 = N136;
  assign metadata_if1[48:44] = (N20)? fetch_scan_i[121:117] : 
                               (N21)? { metadata_if1_r_site_br_, metadata_if1_r_site_jal_, metadata_if1_r_site_jalr_, metadata_if1_r_site_call_, metadata_if1_r_site_return_ } : 1'b0;
  assign N20 = fetch_yumi_i;
  assign N21 = N138;
  assign pc_if1 = (N22)? ntaken_tgt_lo : 
                  (N23)? { pc_if1_aligned, pc_if1_r } : 1'b0;
  assign N22 = fetch_catchup_i;
  assign N23 = N139;
  assign metadata_if2_n = (N24)? if2_br_metadata_fwd_o : 
                          (N25)? metadata_if1 : 1'b0;
  assign N24 = fetch_startup_i;
  assign N25 = N140;
  assign bht_r_ghist_li = (N26)? redirect_br_metadata_fwd_i[1:0] : 
                          (N146)? { ghistory_r[0:0], linear_miss } : 
                          (N144)? ghistory_r : 1'b0;
  assign N26 = N142;
  assign N27 = ovr_o | redirect_v_i;
  assign N28 = ~N27;
  assign N29 = N147 | ovr_jmp;
  assign N147 = ovr_ret | ovr_btaken;
  assign N30 = ovr_btaken | ovr_jmp;
  assign N31 = N30 | ovr_ret;
  assign N32 = ovr_rebase | N31;
  assign N33 = ~N32;
  assign N73 = ~btb_taken;
  assign N113 = ~redirect_v_i;
  assign N114 = ovr_o & N113;
  assign N115 = ~ovr_ret;
  assign N116 = N30 & N115;
  assign N117 = ~N30;
  assign N118 = N115 & N117;
  assign N119 = ovr_rebase & N118;
  assign btb_w_v_li = N163 | N165;
  assign N163 = N161 | N162;
  assign N161 = N155 | N160;
  assign N155 = N152 | N154;
  assign N152 = N150 & N151;
  assign N150 = N148 & N149;
  assign N148 = redirect_br_v_i & redirect_br_taken_i;
  assign N149 = ~redirect_br_metadata_fwd_i[42];
  assign N151 = ~redirect_br_metadata_fwd_i[43];
  assign N154 = N153 & N151;
  assign N153 = N148 & redirect_br_metadata_fwd_i[42];
  assign N160 = N158 & N159;
  assign N158 = N156 & N157;
  assign N156 = attaboy_v_i & attaboy_taken_i;
  assign N157 = ~attaboy_br_metadata_fwd_i[42];
  assign N159 = ~attaboy_br_metadata_fwd_i[43];
  assign N162 = N153 & redirect_br_metadata_fwd_i[43];
  assign N165 = N164 & redirect_br_metadata_fwd_i[42];
  assign N164 = redirect_br_v_i & redirect_br_nonbr_i;
  assign btb_w_force_li = redirect_br_v_i | attaboy_force_i;
  assign btb_clr_li = N168 | N170;
  assign N168 = N167 & redirect_br_metadata_fwd_i[43];
  assign N167 = N166 & redirect_br_metadata_fwd_i[42];
  assign N166 = redirect_br_v_i & redirect_br_taken_i;
  assign N170 = N169 & redirect_br_metadata_fwd_i[42];
  assign N169 = redirect_br_v_i & redirect_br_nonbr_i;
  assign N120 = ~redirect_br_v_i;
  assign N121 = redirect_br_v_i;
  assign N122 = redirect_br_metadata_fwd_i[47] | redirect_br_metadata_fwd_i[46];
  assign N123 = attaboy_br_metadata_fwd_i[47] | attaboy_br_metadata_fwd_i[46];
  assign N124 = ~redirect_br_v_i;
  assign N125 = redirect_br_v_i;
  assign N126 = ~redirect_br_v_i;
  assign N127 = redirect_br_v_i;
  assign N128 = ~redirect_br_v_i;
  assign N129 = redirect_br_v_i;
  assign bht_w_v_li = N171 | N172;
  assign N171 = redirect_br_v_i & redirect_br_metadata_fwd_i[48];
  assign N172 = attaboy_v_i & attaboy_br_metadata_fwd_i[48];
  assign bht_w_force_li = redirect_br_v_i | attaboy_force_i;
  assign N130 = ~redirect_br_v_i;
  assign N131 = redirect_br_v_i;
  assign N132 = ~redirect_br_v_i;
  assign N133 = redirect_br_v_i;
  assign N134 = ~redirect_br_v_i;
  assign N135 = redirect_br_v_i;
  assign N136 = ~redirect_br_v_i;
  assign N137 = redirect_br_v_i;
  assign N138 = ~fetch_yumi_i;
  assign N139 = ~fetch_catchup_i;
  assign btb_taken = btb_br_tgt_v_lo & N173;
  assign N173 = bht_pred_lo | btb_br_tgt_jmp_lo;
  assign N140 = ~fetch_startup_i;
  assign _2_net_ = icache_tv_we_i | fetch_catchup_i;
  assign icache_hit_yumi_o = if2_hit_v_o & if2_yumi_i;
  assign ras_call_li = fetch_yumi_i & fetch_scan_i[118];
  assign ras_return_li = fetch_yumi_i & fetch_scan_i[117];
  assign rebase_miss = ~linear_miss;
  assign ovr_ret = N174 & ras_valid_lo;
  assign N174 = btb_miss_ras & fetch_scan_i[117];
  assign ovr_btaken = N175 & pred_if1_r;
  assign N175 = btb_miss_br & fetch_scan_i[121];
  assign ovr_jmp = btb_miss_br & fetch_scan_i[120];
  assign ovr_linear = linear_miss & fetch_linear_i;
  assign ovr_rebase = rebase_miss & fetch_rebase_i;
  assign ovr_o = N178 | ovr_rebase;
  assign N178 = N177 | ovr_linear;
  assign N177 = N176 | ovr_ret;
  assign N176 = ovr_btaken | ovr_jmp;
  assign fetch_taken_o = N180 | ovr_jmp;
  assign N180 = N179 | ovr_btaken;
  assign N179 = linear_miss | ovr_ret;
  assign attaboy_yumi_o = N184 & N187;
  assign N184 = attaboy_v_i & N183;
  assign N183 = ~N182;
  assign N182 = bht_w_v_li & N181;
  assign N181 = ~bht_w_yumi_lo;
  assign N187 = ~N186;
  assign N186 = btb_w_v_li & N185;
  assign N185 = ~btb_w_yumi_lo;
  assign init_done_o = N188 & ras_init_done_lo;
  assign N188 = bht_init_done_lo & btb_init_done_lo;
  assign N141 = metadata_if1[48] & N189;
  assign N189 = ~ovr_o;
  assign N142 = redirect_br_v_i;
  assign N143 = N141 | N142;
  assign N144 = ~N143;
  assign N145 = ~N142;
  assign N146 = N141 & N145;
  assign ghistory_w_v = redirect_br_v_i | icache_tv_we_i;

endmodule



module bsg_dff_reset_en_width_p59
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [58:0] data_i;
  output [58:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [58:0] data_o;
  wire N0,N1,N2;
  reg data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,data_o_55_sv2v_reg,
  data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,data_o_51_sv2v_reg,
  data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,data_o_47_sv2v_reg,
  data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,data_o_43_sv2v_reg,
  data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,
  data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,
  data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,
  data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,
  data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,
  data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,
  data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,
  data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,
  data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_58_sv2v_reg <= 1'b0;
      data_o_57_sv2v_reg <= 1'b0;
      data_o_56_sv2v_reg <= 1'b0;
      data_o_55_sv2v_reg <= 1'b0;
      data_o_54_sv2v_reg <= 1'b0;
      data_o_53_sv2v_reg <= 1'b0;
      data_o_52_sv2v_reg <= 1'b0;
      data_o_51_sv2v_reg <= 1'b0;
      data_o_50_sv2v_reg <= 1'b0;
      data_o_49_sv2v_reg <= 1'b0;
      data_o_48_sv2v_reg <= 1'b0;
      data_o_47_sv2v_reg <= 1'b0;
      data_o_46_sv2v_reg <= 1'b0;
      data_o_45_sv2v_reg <= 1'b0;
      data_o_44_sv2v_reg <= 1'b0;
      data_o_43_sv2v_reg <= 1'b0;
      data_o_42_sv2v_reg <= 1'b0;
      data_o_41_sv2v_reg <= 1'b0;
      data_o_40_sv2v_reg <= 1'b0;
      data_o_39_sv2v_reg <= 1'b0;
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_rotate_left_width_p36
(
  data_i,
  rot_i,
  o
);

  input [35:0] data_i;
  input [5:0] rot_i;
  output [35:0] o;
  wire [35:0] o;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,
  sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,
  sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,sv2v_dc_21,sv2v_dc_22,
  sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,sv2v_dc_27,sv2v_dc_28,sv2v_dc_29,
  sv2v_dc_30,sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,sv2v_dc_34,sv2v_dc_35,sv2v_dc_36;
  assign { o, sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36 } = { data_i, data_i } << rot_i;

endmodule



module bsg_dff_en_0000001b
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [26:0] data_i;
  output [26:0] data_o;
  input clk_i;
  input en_i;
  wire [26:0] data_o;
  reg data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,
  data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,
  data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,
  data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_en_width_p1
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [0:0] data_o;
  wire N0,N1,N2;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_cam_1r1w_tag_array_0000001b_00000008
(
  clk_i,
  reset_i,
  w_v_i,
  w_set_not_clear_i,
  w_tag_i,
  w_empty_o,
  r_v_i,
  r_tag_i,
  r_match_o
);

  input [7:0] w_v_i;
  input [26:0] w_tag_i;
  output [7:0] w_empty_o;
  input [26:0] r_tag_i;
  output [7:0] r_match_o;
  input clk_i;
  input reset_i;
  input w_set_not_clear_i;
  input r_v_i;
  wire [7:0] w_empty_o,r_match_o,v_r;
  wire _0_net_,N0,_1_net_,N1,_2_net_,N2,_3_net_,N3,_4_net_,N4,_5_net_,N5,_6_net_,N6,
  _7_net_,N7,N8,N9,N10,N11,N12,N13,N14,N15;
  wire [215:0] tag_r;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_0_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[0]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[0])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_0_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_0_net_),
    .data_o(tag_r[26:0])
  );

  assign N0 = tag_r[26:0] == r_tag_i;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_1_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[1]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[1])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_1_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_1_net_),
    .data_o(tag_r[53:27])
  );

  assign N1 = tag_r[53:27] == r_tag_i;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_2_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[2]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[2])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_2_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_2_net_),
    .data_o(tag_r[80:54])
  );

  assign N2 = tag_r[80:54] == r_tag_i;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_3_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[3]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[3])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_3_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_3_net_),
    .data_o(tag_r[107:81])
  );

  assign N3 = tag_r[107:81] == r_tag_i;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_4_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[4]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[4])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_4_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_4_net_),
    .data_o(tag_r[134:108])
  );

  assign N4 = tag_r[134:108] == r_tag_i;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_5_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[5]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[5])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_5_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_5_net_),
    .data_o(tag_r[161:135])
  );

  assign N5 = tag_r[161:135] == r_tag_i;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_6_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[6]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[6])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_6_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_6_net_),
    .data_o(tag_r[188:162])
  );

  assign N6 = tag_r[188:162] == r_tag_i;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_7_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[7]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[7])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_7_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_7_net_),
    .data_o(tag_r[215:189])
  );

  assign N7 = tag_r[215:189] == r_tag_i;
  assign _0_net_ = w_v_i[0] & w_set_not_clear_i;
  assign r_match_o[0] = N8 & N0;
  assign N8 = r_v_i & v_r[0];
  assign w_empty_o[0] = ~v_r[0];
  assign _1_net_ = w_v_i[1] & w_set_not_clear_i;
  assign r_match_o[1] = N9 & N1;
  assign N9 = r_v_i & v_r[1];
  assign w_empty_o[1] = ~v_r[1];
  assign _2_net_ = w_v_i[2] & w_set_not_clear_i;
  assign r_match_o[2] = N10 & N2;
  assign N10 = r_v_i & v_r[2];
  assign w_empty_o[2] = ~v_r[2];
  assign _3_net_ = w_v_i[3] & w_set_not_clear_i;
  assign r_match_o[3] = N11 & N3;
  assign N11 = r_v_i & v_r[3];
  assign w_empty_o[3] = ~v_r[3];
  assign _4_net_ = w_v_i[4] & w_set_not_clear_i;
  assign r_match_o[4] = N12 & N4;
  assign N12 = r_v_i & v_r[4];
  assign w_empty_o[4] = ~v_r[4];
  assign _5_net_ = w_v_i[5] & w_set_not_clear_i;
  assign r_match_o[5] = N13 & N5;
  assign N13 = r_v_i & v_r[5];
  assign w_empty_o[5] = ~v_r[5];
  assign _6_net_ = w_v_i[6] & w_set_not_clear_i;
  assign r_match_o[6] = N14 & N6;
  assign N14 = r_v_i & v_r[6];
  assign w_empty_o[6] = ~v_r[6];
  assign _7_net_ = w_v_i[7] & w_set_not_clear_i;
  assign r_match_o[7] = N15 & N7;
  assign N15 = r_v_i & v_r[7];
  assign w_empty_o[7] = ~v_r[7];

endmodule



module bsg_dff_reset_en_00000007
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [6:0] data_i;
  output [6:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [6:0] data_o;
  wire N0,N1,N2;
  reg data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mux_width_p1_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [1:0] data_i;
  input [0:0] sel_i;
  output [0:0] data_o;
  wire [0:0] data_o;
  wire N0,N1;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[1] : 1'b0;
  assign N0 = sel_i[0];
  assign N1 = ~sel_i[0];

endmodule



module bsg_mux_width_p1_els_p4
(
  data_i,
  sel_i,
  data_o
);

  input [3:0] data_i;
  input [1:0] sel_i;
  output [0:0] data_o;
  wire [0:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[1] : 
                     (N3)? data_i[2] : 
                     (N5)? data_i[3] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_lru_pseudo_tree_encode_00000008
(
  lru_i,
  way_id_o
);

  input [6:0] lru_i;
  output [2:0] way_id_o;
  wire [2:0] way_id_o;
  wire way_id_o_2_;
  assign way_id_o_2_ = lru_i[0];
  assign way_id_o[2] = way_id_o_2_;

  bsg_mux_width_p1_els_p2
  \lru.rank_1_.nz.mux 
  (
    .data_i(lru_i[2:1]),
    .sel_i(way_id_o_2_),
    .data_o(way_id_o[1])
  );


  bsg_mux_width_p1_els_p4
  \lru.rank_2_.nz.mux 
  (
    .data_i(lru_i[6:3]),
    .sel_i({ way_id_o_2_, way_id_o[1:1] }),
    .data_o(way_id_o[0])
  );


endmodule



module bsg_scan_00000008_1_1
(
  i,
  o
);

  input [7:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__7_,t_1__6_,
  t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__7_ = i[0] | 1'b0;
  assign t_1__6_ = i[1] | i[0];
  assign t_1__5_ = i[2] | i[1];
  assign t_1__4_ = i[3] | i[2];
  assign t_1__3_ = i[4] | i[3];
  assign t_1__2_ = i[5] | i[4];
  assign t_1__1_ = i[6] | i[5];
  assign t_1__0_ = i[7] | i[6];
  assign t_2__7_ = t_1__7_ | 1'b0;
  assign t_2__6_ = t_1__6_ | 1'b0;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign o[0] = t_2__7_ | 1'b0;
  assign o[1] = t_2__6_ | 1'b0;
  assign o[2] = t_2__5_ | 1'b0;
  assign o[3] = t_2__4_ | 1'b0;
  assign o[4] = t_2__3_ | t_2__7_;
  assign o[5] = t_2__2_ | t_2__6_;
  assign o[6] = t_2__1_ | t_2__5_;
  assign o[7] = t_2__0_ | t_2__4_;

endmodule



module bsg_priority_encode_one_hot_out_00000008_1
(
  i,
  o,
  v_o
);

  input [7:0] i;
  output [7:0] o;
  output v_o;
  wire [7:0] o;
  wire v_o,N0,N1,N2,N3,N4,N5,N6;
  wire [6:1] scan_lo;

  bsg_scan_00000008_1_1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, scan_lo, o[0:0] })
  );

  assign o[7] = v_o & N0;
  assign N0 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N1;
  assign N1 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N2;
  assign N2 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N3;
  assign N3 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N4;
  assign N4 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N5;
  assign N5 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N6;
  assign N6 = ~o[0];

endmodule



module bsg_encode_one_hot_00000008_1
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o,v_2__0_,v_1__6_,v_1__4_,v_1__2_,v_1__0_,addr_2__4_,addr_2__0_;
  assign v_1__0_ = i[1] | i[0];
  assign v_1__2_ = i[3] | i[2];
  assign v_1__4_ = i[5] | i[4];
  assign v_1__6_ = i[7] | i[6];
  assign v_2__0_ = v_1__2_ | v_1__0_;
  assign addr_2__0_ = i[1] | i[3];
  assign addr_o[2] = v_1__6_ | v_1__4_;
  assign addr_2__4_ = i[5] | i[7];
  assign v_o = addr_o[2] | v_2__0_;
  assign addr_o[1] = v_1__2_ | v_1__6_;
  assign addr_o[0] = addr_2__0_ | addr_2__4_;

endmodule



module bsg_priority_encode_00000008_1
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [7:0] enc_lo;

  bsg_priority_encode_one_hot_out_00000008_1
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_00000008_1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o)
  );


endmodule



module bsg_decode_00000008
(
  i,
  o
);

  input [2:0] i;
  output [7:0] o;
  wire [7:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_encode_one_hot_00000008
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o,v_2__0_,v_1__6_,v_1__4_,v_1__2_,v_1__0_,addr_2__4_,addr_2__0_;
  assign v_1__0_ = i[1] | i[0];
  assign v_1__2_ = i[3] | i[2];
  assign v_1__4_ = i[5] | i[4];
  assign v_1__6_ = i[7] | i[6];
  assign v_2__0_ = v_1__2_ | v_1__0_;
  assign addr_2__0_ = i[1] | i[3];
  assign addr_o[2] = v_1__6_ | v_1__4_;
  assign addr_2__4_ = i[5] | i[7];
  assign v_o = addr_o[2] | v_2__0_;
  assign addr_o[1] = v_1__2_ | v_1__6_;
  assign addr_o[0] = addr_2__0_ | addr_2__4_;

endmodule



module bsg_lru_pseudo_tree_decode_00000008
(
  way_id_i,
  data_o,
  mask_o
);

  input [2:0] way_id_i;
  output [6:0] data_o;
  output [6:0] mask_o;
  wire [6:0] data_o,mask_o;
  wire N0,N1,N2;
  assign mask_o[0] = 1'b1;
  assign data_o[0] = 1'b1 & N0;
  assign N0 = ~way_id_i[2];
  assign mask_o[1] = 1'b1 & N0;
  assign data_o[1] = mask_o[1] & N1;
  assign N1 = ~way_id_i[1];
  assign mask_o[2] = 1'b1 & way_id_i[2];
  assign data_o[2] = mask_o[2] & N1;
  assign mask_o[3] = mask_o[1] & N1;
  assign data_o[3] = mask_o[3] & N2;
  assign N2 = ~way_id_i[0];
  assign mask_o[4] = mask_o[1] & way_id_i[1];
  assign data_o[4] = mask_o[4] & N2;
  assign mask_o[5] = mask_o[2] & N1;
  assign data_o[5] = mask_o[5] & N2;
  assign mask_o[6] = mask_o[2] & way_id_i[1];
  assign data_o[6] = mask_o[6] & N2;

endmodule



module bsg_mux_segmented_00000007_1
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [6:0] data0_i;
  input [6:0] data1_i;
  input [6:0] sel_i;
  output [6:0] data_o;
  wire [6:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;
  assign data_o[0] = (N0)? data1_i[0] : 
                     (N7)? data0_i[0] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[1] = (N1)? data1_i[1] : 
                     (N8)? data0_i[1] : 1'b0;
  assign N1 = sel_i[1];
  assign data_o[2] = (N2)? data1_i[2] : 
                     (N9)? data0_i[2] : 1'b0;
  assign N2 = sel_i[2];
  assign data_o[3] = (N3)? data1_i[3] : 
                     (N10)? data0_i[3] : 1'b0;
  assign N3 = sel_i[3];
  assign data_o[4] = (N4)? data1_i[4] : 
                     (N11)? data0_i[4] : 1'b0;
  assign N4 = sel_i[4];
  assign data_o[5] = (N5)? data1_i[5] : 
                     (N12)? data0_i[5] : 1'b0;
  assign N5 = sel_i[5];
  assign data_o[6] = (N6)? data1_i[6] : 
                     (N13)? data0_i[6] : 1'b0;
  assign N6 = sel_i[6];
  assign N7 = ~sel_i[0];
  assign N8 = ~sel_i[1];
  assign N9 = ~sel_i[2];
  assign N10 = ~sel_i[3];
  assign N11 = ~sel_i[4];
  assign N12 = ~sel_i[5];
  assign N13 = ~sel_i[6];

endmodule



module bsg_mux_bitwise_00000007
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [6:0] data0_i;
  input [6:0] data1_i;
  input [6:0] sel_i;
  output [6:0] data_o;
  wire [6:0] data_o;

  bsg_mux_segmented_00000007_1
  mux_segmented
  (
    .data0_i(data0_i),
    .data1_i(data1_i),
    .sel_i(sel_i),
    .data_o(data_o)
  );


endmodule



module bsg_cam_1r1w_replacement_00000008
(
  clk_i,
  reset_i,
  read_v_i,
  alloc_v_i,
  alloc_empty_i,
  alloc_v_o
);

  input [7:0] read_v_i;
  input [7:0] alloc_empty_i;
  output [7:0] alloc_v_o;
  input clk_i;
  input reset_i;
  input alloc_v_i;
  wire [7:0] alloc_v_o;
  wire N0,N1,\lru.read_v_li ,\lru.lru_touch_li ,\lru.empty_way_v_lo ,N2,N3,N4,N5,N6,N7,
  N8;
  wire [6:0] \lru.lru_r ,\lru.read_update_data_lo ,\lru.read_update_mask_lo ,
  \lru.read_sel_lo ,\lru.read_update_lo ,\lru.alloc_update_data_lo ,\lru.alloc_update_mask_lo ,
  \lru.alloc_sel_lo ,\lru.alloc_update_lo ;
  wire [2:0] \lru.lru_way_lo ,\lru.empty_way_lo ,\lru.way_lo ,\lru.read_way_li ;

  bsg_dff_reset_en_00000007
  \lru.lru_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(\lru.lru_touch_li ),
    .data_i(\lru.alloc_update_lo ),
    .data_o(\lru.lru_r )
  );


  bsg_lru_pseudo_tree_encode_00000008
  \lru.lru_encoder 
  (
    .lru_i(\lru.lru_r ),
    .way_id_o(\lru.lru_way_lo )
  );


  bsg_priority_encode_00000008_1
  \lru.empty_encoder 
  (
    .i(alloc_empty_i),
    .addr_o(\lru.empty_way_lo ),
    .v_o(\lru.empty_way_v_lo )
  );


  bsg_decode_00000008
  \lru.way_decoder 
  (
    .i(\lru.way_lo ),
    .o(alloc_v_o)
  );


  bsg_encode_one_hot_00000008
  \lru.read_way_encoder 
  (
    .i(read_v_i),
    .addr_o(\lru.read_way_li )
  );


  bsg_lru_pseudo_tree_decode_00000008
  \lru.read_decoder 
  (
    .way_id_i(\lru.read_way_li ),
    .data_o(\lru.read_update_data_lo ),
    .mask_o(\lru.read_update_mask_lo )
  );


  bsg_mux_bitwise_00000007
  \lru.read_update_mux 
  (
    .data0_i(\lru.lru_r ),
    .data1_i(\lru.read_update_data_lo ),
    .sel_i(\lru.read_sel_lo ),
    .data_o(\lru.read_update_lo )
  );


  bsg_lru_pseudo_tree_decode_00000008
  \lru.alloc_decoder 
  (
    .way_id_i(\lru.way_lo ),
    .data_o(\lru.alloc_update_data_lo ),
    .mask_o(\lru.alloc_update_mask_lo )
  );


  bsg_mux_bitwise_00000007
  \lru.alloc_update_mux 
  (
    .data0_i(\lru.read_update_lo ),
    .data1_i(\lru.alloc_update_data_lo ),
    .sel_i(\lru.alloc_sel_lo ),
    .data_o(\lru.alloc_update_lo )
  );

  assign \lru.way_lo  = (N0)? \lru.empty_way_lo  : 
                        (N1)? \lru.lru_way_lo  : 1'b0;
  assign N0 = \lru.empty_way_v_lo ;
  assign N1 = N2;
  assign \lru.read_v_li  = N8 | read_v_i[0];
  assign N8 = N7 | read_v_i[1];
  assign N7 = N6 | read_v_i[2];
  assign N6 = N5 | read_v_i[3];
  assign N5 = N4 | read_v_i[4];
  assign N4 = N3 | read_v_i[5];
  assign N3 = read_v_i[7] | read_v_i[6];
  assign \lru.lru_touch_li  = \lru.read_v_li  | alloc_v_i;
  assign N2 = ~\lru.empty_way_v_lo ;
  assign \lru.read_sel_lo [6] = \lru.read_update_mask_lo [6] & \lru.read_v_li ;
  assign \lru.read_sel_lo [5] = \lru.read_update_mask_lo [5] & \lru.read_v_li ;
  assign \lru.read_sel_lo [4] = \lru.read_update_mask_lo [4] & \lru.read_v_li ;
  assign \lru.read_sel_lo [3] = \lru.read_update_mask_lo [3] & \lru.read_v_li ;
  assign \lru.read_sel_lo [2] = \lru.read_update_mask_lo [2] & \lru.read_v_li ;
  assign \lru.read_sel_lo [1] = \lru.read_update_mask_lo [1] & \lru.read_v_li ;
  assign \lru.read_sel_lo [0] = \lru.read_update_mask_lo [0] & \lru.read_v_li ;
  assign \lru.alloc_sel_lo [6] = \lru.alloc_update_mask_lo [6] & alloc_v_i;
  assign \lru.alloc_sel_lo [5] = \lru.alloc_update_mask_lo [5] & alloc_v_i;
  assign \lru.alloc_sel_lo [4] = \lru.alloc_update_mask_lo [4] & alloc_v_i;
  assign \lru.alloc_sel_lo [3] = \lru.alloc_update_mask_lo [3] & alloc_v_i;
  assign \lru.alloc_sel_lo [2] = \lru.alloc_update_mask_lo [2] & alloc_v_i;
  assign \lru.alloc_sel_lo [1] = \lru.alloc_update_mask_lo [1] & alloc_v_i;
  assign \lru.alloc_sel_lo [0] = \lru.alloc_update_mask_lo [0] & alloc_v_i;

endmodule



module bsg_cam_1r1w_tag_array_0000001b_00000002
(
  clk_i,
  reset_i,
  w_v_i,
  w_set_not_clear_i,
  w_tag_i,
  w_empty_o,
  r_v_i,
  r_tag_i,
  r_match_o
);

  input [1:0] w_v_i;
  input [26:0] w_tag_i;
  output [1:0] w_empty_o;
  input [26:0] r_tag_i;
  output [1:0] r_match_o;
  input clk_i;
  input reset_i;
  input w_set_not_clear_i;
  input r_v_i;
  wire [1:0] w_empty_o,r_match_o,v_r;
  wire _0_net_,N0,_1_net_,N1,N2,N3;
  wire [53:0] tag_r;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_0_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[0]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[0])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_0_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_0_net_),
    .data_o(tag_r[26:0])
  );

  assign N0 = tag_r[26:0] == r_tag_i;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_1_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[1]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[1])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_1_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_1_net_),
    .data_o(tag_r[53:27])
  );

  assign N1 = tag_r[53:27] == r_tag_i;
  assign _0_net_ = w_v_i[0] & w_set_not_clear_i;
  assign r_match_o[0] = N2 & N0;
  assign N2 = r_v_i & v_r[0];
  assign w_empty_o[0] = ~v_r[0];
  assign _1_net_ = w_v_i[1] & w_set_not_clear_i;
  assign r_match_o[1] = N3 & N1;
  assign N3 = r_v_i & v_r[1];
  assign w_empty_o[1] = ~v_r[1];

endmodule



module bsg_lru_pseudo_tree_encode_00000002
(
  lru_i,
  way_id_o
);

  input [0:0] lru_i;
  output [0:0] way_id_o;
  wire [0:0] way_id_o;
  assign way_id_o[0] = lru_i[0];

endmodule



module bsg_scan_00000002_1_1
(
  i,
  o
);

  input [1:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o[0] = i[0] | 1'b0;
  assign o[1] = i[1] | i[0];

endmodule



module bsg_priority_encode_one_hot_out_00000002_1
(
  i,
  o,
  v_o
);

  input [1:0] i;
  output [1:0] o;
  output v_o;
  wire [1:0] o;
  wire v_o,N0;

  bsg_scan_00000002_1_1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, o[0:0] })
  );

  assign o[1] = v_o & N0;
  assign N0 = ~o[0];

endmodule



module bsg_encode_one_hot_00000002_1
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign addr_o[0] = i[1];
  assign v_o = addr_o[0] | i[0];

endmodule



module bsg_priority_encode_00000002_1
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  wire [1:0] enc_lo;

  bsg_priority_encode_one_hot_out_00000002_1
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_00000002_1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o[0])
  );


endmodule



module bsg_decode_00000002
(
  i,
  o
);

  input [0:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o = { 1'b0, 1'b1 } << i[0];

endmodule



module bsg_encode_one_hot_00000002
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign addr_o[0] = i[1];
  assign v_o = addr_o[0] | i[0];

endmodule



module bsg_lru_pseudo_tree_decode_00000002
(
  way_id_i,
  data_o,
  mask_o
);

  input [0:0] way_id_i;
  output [0:0] data_o;
  output [0:0] mask_o;
  wire [0:0] data_o,mask_o;
  wire N0;
  assign mask_o[0] = 1'b1;
  assign data_o[0] = 1'b1 & N0;
  assign N0 = ~way_id_i[0];

endmodule



module bsg_mux_segmented_00000001_1
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [0:0] data0_i;
  input [0:0] data1_i;
  input [0:0] sel_i;
  output [0:0] data_o;
  wire [0:0] data_o;
  wire N0,N1;
  assign data_o[0] = (N0)? data1_i[0] : 
                     (N1)? data0_i[0] : 1'b0;
  assign N0 = sel_i[0];
  assign N1 = ~sel_i[0];

endmodule



module bsg_mux_bitwise_00000001
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [0:0] data0_i;
  input [0:0] data1_i;
  input [0:0] sel_i;
  output [0:0] data_o;
  wire [0:0] data_o;

  bsg_mux_segmented_00000001_1
  mux_segmented
  (
    .data0_i(data0_i[0]),
    .data1_i(data1_i[0]),
    .sel_i(sel_i[0]),
    .data_o(data_o[0])
  );


endmodule



module bsg_cam_1r1w_replacement_00000002
(
  clk_i,
  reset_i,
  read_v_i,
  alloc_v_i,
  alloc_empty_i,
  alloc_v_o
);

  input [1:0] read_v_i;
  input [1:0] alloc_empty_i;
  output [1:0] alloc_v_o;
  input clk_i;
  input reset_i;
  input alloc_v_i;
  wire [1:0] alloc_v_o;
  wire N0,N1,\lru.read_v_li ,\lru.lru_touch_li ,\lru.empty_way_v_lo ,N2;
  wire [0:0] \lru.lru_r ,\lru.lru_way_lo ,\lru.empty_way_lo ,\lru.way_lo ,\lru.read_way_li ,
  \lru.read_update_data_lo ,\lru.read_update_mask_lo ,\lru.read_sel_lo ,
  \lru.read_update_lo ,\lru.alloc_update_data_lo ,\lru.alloc_update_mask_lo ,
  \lru.alloc_sel_lo ,\lru.alloc_update_lo ;

  bsg_dff_reset_en_width_p1
  \lru.lru_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(\lru.lru_touch_li ),
    .data_i(\lru.alloc_update_lo [0]),
    .data_o(\lru.lru_r [0])
  );


  bsg_lru_pseudo_tree_encode_00000002
  \lru.lru_encoder 
  (
    .lru_i(\lru.lru_r [0]),
    .way_id_o(\lru.lru_way_lo [0])
  );


  bsg_priority_encode_00000002_1
  \lru.empty_encoder 
  (
    .i(alloc_empty_i),
    .addr_o(\lru.empty_way_lo [0]),
    .v_o(\lru.empty_way_v_lo )
  );


  bsg_decode_00000002
  \lru.way_decoder 
  (
    .i(\lru.way_lo [0]),
    .o(alloc_v_o)
  );


  bsg_encode_one_hot_00000002
  \lru.read_way_encoder 
  (
    .i(read_v_i),
    .addr_o(\lru.read_way_li [0])
  );


  bsg_lru_pseudo_tree_decode_00000002
  \lru.read_decoder 
  (
    .way_id_i(\lru.read_way_li [0]),
    .data_o(\lru.read_update_data_lo [0]),
    .mask_o(\lru.read_update_mask_lo [0])
  );


  bsg_mux_bitwise_00000001
  \lru.read_update_mux 
  (
    .data0_i(\lru.lru_r [0]),
    .data1_i(\lru.read_update_data_lo [0]),
    .sel_i(\lru.read_sel_lo [0]),
    .data_o(\lru.read_update_lo [0])
  );


  bsg_lru_pseudo_tree_decode_00000002
  \lru.alloc_decoder 
  (
    .way_id_i(\lru.way_lo [0]),
    .data_o(\lru.alloc_update_data_lo [0]),
    .mask_o(\lru.alloc_update_mask_lo [0])
  );


  bsg_mux_bitwise_00000001
  \lru.alloc_update_mux 
  (
    .data0_i(\lru.read_update_lo [0]),
    .data1_i(\lru.alloc_update_data_lo [0]),
    .sel_i(\lru.alloc_sel_lo [0]),
    .data_o(\lru.alloc_update_lo [0])
  );

  assign \lru.way_lo [0] = (N0)? \lru.empty_way_lo [0] : 
                           (N1)? \lru.lru_way_lo [0] : 1'b0;
  assign N0 = \lru.empty_way_v_lo ;
  assign N1 = N2;
  assign \lru.read_v_li  = read_v_i[1] | read_v_i[0];
  assign \lru.lru_touch_li  = \lru.read_v_li  | alloc_v_i;
  assign N2 = ~\lru.empty_way_v_lo ;
  assign \lru.read_sel_lo [0] = \lru.read_update_mask_lo [0] & \lru.read_v_li ;
  assign \lru.alloc_sel_lo [0] = \lru.alloc_update_mask_lo [0] & alloc_v_i;

endmodule



module bsg_cam_1r1w_tag_array_0000001b_00000001
(
  clk_i,
  reset_i,
  w_v_i,
  w_set_not_clear_i,
  w_tag_i,
  w_empty_o,
  r_v_i,
  r_tag_i,
  r_match_o
);

  input [0:0] w_v_i;
  input [26:0] w_tag_i;
  output [0:0] w_empty_o;
  input [26:0] r_tag_i;
  output [0:0] r_match_o;
  input clk_i;
  input reset_i;
  input w_set_not_clear_i;
  input r_v_i;
  wire [0:0] w_empty_o,r_match_o,v_r;
  wire _0_net_,N0,N1;
  wire [26:0] tag_r;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_0_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[0]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[0])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_0_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_0_net_),
    .data_o(tag_r)
  );

  assign N0 = tag_r == r_tag_i;
  assign _0_net_ = w_v_i[0] & w_set_not_clear_i;
  assign r_match_o[0] = N1 & N0;
  assign N1 = r_v_i & v_r[0];
  assign w_empty_o[0] = ~v_r[0];

endmodule



module bsg_cam_1r1w_replacement_00000001
(
  clk_i,
  reset_i,
  read_v_i,
  alloc_v_i,
  alloc_empty_i,
  alloc_v_o
);

  input [0:0] read_v_i;
  input [0:0] alloc_empty_i;
  output [0:0] alloc_v_o;
  input clk_i;
  input reset_i;
  input alloc_v_i;
  wire [0:0] alloc_v_o;
  assign alloc_v_o[0] = 1'b1;

endmodule



module bsg_dff_en_00000024
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [35:0] data_i;
  output [35:0] data_o;
  input clk_i;
  input en_i;
  wire [35:0] data_o;
  reg data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,
  data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,
  data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,
  data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_width_p18
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [17:0] data_i;
  output [17:0] data_o;
  input clk_i;
  input en_i;
  wire [17:0] data_o;
  reg data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,
  data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mux_one_hot_9_00000009
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [80:0] data_i;
  input [8:0] sel_one_hot_i;
  output [8:0] data_o;
  wire [8:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62;
  wire [80:0] data_masked;
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[1];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[1];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[1];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[1];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[1];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[1];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[1];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[1];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[1];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[2];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[2];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[2];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[2];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[2];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[2];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[2];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[2];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[2];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[3];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[3];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[3];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[3];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[3];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[3];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[3];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[3];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[3];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[4];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[4];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[4];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[4];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[4];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[4];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[4];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[4];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[4];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[5];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[5];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[5];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[5];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[5];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[5];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[5];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[5];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[5];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[6];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[6];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[6];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[6];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[6];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[6];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[6];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[6];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[6];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[7];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[7];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[7];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[7];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[7];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[7];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[7];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[7];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[7];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[8];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[8];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[8];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[8];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[8];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[8];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[8];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[8];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[8];
  assign data_o[0] = N6 | data_masked[0];
  assign N6 = N5 | data_masked[9];
  assign N5 = N4 | data_masked[18];
  assign N4 = N3 | data_masked[27];
  assign N3 = N2 | data_masked[36];
  assign N2 = N1 | data_masked[45];
  assign N1 = N0 | data_masked[54];
  assign N0 = data_masked[72] | data_masked[63];
  assign data_o[1] = N13 | data_masked[1];
  assign N13 = N12 | data_masked[10];
  assign N12 = N11 | data_masked[19];
  assign N11 = N10 | data_masked[28];
  assign N10 = N9 | data_masked[37];
  assign N9 = N8 | data_masked[46];
  assign N8 = N7 | data_masked[55];
  assign N7 = data_masked[73] | data_masked[64];
  assign data_o[2] = N20 | data_masked[2];
  assign N20 = N19 | data_masked[11];
  assign N19 = N18 | data_masked[20];
  assign N18 = N17 | data_masked[29];
  assign N17 = N16 | data_masked[38];
  assign N16 = N15 | data_masked[47];
  assign N15 = N14 | data_masked[56];
  assign N14 = data_masked[74] | data_masked[65];
  assign data_o[3] = N27 | data_masked[3];
  assign N27 = N26 | data_masked[12];
  assign N26 = N25 | data_masked[21];
  assign N25 = N24 | data_masked[30];
  assign N24 = N23 | data_masked[39];
  assign N23 = N22 | data_masked[48];
  assign N22 = N21 | data_masked[57];
  assign N21 = data_masked[75] | data_masked[66];
  assign data_o[4] = N34 | data_masked[4];
  assign N34 = N33 | data_masked[13];
  assign N33 = N32 | data_masked[22];
  assign N32 = N31 | data_masked[31];
  assign N31 = N30 | data_masked[40];
  assign N30 = N29 | data_masked[49];
  assign N29 = N28 | data_masked[58];
  assign N28 = data_masked[76] | data_masked[67];
  assign data_o[5] = N41 | data_masked[5];
  assign N41 = N40 | data_masked[14];
  assign N40 = N39 | data_masked[23];
  assign N39 = N38 | data_masked[32];
  assign N38 = N37 | data_masked[41];
  assign N37 = N36 | data_masked[50];
  assign N36 = N35 | data_masked[59];
  assign N35 = data_masked[77] | data_masked[68];
  assign data_o[6] = N48 | data_masked[6];
  assign N48 = N47 | data_masked[15];
  assign N47 = N46 | data_masked[24];
  assign N46 = N45 | data_masked[33];
  assign N45 = N44 | data_masked[42];
  assign N44 = N43 | data_masked[51];
  assign N43 = N42 | data_masked[60];
  assign N42 = data_masked[78] | data_masked[69];
  assign data_o[7] = N55 | data_masked[7];
  assign N55 = N54 | data_masked[16];
  assign N54 = N53 | data_masked[25];
  assign N53 = N52 | data_masked[34];
  assign N52 = N51 | data_masked[43];
  assign N51 = N50 | data_masked[52];
  assign N50 = N49 | data_masked[61];
  assign N49 = data_masked[79] | data_masked[70];
  assign data_o[8] = N62 | data_masked[8];
  assign N62 = N61 | data_masked[17];
  assign N61 = N60 | data_masked[26];
  assign N60 = N59 | data_masked[35];
  assign N59 = N58 | data_masked[44];
  assign N58 = N57 | data_masked[53];
  assign N57 = N56 | data_masked[62];
  assign N56 = data_masked[80] | data_masked[71];

endmodule



module bsg_mux_one_hot_9_0000000b
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [98:0] data_i;
  input [10:0] sel_one_hot_i;
  output [8:0] data_o;
  wire [8:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80;
  wire [98:0] data_masked;
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[1];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[1];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[1];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[1];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[1];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[1];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[1];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[1];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[1];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[2];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[2];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[2];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[2];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[2];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[2];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[2];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[2];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[2];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[3];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[3];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[3];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[3];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[3];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[3];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[3];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[3];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[3];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[4];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[4];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[4];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[4];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[4];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[4];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[4];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[4];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[4];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[5];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[5];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[5];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[5];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[5];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[5];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[5];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[5];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[5];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[6];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[6];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[6];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[6];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[6];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[6];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[6];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[6];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[6];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[7];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[7];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[7];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[7];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[7];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[7];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[7];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[7];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[7];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[8];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[8];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[8];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[8];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[8];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[8];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[8];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[8];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[8];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[9];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[9];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[9];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[9];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[9];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[9];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[9];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[9];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[9];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[10];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[10];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[10];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[10];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[10];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[10];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[10];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[10];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[10];
  assign data_o[0] = N8 | data_masked[0];
  assign N8 = N7 | data_masked[9];
  assign N7 = N6 | data_masked[18];
  assign N6 = N5 | data_masked[27];
  assign N5 = N4 | data_masked[36];
  assign N4 = N3 | data_masked[45];
  assign N3 = N2 | data_masked[54];
  assign N2 = N1 | data_masked[63];
  assign N1 = N0 | data_masked[72];
  assign N0 = data_masked[90] | data_masked[81];
  assign data_o[1] = N17 | data_masked[1];
  assign N17 = N16 | data_masked[10];
  assign N16 = N15 | data_masked[19];
  assign N15 = N14 | data_masked[28];
  assign N14 = N13 | data_masked[37];
  assign N13 = N12 | data_masked[46];
  assign N12 = N11 | data_masked[55];
  assign N11 = N10 | data_masked[64];
  assign N10 = N9 | data_masked[73];
  assign N9 = data_masked[91] | data_masked[82];
  assign data_o[2] = N26 | data_masked[2];
  assign N26 = N25 | data_masked[11];
  assign N25 = N24 | data_masked[20];
  assign N24 = N23 | data_masked[29];
  assign N23 = N22 | data_masked[38];
  assign N22 = N21 | data_masked[47];
  assign N21 = N20 | data_masked[56];
  assign N20 = N19 | data_masked[65];
  assign N19 = N18 | data_masked[74];
  assign N18 = data_masked[92] | data_masked[83];
  assign data_o[3] = N35 | data_masked[3];
  assign N35 = N34 | data_masked[12];
  assign N34 = N33 | data_masked[21];
  assign N33 = N32 | data_masked[30];
  assign N32 = N31 | data_masked[39];
  assign N31 = N30 | data_masked[48];
  assign N30 = N29 | data_masked[57];
  assign N29 = N28 | data_masked[66];
  assign N28 = N27 | data_masked[75];
  assign N27 = data_masked[93] | data_masked[84];
  assign data_o[4] = N44 | data_masked[4];
  assign N44 = N43 | data_masked[13];
  assign N43 = N42 | data_masked[22];
  assign N42 = N41 | data_masked[31];
  assign N41 = N40 | data_masked[40];
  assign N40 = N39 | data_masked[49];
  assign N39 = N38 | data_masked[58];
  assign N38 = N37 | data_masked[67];
  assign N37 = N36 | data_masked[76];
  assign N36 = data_masked[94] | data_masked[85];
  assign data_o[5] = N53 | data_masked[5];
  assign N53 = N52 | data_masked[14];
  assign N52 = N51 | data_masked[23];
  assign N51 = N50 | data_masked[32];
  assign N50 = N49 | data_masked[41];
  assign N49 = N48 | data_masked[50];
  assign N48 = N47 | data_masked[59];
  assign N47 = N46 | data_masked[68];
  assign N46 = N45 | data_masked[77];
  assign N45 = data_masked[95] | data_masked[86];
  assign data_o[6] = N62 | data_masked[6];
  assign N62 = N61 | data_masked[15];
  assign N61 = N60 | data_masked[24];
  assign N60 = N59 | data_masked[33];
  assign N59 = N58 | data_masked[42];
  assign N58 = N57 | data_masked[51];
  assign N57 = N56 | data_masked[60];
  assign N56 = N55 | data_masked[69];
  assign N55 = N54 | data_masked[78];
  assign N54 = data_masked[96] | data_masked[87];
  assign data_o[7] = N71 | data_masked[7];
  assign N71 = N70 | data_masked[16];
  assign N70 = N69 | data_masked[25];
  assign N69 = N68 | data_masked[34];
  assign N68 = N67 | data_masked[43];
  assign N67 = N66 | data_masked[52];
  assign N66 = N65 | data_masked[61];
  assign N65 = N64 | data_masked[70];
  assign N64 = N63 | data_masked[79];
  assign N63 = data_masked[97] | data_masked[88];
  assign data_o[8] = N80 | data_masked[8];
  assign N80 = N79 | data_masked[17];
  assign N79 = N78 | data_masked[26];
  assign N78 = N77 | data_masked[35];
  assign N77 = N76 | data_masked[44];
  assign N76 = N75 | data_masked[53];
  assign N75 = N74 | data_masked[62];
  assign N74 = N73 | data_masked[71];
  assign N73 = N72 | data_masked[80];
  assign N72 = data_masked[98] | data_masked[89];

endmodule



module bsg_mux_one_hot_18_0000000b
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [197:0] data_i;
  input [10:0] sel_one_hot_i;
  output [17:0] data_o;
  wire [17:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161;
  wire [197:0] data_masked;
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[1];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[1];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[1];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[1];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[1];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[1];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[1];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[1];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[1];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[1];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[1];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[1];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[1];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[1];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[1];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[1];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[1];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[1];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[2];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[2];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[2];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[2];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[2];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[2];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[2];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[2];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[2];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[2];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[2];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[2];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[2];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[2];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[2];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[2];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[2];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[2];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[3];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[3];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[3];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[3];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[3];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[3];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[3];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[3];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[3];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[3];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[3];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[3];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[3];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[3];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[3];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[3];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[3];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[3];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[4];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[4];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[4];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[4];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[4];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[4];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[4];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[4];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[4];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[4];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[4];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[4];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[4];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[4];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[4];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[4];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[4];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[4];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[5];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[5];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[5];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[5];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[5];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[5];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[5];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[5];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[5];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[5];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[5];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[5];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[5];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[5];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[5];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[5];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[5];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[5];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[6];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[6];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[6];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[6];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[6];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[6];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[6];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[6];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[6];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[6];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[6];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[6];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[6];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[6];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[6];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[6];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[6];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[6];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[7];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[7];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[7];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[7];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[7];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[7];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[7];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[7];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[7];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[7];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[7];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[7];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[7];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[7];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[7];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[7];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[7];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[7];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[8];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[8];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[8];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[8];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[8];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[8];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[8];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[8];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[8];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[8];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[8];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[8];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[8];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[8];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[8];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[8];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[8];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[8];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[9];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[9];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[9];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[9];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[9];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[9];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[9];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[9];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[9];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[9];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[9];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[9];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[9];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[9];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[9];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[9];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[9];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[9];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[10];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[10];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[10];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[10];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[10];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[10];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[10];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[10];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[10];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[10];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[10];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[10];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[10];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[10];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[10];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[10];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[10];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[10];
  assign data_o[0] = N8 | data_masked[0];
  assign N8 = N7 | data_masked[18];
  assign N7 = N6 | data_masked[36];
  assign N6 = N5 | data_masked[54];
  assign N5 = N4 | data_masked[72];
  assign N4 = N3 | data_masked[90];
  assign N3 = N2 | data_masked[108];
  assign N2 = N1 | data_masked[126];
  assign N1 = N0 | data_masked[144];
  assign N0 = data_masked[180] | data_masked[162];
  assign data_o[1] = N17 | data_masked[1];
  assign N17 = N16 | data_masked[19];
  assign N16 = N15 | data_masked[37];
  assign N15 = N14 | data_masked[55];
  assign N14 = N13 | data_masked[73];
  assign N13 = N12 | data_masked[91];
  assign N12 = N11 | data_masked[109];
  assign N11 = N10 | data_masked[127];
  assign N10 = N9 | data_masked[145];
  assign N9 = data_masked[181] | data_masked[163];
  assign data_o[2] = N26 | data_masked[2];
  assign N26 = N25 | data_masked[20];
  assign N25 = N24 | data_masked[38];
  assign N24 = N23 | data_masked[56];
  assign N23 = N22 | data_masked[74];
  assign N22 = N21 | data_masked[92];
  assign N21 = N20 | data_masked[110];
  assign N20 = N19 | data_masked[128];
  assign N19 = N18 | data_masked[146];
  assign N18 = data_masked[182] | data_masked[164];
  assign data_o[3] = N35 | data_masked[3];
  assign N35 = N34 | data_masked[21];
  assign N34 = N33 | data_masked[39];
  assign N33 = N32 | data_masked[57];
  assign N32 = N31 | data_masked[75];
  assign N31 = N30 | data_masked[93];
  assign N30 = N29 | data_masked[111];
  assign N29 = N28 | data_masked[129];
  assign N28 = N27 | data_masked[147];
  assign N27 = data_masked[183] | data_masked[165];
  assign data_o[4] = N44 | data_masked[4];
  assign N44 = N43 | data_masked[22];
  assign N43 = N42 | data_masked[40];
  assign N42 = N41 | data_masked[58];
  assign N41 = N40 | data_masked[76];
  assign N40 = N39 | data_masked[94];
  assign N39 = N38 | data_masked[112];
  assign N38 = N37 | data_masked[130];
  assign N37 = N36 | data_masked[148];
  assign N36 = data_masked[184] | data_masked[166];
  assign data_o[5] = N53 | data_masked[5];
  assign N53 = N52 | data_masked[23];
  assign N52 = N51 | data_masked[41];
  assign N51 = N50 | data_masked[59];
  assign N50 = N49 | data_masked[77];
  assign N49 = N48 | data_masked[95];
  assign N48 = N47 | data_masked[113];
  assign N47 = N46 | data_masked[131];
  assign N46 = N45 | data_masked[149];
  assign N45 = data_masked[185] | data_masked[167];
  assign data_o[6] = N62 | data_masked[6];
  assign N62 = N61 | data_masked[24];
  assign N61 = N60 | data_masked[42];
  assign N60 = N59 | data_masked[60];
  assign N59 = N58 | data_masked[78];
  assign N58 = N57 | data_masked[96];
  assign N57 = N56 | data_masked[114];
  assign N56 = N55 | data_masked[132];
  assign N55 = N54 | data_masked[150];
  assign N54 = data_masked[186] | data_masked[168];
  assign data_o[7] = N71 | data_masked[7];
  assign N71 = N70 | data_masked[25];
  assign N70 = N69 | data_masked[43];
  assign N69 = N68 | data_masked[61];
  assign N68 = N67 | data_masked[79];
  assign N67 = N66 | data_masked[97];
  assign N66 = N65 | data_masked[115];
  assign N65 = N64 | data_masked[133];
  assign N64 = N63 | data_masked[151];
  assign N63 = data_masked[187] | data_masked[169];
  assign data_o[8] = N80 | data_masked[8];
  assign N80 = N79 | data_masked[26];
  assign N79 = N78 | data_masked[44];
  assign N78 = N77 | data_masked[62];
  assign N77 = N76 | data_masked[80];
  assign N76 = N75 | data_masked[98];
  assign N75 = N74 | data_masked[116];
  assign N74 = N73 | data_masked[134];
  assign N73 = N72 | data_masked[152];
  assign N72 = data_masked[188] | data_masked[170];
  assign data_o[9] = N89 | data_masked[9];
  assign N89 = N88 | data_masked[27];
  assign N88 = N87 | data_masked[45];
  assign N87 = N86 | data_masked[63];
  assign N86 = N85 | data_masked[81];
  assign N85 = N84 | data_masked[99];
  assign N84 = N83 | data_masked[117];
  assign N83 = N82 | data_masked[135];
  assign N82 = N81 | data_masked[153];
  assign N81 = data_masked[189] | data_masked[171];
  assign data_o[10] = N98 | data_masked[10];
  assign N98 = N97 | data_masked[28];
  assign N97 = N96 | data_masked[46];
  assign N96 = N95 | data_masked[64];
  assign N95 = N94 | data_masked[82];
  assign N94 = N93 | data_masked[100];
  assign N93 = N92 | data_masked[118];
  assign N92 = N91 | data_masked[136];
  assign N91 = N90 | data_masked[154];
  assign N90 = data_masked[190] | data_masked[172];
  assign data_o[11] = N107 | data_masked[11];
  assign N107 = N106 | data_masked[29];
  assign N106 = N105 | data_masked[47];
  assign N105 = N104 | data_masked[65];
  assign N104 = N103 | data_masked[83];
  assign N103 = N102 | data_masked[101];
  assign N102 = N101 | data_masked[119];
  assign N101 = N100 | data_masked[137];
  assign N100 = N99 | data_masked[155];
  assign N99 = data_masked[191] | data_masked[173];
  assign data_o[12] = N116 | data_masked[12];
  assign N116 = N115 | data_masked[30];
  assign N115 = N114 | data_masked[48];
  assign N114 = N113 | data_masked[66];
  assign N113 = N112 | data_masked[84];
  assign N112 = N111 | data_masked[102];
  assign N111 = N110 | data_masked[120];
  assign N110 = N109 | data_masked[138];
  assign N109 = N108 | data_masked[156];
  assign N108 = data_masked[192] | data_masked[174];
  assign data_o[13] = N125 | data_masked[13];
  assign N125 = N124 | data_masked[31];
  assign N124 = N123 | data_masked[49];
  assign N123 = N122 | data_masked[67];
  assign N122 = N121 | data_masked[85];
  assign N121 = N120 | data_masked[103];
  assign N120 = N119 | data_masked[121];
  assign N119 = N118 | data_masked[139];
  assign N118 = N117 | data_masked[157];
  assign N117 = data_masked[193] | data_masked[175];
  assign data_o[14] = N134 | data_masked[14];
  assign N134 = N133 | data_masked[32];
  assign N133 = N132 | data_masked[50];
  assign N132 = N131 | data_masked[68];
  assign N131 = N130 | data_masked[86];
  assign N130 = N129 | data_masked[104];
  assign N129 = N128 | data_masked[122];
  assign N128 = N127 | data_masked[140];
  assign N127 = N126 | data_masked[158];
  assign N126 = data_masked[194] | data_masked[176];
  assign data_o[15] = N143 | data_masked[15];
  assign N143 = N142 | data_masked[33];
  assign N142 = N141 | data_masked[51];
  assign N141 = N140 | data_masked[69];
  assign N140 = N139 | data_masked[87];
  assign N139 = N138 | data_masked[105];
  assign N138 = N137 | data_masked[123];
  assign N137 = N136 | data_masked[141];
  assign N136 = N135 | data_masked[159];
  assign N135 = data_masked[195] | data_masked[177];
  assign data_o[16] = N152 | data_masked[16];
  assign N152 = N151 | data_masked[34];
  assign N151 = N150 | data_masked[52];
  assign N150 = N149 | data_masked[70];
  assign N149 = N148 | data_masked[88];
  assign N148 = N147 | data_masked[106];
  assign N147 = N146 | data_masked[124];
  assign N146 = N145 | data_masked[142];
  assign N145 = N144 | data_masked[160];
  assign N144 = data_masked[196] | data_masked[178];
  assign data_o[17] = N161 | data_masked[17];
  assign N161 = N160 | data_masked[35];
  assign N160 = N159 | data_masked[53];
  assign N159 = N158 | data_masked[71];
  assign N158 = N157 | data_masked[89];
  assign N157 = N156 | data_masked[107];
  assign N156 = N155 | data_masked[125];
  assign N155 = N154 | data_masked[143];
  assign N154 = N153 | data_masked[161];
  assign N153 = data_masked[197] | data_masked[179];

endmodule



module bsg_popcount_width_p3
(
  i,
  o
);

  input [2:0] i;
  output [1:0] o;
  wire [1:0] o;
  wire N0,N1,N2,N3,N4;
  assign o[0] = N0 ^ i[0];
  assign N0 = i[2] ^ i[1];
  assign o[1] = N3 | N4;
  assign N3 = N1 | N2;
  assign N1 = i[1] & i[0];
  assign N2 = i[2] & i[1];
  assign N4 = i[0] & i[2];

endmodule



module bsg_rotate_right_width_p36
(
  data_i,
  rot_i,
  o
);

  input [35:0] data_i;
  input [5:0] rot_i;
  output [35:0] o;
  wire [35:0] o;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,
  sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,
  sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,sv2v_dc_21,sv2v_dc_22,
  sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,sv2v_dc_27,sv2v_dc_28,sv2v_dc_29,
  sv2v_dc_30,sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,sv2v_dc_34,sv2v_dc_35,sv2v_dc_36;
  assign { sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36, o } = { data_i, data_i } >> rot_i;

endmodule



module bp_tlb_00_00000001_00000002_00000008
(
  clk_i,
  reset_i,
  fence_i,
  v_i,
  w_i,
  vtag_i,
  entry_i,
  v_o,
  entry_o
);

  input [26:0] vtag_i;
  input [35:0] entry_i;
  output [35:0] entry_o;
  input clk_i;
  input reset_i;
  input fence_i;
  input v_i;
  input w_i;
  output v_o;
  wire [35:0] entry_o,entry_shifted,data_2m_high_r,r_entry;
  wire v_o,w_v_li,fill_gigapage,fill_megapage,fill_kilopage,flush_4k_li,_1_net_,
  any_match_4k_lo,flush_2m_li,_3_net_,any_match_2m_lo,_5_net_,_21_net__8_,N0,N1,N3,N4,N5,
  N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26;
  wire [26:0] vtag_r;
  wire [7:0] repl_way_4k_lo,tag_4k_w_v_li,tag_empty_4k_lo,tag_r_match_4k_lo,mem_4k_w_v_li;
  wire [1:0] repl_way_2m_lo,tag_2m_w_v_li,tag_empty_2m_lo,tag_r_match_2m_lo,mem_2m_w_v_li,
  match_cnt;
  wire [0:0] repl_way_1g_lo,tag_1g_w_v_li,tag_empty_1g_lo,tag_r_match_1g_lo,mem_1g_w_v_li;
  wire [143:0] data_4k_high_r;
  wire [71:0] data_4k_med_r,data_4k_low_r;
  wire [17:0] data_2m_med_r,data_1g_high_r;

  bsg_rotate_left_width_p36
  entry_shift
  (
    .data_i(entry_i),
    .rot_i({ 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0 }),
    .o(entry_shifted)
  );


  bsg_dff_en_0000001b
  vtag_reg
  (
    .clk_i(clk_i),
    .data_i(vtag_i),
    .en_i(v_i),
    .data_o(vtag_r)
  );


  bsg_cam_1r1w_tag_array_0000001b_00000008
  tag_array_4k
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(tag_4k_w_v_li),
    .w_set_not_clear_i(_1_net_),
    .w_tag_i(vtag_i),
    .w_empty_o(tag_empty_4k_lo),
    .r_v_i(1'b1),
    .r_tag_i(vtag_r),
    .r_match_o(tag_r_match_4k_lo)
  );


  bsg_cam_1r1w_replacement_00000008
  replacement_4k
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .read_v_i(tag_r_match_4k_lo),
    .alloc_v_i(fill_kilopage),
    .alloc_empty_i(tag_empty_4k_lo),
    .alloc_v_o(repl_way_4k_lo)
  );


  bsg_cam_1r1w_tag_array_0000001b_00000002
  tag_array_2m
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(tag_2m_w_v_li),
    .w_set_not_clear_i(_3_net_),
    .w_tag_i(vtag_i),
    .w_empty_o(tag_empty_2m_lo),
    .r_v_i(1'b1),
    .r_tag_i(vtag_r),
    .r_match_o(tag_r_match_2m_lo)
  );


  bsg_cam_1r1w_replacement_00000002
  replacement_2m
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .read_v_i(tag_r_match_2m_lo),
    .alloc_v_i(fill_megapage),
    .alloc_empty_i(tag_empty_2m_lo),
    .alloc_v_o(repl_way_2m_lo)
  );


  bsg_cam_1r1w_tag_array_0000001b_00000001
  tag_array_1g
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(tag_1g_w_v_li[0]),
    .w_set_not_clear_i(_5_net_),
    .w_tag_i(vtag_i),
    .w_empty_o(tag_empty_1g_lo[0]),
    .r_v_i(1'b1),
    .r_tag_i(vtag_r),
    .r_match_o(tag_r_match_1g_lo[0])
  );


  bsg_cam_1r1w_replacement_00000001
  replacement_1g
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .read_v_i(tag_r_match_1g_lo[0]),
    .alloc_v_i(fill_gigapage),
    .alloc_empty_i(tag_empty_1g_lo[0]),
    .alloc_v_o(repl_way_1g_lo[0])
  );


  bsg_dff_en_00000024
  \mem_array_4k_0_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted),
    .en_i(mem_4k_w_v_li[0]),
    .data_o({ data_4k_high_r[17:0], data_4k_med_r[8:0], data_4k_low_r[8:0] })
  );


  bsg_dff_en_00000024
  \mem_array_4k_1_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted),
    .en_i(mem_4k_w_v_li[1]),
    .data_o({ data_4k_high_r[35:18], data_4k_med_r[17:9], data_4k_low_r[17:9] })
  );


  bsg_dff_en_00000024
  \mem_array_4k_2_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted),
    .en_i(mem_4k_w_v_li[2]),
    .data_o({ data_4k_high_r[53:36], data_4k_med_r[26:18], data_4k_low_r[26:18] })
  );


  bsg_dff_en_00000024
  \mem_array_4k_3_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted),
    .en_i(mem_4k_w_v_li[3]),
    .data_o({ data_4k_high_r[71:54], data_4k_med_r[35:27], data_4k_low_r[35:27] })
  );


  bsg_dff_en_00000024
  \mem_array_4k_4_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted),
    .en_i(mem_4k_w_v_li[4]),
    .data_o({ data_4k_high_r[89:72], data_4k_med_r[44:36], data_4k_low_r[44:36] })
  );


  bsg_dff_en_00000024
  \mem_array_4k_5_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted),
    .en_i(mem_4k_w_v_li[5]),
    .data_o({ data_4k_high_r[107:90], data_4k_med_r[53:45], data_4k_low_r[53:45] })
  );


  bsg_dff_en_00000024
  \mem_array_4k_6_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted),
    .en_i(mem_4k_w_v_li[6]),
    .data_o({ data_4k_high_r[125:108], data_4k_med_r[62:54], data_4k_low_r[62:54] })
  );


  bsg_dff_en_00000024
  \mem_array_4k_7_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted),
    .en_i(mem_4k_w_v_li[7]),
    .data_o({ data_4k_high_r[143:126], data_4k_med_r[71:63], data_4k_low_r[71:63] })
  );


  bsg_dff_en_0000001b
  \genblk2.mem_array_2m_0_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted[35:9]),
    .en_i(mem_2m_w_v_li[0]),
    .data_o({ data_2m_high_r[17:0], data_2m_med_r[8:0] })
  );


  bsg_dff_en_0000001b
  \genblk2.mem_array_2m_1_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted[35:9]),
    .en_i(mem_2m_w_v_li[1]),
    .data_o({ data_2m_high_r[35:18], data_2m_med_r[17:9] })
  );


  bsg_dff_en_width_p18
  \genblk3.mem_array_1g_0_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted[35:18]),
    .en_i(mem_1g_w_v_li[0]),
    .data_o(data_1g_high_r)
  );


  bsg_mux_one_hot_9_00000009
  one_hot_sel_low
  (
    .data_i({ vtag_r[8:0], data_4k_low_r }),
    .sel_one_hot_i({ _21_net__8_, tag_r_match_4k_lo }),
    .data_o(r_entry[8:0])
  );


  bsg_mux_one_hot_9_0000000b
  one_hot_sel_med
  (
    .data_i({ vtag_r[17:9], data_2m_med_r, data_4k_med_r }),
    .sel_one_hot_i({ tag_r_match_1g_lo[0:0], tag_r_match_2m_lo, tag_r_match_4k_lo }),
    .data_o(r_entry[17:9])
  );


  bsg_mux_one_hot_18_0000000b
  one_hot_sel_high
  (
    .data_i({ data_1g_high_r, data_2m_high_r, data_4k_high_r }),
    .sel_one_hot_i({ tag_r_match_1g_lo[0:0], tag_r_match_2m_lo, tag_r_match_4k_lo }),
    .data_o(r_entry[35:18])
  );


  bsg_popcount_width_p3
  mpc
  (
    .i({ tag_r_match_1g_lo[0:0], any_match_2m_lo, any_match_4k_lo }),
    .o(match_cnt)
  );


  bsg_rotate_right_width_p36
  entry_unshift
  (
    .data_i(r_entry),
    .rot_i({ 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0 }),
    .o(entry_o)
  );

  assign N0 = ~match_cnt[0];
  assign N1 = N0 | match_cnt[1];
  assign v_o = ~N1;
  assign w_v_li = v_i & w_i;
  assign fill_gigapage = w_v_li & entry_i[7];
  assign fill_megapage = w_v_li & entry_i[6];
  assign fill_kilopage = N4 & N5;
  assign N4 = w_v_li & N3;
  assign N3 = ~fill_gigapage;
  assign N5 = ~fill_megapage;
  assign tag_4k_w_v_li[7] = N6 | flush_4k_li;
  assign N6 = fill_kilopage & repl_way_4k_lo[7];
  assign tag_4k_w_v_li[6] = N7 | flush_4k_li;
  assign N7 = fill_kilopage & repl_way_4k_lo[6];
  assign tag_4k_w_v_li[5] = N8 | flush_4k_li;
  assign N8 = fill_kilopage & repl_way_4k_lo[5];
  assign tag_4k_w_v_li[4] = N9 | flush_4k_li;
  assign N9 = fill_kilopage & repl_way_4k_lo[4];
  assign tag_4k_w_v_li[3] = N10 | flush_4k_li;
  assign N10 = fill_kilopage & repl_way_4k_lo[3];
  assign tag_4k_w_v_li[2] = N11 | flush_4k_li;
  assign N11 = fill_kilopage & repl_way_4k_lo[2];
  assign tag_4k_w_v_li[1] = N12 | flush_4k_li;
  assign N12 = fill_kilopage & repl_way_4k_lo[1];
  assign tag_4k_w_v_li[0] = N13 | flush_4k_li;
  assign N13 = fill_kilopage & repl_way_4k_lo[0];
  assign _1_net_ = ~flush_4k_li;
  assign any_match_4k_lo = N19 | tag_r_match_4k_lo[0];
  assign N19 = N18 | tag_r_match_4k_lo[1];
  assign N18 = N17 | tag_r_match_4k_lo[2];
  assign N17 = N16 | tag_r_match_4k_lo[3];
  assign N16 = N15 | tag_r_match_4k_lo[4];
  assign N15 = N14 | tag_r_match_4k_lo[5];
  assign N14 = tag_r_match_4k_lo[7] | tag_r_match_4k_lo[6];
  assign tag_2m_w_v_li[1] = N20 | flush_2m_li;
  assign N20 = fill_megapage & repl_way_2m_lo[1];
  assign tag_2m_w_v_li[0] = N21 | flush_2m_li;
  assign N21 = fill_megapage & repl_way_2m_lo[0];
  assign _3_net_ = ~flush_2m_li;
  assign any_match_2m_lo = tag_r_match_2m_lo[1] | tag_r_match_2m_lo[0];
  assign tag_1g_w_v_li[0] = N22 | fence_i;
  assign N22 = fill_gigapage & repl_way_1g_lo[0];
  assign _5_net_ = ~fence_i;
  assign mem_4k_w_v_li[7] = fill_kilopage & repl_way_4k_lo[7];
  assign mem_4k_w_v_li[6] = fill_kilopage & repl_way_4k_lo[6];
  assign mem_4k_w_v_li[5] = fill_kilopage & repl_way_4k_lo[5];
  assign mem_4k_w_v_li[4] = fill_kilopage & repl_way_4k_lo[4];
  assign mem_4k_w_v_li[3] = fill_kilopage & repl_way_4k_lo[3];
  assign mem_4k_w_v_li[2] = fill_kilopage & repl_way_4k_lo[2];
  assign mem_4k_w_v_li[1] = fill_kilopage & repl_way_4k_lo[1];
  assign mem_4k_w_v_li[0] = fill_kilopage & repl_way_4k_lo[0];
  assign mem_2m_w_v_li[1] = fill_megapage & repl_way_2m_lo[1];
  assign mem_2m_w_v_li[0] = fill_megapage & repl_way_2m_lo[0];
  assign mem_1g_w_v_li[0] = fill_gigapage & repl_way_1g_lo[0];
  assign _21_net__8_ = tag_r_match_1g_lo[0] | any_match_2m_lo;
  assign flush_4k_li = N24 | N25;
  assign N24 = fence_i | N23;
  assign N23 = tag_r_match_1g_lo[0] & any_match_4k_lo;
  assign N25 = any_match_2m_lo & any_match_4k_lo;
  assign flush_2m_li = fence_i | N26;
  assign N26 = tag_r_match_1g_lo[0] & any_match_2m_lo;

endmodule



module bsg_dff_width_p1
(
  clk_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  wire [0:0] data_o;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_width_p37_harden_p0_strength_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [36:0] data_i;
  output [36:0] data_o;
  input clk_i;
  input en_i;
  wire [36:0] data_o;
  reg data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,
  data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,
  data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,
  data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,
  data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,
  data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,
  data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,
  data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_bypass_width_p37
(
  clk_i,
  en_i,
  data_i,
  data_o
);

  input [36:0] data_i;
  output [36:0] data_o;
  input clk_i;
  input en_i;
  wire [36:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_en_width_p37_harden_p0_strength_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(en_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_dff_sync_read_width_p37_bypass_p1
(
  clk_i,
  reset_i,
  v_n_i,
  data_i,
  data_o
);

  input [36:0] data_i;
  output [36:0] data_o;
  input clk_i;
  input reset_i;
  input v_n_i;
  wire [36:0] data_o;
  wire v_r;

  bsg_dff_width_p1
  v_reg
  (
    .clk_i(clk_i),
    .data_i(v_n_i),
    .data_o(v_r)
  );


  bsg_dff_en_bypass_width_p37
  \bypass.data_reg 
  (
    .clk_i(clk_i),
    .en_i(v_r),
    .data_i(data_i),
    .data_o(data_o)
  );


endmodule



module bp_pma_00
(
  clk_i,
  reset_i,
  ptag_i,
  uncached_mode_i,
  nonspec_mode_i,
  uncached_o,
  nonidem_o,
  dram_o
);

  input [27:0] ptag_i;
  input clk_i;
  input reset_i;
  input uncached_mode_i;
  input nonspec_mode_i;
  output uncached_o;
  output nonidem_o;
  output dram_o;
  wire uncached_o,nonidem_o,dram_o,is_local_addr,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,
  N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;
  assign N0 = ptag_i[26] | ptag_i[27];
  assign N1 = ptag_i[25] | N0;
  assign N2 = ptag_i[24] | N1;
  assign N3 = ptag_i[23] | N2;
  assign N4 = ptag_i[22] | N3;
  assign N5 = ptag_i[21] | N4;
  assign N6 = ptag_i[20] | N5;
  assign is_local_addr = ~N14;
  assign N14 = N13 | ptag_i[19];
  assign N13 = N12 | ptag_i[20];
  assign N12 = N11 | ptag_i[21];
  assign N11 = N10 | ptag_i[22];
  assign N10 = N9 | ptag_i[23];
  assign N9 = N8 | ptag_i[24];
  assign N8 = N7 | ptag_i[25];
  assign N7 = ptag_i[27] | ptag_i[26];
  assign uncached_o = N16 | uncached_mode_i;
  assign N16 = N15 | is_local_addr;
  assign N15 = N6 | N5;
  assign nonidem_o = N19 | nonspec_mode_i;
  assign N19 = N18 | uncached_mode_i;
  assign N18 = N17 | is_local_addr;
  assign N17 = N6 | N5;
  assign dram_o = N22 & N23;
  assign N22 = N20 & N21;
  assign N20 = ~is_local_addr;
  assign N21 = ~N5;
  assign N23 = ~N6;

endmodule



module bp_mmu_00_00000008_00000002_00000001_1
(
  clk_i,
  reset_i,
  flush_i,
  fence_i,
  priv_mode_i,
  trans_en_i,
  sum_i,
  mxr_i,
  uncached_mode_i,
  nonspec_mode_i,
  hio_mask_i,
  w_v_i,
  w_vtag_i,
  w_entry_i,
  r_v_i,
  r_instr_i,
  r_load_i,
  r_store_i,
  r_eaddr_i,
  r_size_i,
  r_cbo_i,
  r_ptw_i,
  r_v_o,
  r_ptag_o,
  r_instr_miss_o,
  r_load_miss_o,
  r_store_miss_o,
  r_uncached_o,
  r_nonidem_o,
  r_dram_o,
  r_instr_access_fault_o,
  r_load_access_fault_o,
  r_store_access_fault_o,
  r_instr_misaligned_o,
  r_load_misaligned_o,
  r_store_misaligned_o,
  r_instr_page_fault_o,
  r_load_page_fault_o,
  r_store_page_fault_o
);

  input [1:0] priv_mode_i;
  input [6:0] hio_mask_i;
  input [26:0] w_vtag_i;
  input [35:0] w_entry_i;
  input [63:0] r_eaddr_i;
  input [1:0] r_size_i;
  output [27:0] r_ptag_o;
  input clk_i;
  input reset_i;
  input flush_i;
  input fence_i;
  input trans_en_i;
  input sum_i;
  input mxr_i;
  input uncached_mode_i;
  input nonspec_mode_i;
  input w_v_i;
  input r_v_i;
  input r_instr_i;
  input r_load_i;
  input r_store_i;
  input r_cbo_i;
  input r_ptw_i;
  output r_v_o;
  output r_instr_miss_o;
  output r_load_miss_o;
  output r_store_miss_o;
  output r_uncached_o;
  output r_nonidem_o;
  output r_dram_o;
  output r_instr_access_fault_o;
  output r_load_access_fault_o;
  output r_store_access_fault_o;
  output r_instr_misaligned_o;
  output r_load_misaligned_o;
  output r_store_misaligned_o;
  output r_instr_page_fault_o;
  output r_load_page_fault_o;
  output r_store_page_fault_o;
  wire [27:0] r_ptag_o;
  wire r_v_o,r_instr_miss_o,r_load_miss_o,r_store_miss_o,r_uncached_o,r_nonidem_o,
  r_dram_o,r_instr_access_fault_o,r_load_access_fault_o,r_store_access_fault_o,
  r_instr_misaligned_o,r_load_misaligned_o,r_store_misaligned_o,r_instr_page_fault_o,
  r_load_page_fault_o,r_store_page_fault_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,
  N13,N14,N15,N16,N17,N18,N19,N20,r_misaligned,N21,N22,N23,trans_li,trans_r,
  r_misaligned_r,r_instr_r,r_load_r,r_store_r,r_cbo_r,r_ptw_r,r_v_r,tlb_r_v_li,tlb_v_li,
  N24,N25,tlb_r_v_lo,tlb_r_v_r,passthrough_entry_ptag__27_,
  passthrough_entry_ptag__26_,passthrough_entry_ptag__25_,passthrough_entry_ptag__24_,
  passthrough_entry_ptag__23_,passthrough_entry_ptag__22_,passthrough_entry_ptag__21_,
  passthrough_entry_ptag__20_,passthrough_entry_ptag__19_,passthrough_entry_ptag__18_,
  passthrough_entry_ptag__17_,passthrough_entry_ptag__16_,passthrough_entry_ptag__15_,
  passthrough_entry_ptag__14_,passthrough_entry_ptag__13_,passthrough_entry_ptag__12_,
  passthrough_entry_ptag__11_,passthrough_entry_ptag__10_,passthrough_entry_ptag__9_,
  passthrough_entry_ptag__8_,passthrough_entry_ptag__7_,passthrough_entry_ptag__6_,
  passthrough_entry_ptag__5_,passthrough_entry_ptag__4_,passthrough_entry_ptag__3_,
  passthrough_entry_ptag__2_,passthrough_entry_ptag__1_,
  passthrough_entry_ptag__0_,tlb_entry_lo_d_,tlb_entry_lo_u_,tlb_entry_lo_x_,tlb_entry_lo_w_,
  tlb_entry_lo_r_,N26,tlb_v_lo,eaddr_fault_v,cached_fault_v,hio_fault_v,instr_access_fault_v,
  load_access_fault_v,store_access_fault_v,any_access_fault_v,instr_exe_page_fault_v,
  instr_priv_page_fault_v,data_priv_page_fault,data_read_page_fault,
  data_write_page_fault,instr_page_fault_v,load_page_fault_v,store_page_fault_v,any_page_fault_v,
  any_fault_v,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,
  N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,
  N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,
  N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,
  N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,
  N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134;
  wire [51:28] r_etag_r;
  wire [26:0] tlb_vtag_li;
  wire [35:0] tlb_r_entry_lo,tlb_r_entry_r;
  assign N11 = N9 & N10;
  assign N14 = r_size_i[1] | N13;
  assign N17 = N16 | r_size_i[0];
  assign N19 = r_size_i[1] & r_size_i[0];
  assign N20 = N16 & N13;

  bsg_dff_reset_en_width_p59
  read_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(r_v_i),
    .data_i({ trans_li, r_misaligned, r_instr_i, r_load_i, r_store_i, r_cbo_i, r_ptw_i, r_eaddr_i[63:12] }),
    .data_o({ trans_r, r_misaligned_r, r_instr_r, r_load_r, r_store_r, r_cbo_r, r_ptw_r, r_etag_r, passthrough_entry_ptag__27_, passthrough_entry_ptag__26_, passthrough_entry_ptag__25_, passthrough_entry_ptag__24_, passthrough_entry_ptag__23_, passthrough_entry_ptag__22_, passthrough_entry_ptag__21_, passthrough_entry_ptag__20_, passthrough_entry_ptag__19_, passthrough_entry_ptag__18_, passthrough_entry_ptag__17_, passthrough_entry_ptag__16_, passthrough_entry_ptag__15_, passthrough_entry_ptag__14_, passthrough_entry_ptag__13_, passthrough_entry_ptag__12_, passthrough_entry_ptag__11_, passthrough_entry_ptag__10_, passthrough_entry_ptag__9_, passthrough_entry_ptag__8_, passthrough_entry_ptag__7_, passthrough_entry_ptag__6_, passthrough_entry_ptag__5_, passthrough_entry_ptag__4_, passthrough_entry_ptag__3_, passthrough_entry_ptag__2_, passthrough_entry_ptag__1_, passthrough_entry_ptag__0_ })
  );


  bsg_dff_reset_set_clear_width_p1
  r_v_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .set_i(r_v_i),
    .clear_i(flush_i),
    .data_o(r_v_r)
  );


  bp_tlb_00_00000001_00000002_00000008
  tlb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .fence_i(fence_i),
    .v_i(tlb_v_li),
    .w_i(w_v_i),
    .vtag_i(tlb_vtag_li),
    .entry_i(w_entry_i),
    .v_o(tlb_r_v_lo),
    .entry_o(tlb_r_entry_lo)
  );


  bsg_dff_sync_read_width_p37_bypass_p1
  entry_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_n_i(tlb_r_v_li),
    .data_i({ tlb_r_v_lo, tlb_r_entry_lo }),
    .data_o({ tlb_r_v_r, tlb_r_entry_r })
  );


  bp_pma_00
  pma
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ptag_i(r_ptag_o),
    .uncached_mode_i(uncached_mode_i),
    .nonspec_mode_i(nonspec_mode_i),
    .uncached_o(r_uncached_o),
    .nonidem_o(r_nonidem_o),
    .dram_o(r_dram_o)
  );

  assign N27 = r_ptag_o[26] | r_ptag_o[27];
  assign N28 = r_ptag_o[25] | N27;
  assign N29 = r_ptag_o[24] | N28;
  assign N30 = r_ptag_o[23] | N29;
  assign N31 = r_ptag_o[22] | N30;
  assign N32 = r_ptag_o[21] | N31;
  assign N33 = ~priv_mode_i[0];
  assign N34 = N33 | priv_mode_i[1];
  assign N35 = ~N34;
  assign N36 = priv_mode_i[0] | priv_mode_i[1];
  assign N37 = ~N36;
  assign N23 = (N0)? r_eaddr_i[0] : 
               (N1)? N21 : 
               (N2)? N22 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = N15;
  assign N1 = N18;
  assign N2 = N19;
  assign N3 = N20;
  assign r_misaligned = (N4)? N23 : 
                        (N12)? 1'b0 : 1'b0;
  assign N4 = N11;
  assign tlb_vtag_li = (N5)? w_vtag_i : 
                       (N6)? r_eaddr_i[38:12] : 1'b0;
  assign N5 = N25;
  assign N6 = N24;
  assign { r_ptag_o, tlb_entry_lo_d_, tlb_entry_lo_u_, tlb_entry_lo_x_, tlb_entry_lo_w_, tlb_entry_lo_r_ } = (N7)? { tlb_r_entry_r[35:8], tlb_r_entry_r[4:0] } : 
                                                                                                             (N8)? { passthrough_entry_ptag__27_, passthrough_entry_ptag__26_, passthrough_entry_ptag__25_, passthrough_entry_ptag__24_, passthrough_entry_ptag__23_, passthrough_entry_ptag__22_, passthrough_entry_ptag__21_, passthrough_entry_ptag__20_, passthrough_entry_ptag__19_, passthrough_entry_ptag__18_, passthrough_entry_ptag__17_, passthrough_entry_ptag__16_, passthrough_entry_ptag__15_, passthrough_entry_ptag__14_, passthrough_entry_ptag__13_, passthrough_entry_ptag__12_, passthrough_entry_ptag__11_, passthrough_entry_ptag__10_, passthrough_entry_ptag__9_, passthrough_entry_ptag__8_, passthrough_entry_ptag__7_, passthrough_entry_ptag__6_, passthrough_entry_ptag__5_, passthrough_entry_ptag__4_, passthrough_entry_ptag__3_, passthrough_entry_ptag__2_, passthrough_entry_ptag__1_, passthrough_entry_ptag__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N7 = trans_r;
  assign N8 = N26;
  assign tlb_v_lo = (N7)? tlb_r_v_r : 
                    (N8)? r_v_r : 1'b0;
  assign N9 = ~r_ptw_i;
  assign N10 = ~r_cbo_i;
  assign N12 = ~N11;
  assign N13 = ~r_size_i[0];
  assign N15 = ~N14;
  assign N16 = ~r_size_i[1];
  assign N18 = ~N17;
  assign N21 = r_eaddr_i[1] | r_eaddr_i[0];
  assign N22 = N38 | r_eaddr_i[0];
  assign N38 = r_eaddr_i[2] | r_eaddr_i[1];
  assign trans_li = trans_en_i & N39;
  assign N39 = ~r_ptw_i;
  assign tlb_r_v_li = r_v_i | flush_i;
  assign tlb_v_li = tlb_r_v_li | w_v_i;
  assign N24 = ~w_v_i;
  assign N25 = w_v_i;
  assign N26 = ~trans_r;
  assign eaddr_fault_v = N65 & N90;
  assign N65 = ~N64;
  assign N64 = N63 & passthrough_entry_ptag__26_;
  assign N63 = N62 & passthrough_entry_ptag__27_;
  assign N62 = N61 & r_etag_r[28];
  assign N61 = N60 & r_etag_r[29];
  assign N60 = N59 & r_etag_r[30];
  assign N59 = N58 & r_etag_r[31];
  assign N58 = N57 & r_etag_r[32];
  assign N57 = N56 & r_etag_r[33];
  assign N56 = N55 & r_etag_r[34];
  assign N55 = N54 & r_etag_r[35];
  assign N54 = N53 & r_etag_r[36];
  assign N53 = N52 & r_etag_r[37];
  assign N52 = N51 & r_etag_r[38];
  assign N51 = N50 & r_etag_r[39];
  assign N50 = N49 & r_etag_r[40];
  assign N49 = N48 & r_etag_r[41];
  assign N48 = N47 & r_etag_r[42];
  assign N47 = N46 & r_etag_r[43];
  assign N46 = N45 & r_etag_r[44];
  assign N45 = N44 & r_etag_r[45];
  assign N44 = N43 & r_etag_r[46];
  assign N43 = N42 & r_etag_r[47];
  assign N42 = N41 & r_etag_r[48];
  assign N41 = N40 & r_etag_r[49];
  assign N40 = r_etag_r[51] & r_etag_r[50];
  assign N90 = N89 | passthrough_entry_ptag__26_;
  assign N89 = N88 | passthrough_entry_ptag__27_;
  assign N88 = N87 | r_etag_r[28];
  assign N87 = N86 | r_etag_r[29];
  assign N86 = N85 | r_etag_r[30];
  assign N85 = N84 | r_etag_r[31];
  assign N84 = N83 | r_etag_r[32];
  assign N83 = N82 | r_etag_r[33];
  assign N82 = N81 | r_etag_r[34];
  assign N81 = N80 | r_etag_r[35];
  assign N80 = N79 | r_etag_r[36];
  assign N79 = N78 | r_etag_r[37];
  assign N78 = N77 | r_etag_r[38];
  assign N77 = N76 | r_etag_r[39];
  assign N76 = N75 | r_etag_r[40];
  assign N75 = N74 | r_etag_r[41];
  assign N74 = N73 | r_etag_r[42];
  assign N73 = N72 | r_etag_r[43];
  assign N72 = N71 | r_etag_r[44];
  assign N71 = N70 | r_etag_r[45];
  assign N70 = N69 | r_etag_r[46];
  assign N69 = N68 | r_etag_r[47];
  assign N68 = N67 | r_etag_r[48];
  assign N67 = N66 | r_etag_r[49];
  assign N66 = r_etag_r[51] | r_etag_r[50];
  assign cached_fault_v = N91 & r_uncached_o;
  assign N91 = r_cbo_r & tlb_v_lo;
  assign hio_fault_v = N93 | N96;
  assign N93 = N92 & N32;
  assign N92 = r_instr_r & tlb_v_lo;
  assign N96 = N94 & N95;
  assign N94 = tlb_v_lo & r_ptag_o[21];
  assign N95 = ~hio_mask_i[0];
  assign instr_access_fault_v = r_instr_r & hio_fault_v;
  assign load_access_fault_v = r_load_r & cached_fault_v;
  assign store_access_fault_v = r_store_r & cached_fault_v;
  assign any_access_fault_v = N97 | store_access_fault_v;
  assign N97 = instr_access_fault_v | load_access_fault_v;
  assign instr_exe_page_fault_v = tlb_v_lo & N98;
  assign N98 = ~tlb_entry_lo_x_;
  assign instr_priv_page_fault_v = tlb_v_lo & N102;
  assign N102 = N99 | N101;
  assign N99 = N35 & tlb_entry_lo_u_;
  assign N101 = N37 & N100;
  assign N100 = ~tlb_entry_lo_u_;
  assign data_priv_page_fault = tlb_v_lo & N107;
  assign N107 = N105 | N106;
  assign N105 = N104 & tlb_entry_lo_u_;
  assign N104 = N35 & N103;
  assign N103 = ~sum_i;
  assign N106 = N37 & N100;
  assign data_read_page_fault = tlb_v_lo & N110;
  assign N110 = ~N109;
  assign N109 = tlb_entry_lo_r_ | N108;
  assign N108 = tlb_entry_lo_x_ & mxr_i;
  assign data_write_page_fault = tlb_v_lo & N112;
  assign N112 = ~N111;
  assign N111 = tlb_entry_lo_w_ & tlb_entry_lo_d_;
  assign instr_page_fault_v = N113 & N115;
  assign N113 = trans_r & r_instr_r;
  assign N115 = N114 | eaddr_fault_v;
  assign N114 = instr_priv_page_fault_v | instr_exe_page_fault_v;
  assign load_page_fault_v = N116 & N118;
  assign N116 = trans_r & r_load_r;
  assign N118 = N117 | eaddr_fault_v;
  assign N117 = data_priv_page_fault | data_read_page_fault;
  assign store_page_fault_v = N119 & N121;
  assign N119 = trans_r & r_store_r;
  assign N121 = N120 | eaddr_fault_v;
  assign N120 = data_priv_page_fault | data_write_page_fault;
  assign any_page_fault_v = N122 | store_page_fault_v;
  assign N122 = instr_page_fault_v | load_page_fault_v;
  assign any_fault_v = any_access_fault_v | any_page_fault_v;
  assign r_v_o = N123 & N124;
  assign N123 = r_v_r & tlb_v_lo;
  assign N124 = ~any_fault_v;
  assign r_instr_miss_o = N127 & r_instr_r;
  assign N127 = N126 & N124;
  assign N126 = r_v_r & N125;
  assign N125 = ~tlb_v_lo;
  assign r_load_miss_o = N129 & r_load_r;
  assign N129 = N128 & N124;
  assign N128 = r_v_r & N125;
  assign r_store_miss_o = N131 & r_store_r;
  assign N131 = N130 & N124;
  assign N130 = r_v_r & N125;
  assign r_instr_misaligned_o = N132 & r_instr_r;
  assign N132 = r_v_r & r_misaligned_r;
  assign r_load_misaligned_o = N133 & r_load_r;
  assign N133 = r_v_r & r_misaligned_r;
  assign r_store_misaligned_o = N134 & r_store_r;
  assign N134 = r_v_r & r_misaligned_r;
  assign r_instr_access_fault_o = r_v_r & instr_access_fault_v;
  assign r_load_access_fault_o = r_v_r & load_access_fault_v;
  assign r_store_access_fault_o = r_v_r & store_access_fault_v;
  assign r_instr_page_fault_o = r_v_r & instr_page_fault_v;
  assign r_load_page_fault_o = r_v_r & load_page_fault_v;
  assign r_store_page_fault_o = r_v_r & store_page_fault_v;

endmodule



module bsg_mem_1rw_sync_mask_write_bit_000000b8_00000040_1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [183:0] data_i;
  input [5:0] addr_i;
  input [183:0] w_mask_i;
  output [183:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [183:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_mem_1rw_sync_00000040_00000200_1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_i,
  data_o
);

  input [63:0] data_i;
  input [8:0] addr_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [63:0] data_o;

  bsg_mem_1rw_sync_synth
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_dff_reset_en_0000002a
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [41:0] data_i;
  output [41:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [41:0] data_o;
  wire N0,N1,N2;
  reg data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,
  data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,
  data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,
  data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,
  data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,
  data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,
  data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,
  data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,
  data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_41_sv2v_reg <= 1'b0;
      data_o_40_sv2v_reg <= 1'b0;
      data_o_39_sv2v_reg <= 1'b0;
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mux_0000021c_2
(
  data_i,
  sel_i,
  data_o
);

  input [1079:0] data_i;
  input [0:0] sel_i;
  output [539:0] data_o;
  wire [539:0] data_o;
  wire N0,N1;
  assign data_o[539] = (N1)? data_i[539] : 
                       (N0)? data_i[1079] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[538] = (N1)? data_i[538] : 
                       (N0)? data_i[1078] : 1'b0;
  assign data_o[537] = (N1)? data_i[537] : 
                       (N0)? data_i[1077] : 1'b0;
  assign data_o[536] = (N1)? data_i[536] : 
                       (N0)? data_i[1076] : 1'b0;
  assign data_o[535] = (N1)? data_i[535] : 
                       (N0)? data_i[1075] : 1'b0;
  assign data_o[534] = (N1)? data_i[534] : 
                       (N0)? data_i[1074] : 1'b0;
  assign data_o[533] = (N1)? data_i[533] : 
                       (N0)? data_i[1073] : 1'b0;
  assign data_o[532] = (N1)? data_i[532] : 
                       (N0)? data_i[1072] : 1'b0;
  assign data_o[531] = (N1)? data_i[531] : 
                       (N0)? data_i[1071] : 1'b0;
  assign data_o[530] = (N1)? data_i[530] : 
                       (N0)? data_i[1070] : 1'b0;
  assign data_o[529] = (N1)? data_i[529] : 
                       (N0)? data_i[1069] : 1'b0;
  assign data_o[528] = (N1)? data_i[528] : 
                       (N0)? data_i[1068] : 1'b0;
  assign data_o[527] = (N1)? data_i[527] : 
                       (N0)? data_i[1067] : 1'b0;
  assign data_o[526] = (N1)? data_i[526] : 
                       (N0)? data_i[1066] : 1'b0;
  assign data_o[525] = (N1)? data_i[525] : 
                       (N0)? data_i[1065] : 1'b0;
  assign data_o[524] = (N1)? data_i[524] : 
                       (N0)? data_i[1064] : 1'b0;
  assign data_o[523] = (N1)? data_i[523] : 
                       (N0)? data_i[1063] : 1'b0;
  assign data_o[522] = (N1)? data_i[522] : 
                       (N0)? data_i[1062] : 1'b0;
  assign data_o[521] = (N1)? data_i[521] : 
                       (N0)? data_i[1061] : 1'b0;
  assign data_o[520] = (N1)? data_i[520] : 
                       (N0)? data_i[1060] : 1'b0;
  assign data_o[519] = (N1)? data_i[519] : 
                       (N0)? data_i[1059] : 1'b0;
  assign data_o[518] = (N1)? data_i[518] : 
                       (N0)? data_i[1058] : 1'b0;
  assign data_o[517] = (N1)? data_i[517] : 
                       (N0)? data_i[1057] : 1'b0;
  assign data_o[516] = (N1)? data_i[516] : 
                       (N0)? data_i[1056] : 1'b0;
  assign data_o[515] = (N1)? data_i[515] : 
                       (N0)? data_i[1055] : 1'b0;
  assign data_o[514] = (N1)? data_i[514] : 
                       (N0)? data_i[1054] : 1'b0;
  assign data_o[513] = (N1)? data_i[513] : 
                       (N0)? data_i[1053] : 1'b0;
  assign data_o[512] = (N1)? data_i[512] : 
                       (N0)? data_i[1052] : 1'b0;
  assign data_o[511] = (N1)? data_i[511] : 
                       (N0)? data_i[1051] : 1'b0;
  assign data_o[510] = (N1)? data_i[510] : 
                       (N0)? data_i[1050] : 1'b0;
  assign data_o[509] = (N1)? data_i[509] : 
                       (N0)? data_i[1049] : 1'b0;
  assign data_o[508] = (N1)? data_i[508] : 
                       (N0)? data_i[1048] : 1'b0;
  assign data_o[507] = (N1)? data_i[507] : 
                       (N0)? data_i[1047] : 1'b0;
  assign data_o[506] = (N1)? data_i[506] : 
                       (N0)? data_i[1046] : 1'b0;
  assign data_o[505] = (N1)? data_i[505] : 
                       (N0)? data_i[1045] : 1'b0;
  assign data_o[504] = (N1)? data_i[504] : 
                       (N0)? data_i[1044] : 1'b0;
  assign data_o[503] = (N1)? data_i[503] : 
                       (N0)? data_i[1043] : 1'b0;
  assign data_o[502] = (N1)? data_i[502] : 
                       (N0)? data_i[1042] : 1'b0;
  assign data_o[501] = (N1)? data_i[501] : 
                       (N0)? data_i[1041] : 1'b0;
  assign data_o[500] = (N1)? data_i[500] : 
                       (N0)? data_i[1040] : 1'b0;
  assign data_o[499] = (N1)? data_i[499] : 
                       (N0)? data_i[1039] : 1'b0;
  assign data_o[498] = (N1)? data_i[498] : 
                       (N0)? data_i[1038] : 1'b0;
  assign data_o[497] = (N1)? data_i[497] : 
                       (N0)? data_i[1037] : 1'b0;
  assign data_o[496] = (N1)? data_i[496] : 
                       (N0)? data_i[1036] : 1'b0;
  assign data_o[495] = (N1)? data_i[495] : 
                       (N0)? data_i[1035] : 1'b0;
  assign data_o[494] = (N1)? data_i[494] : 
                       (N0)? data_i[1034] : 1'b0;
  assign data_o[493] = (N1)? data_i[493] : 
                       (N0)? data_i[1033] : 1'b0;
  assign data_o[492] = (N1)? data_i[492] : 
                       (N0)? data_i[1032] : 1'b0;
  assign data_o[491] = (N1)? data_i[491] : 
                       (N0)? data_i[1031] : 1'b0;
  assign data_o[490] = (N1)? data_i[490] : 
                       (N0)? data_i[1030] : 1'b0;
  assign data_o[489] = (N1)? data_i[489] : 
                       (N0)? data_i[1029] : 1'b0;
  assign data_o[488] = (N1)? data_i[488] : 
                       (N0)? data_i[1028] : 1'b0;
  assign data_o[487] = (N1)? data_i[487] : 
                       (N0)? data_i[1027] : 1'b0;
  assign data_o[486] = (N1)? data_i[486] : 
                       (N0)? data_i[1026] : 1'b0;
  assign data_o[485] = (N1)? data_i[485] : 
                       (N0)? data_i[1025] : 1'b0;
  assign data_o[484] = (N1)? data_i[484] : 
                       (N0)? data_i[1024] : 1'b0;
  assign data_o[483] = (N1)? data_i[483] : 
                       (N0)? data_i[1023] : 1'b0;
  assign data_o[482] = (N1)? data_i[482] : 
                       (N0)? data_i[1022] : 1'b0;
  assign data_o[481] = (N1)? data_i[481] : 
                       (N0)? data_i[1021] : 1'b0;
  assign data_o[480] = (N1)? data_i[480] : 
                       (N0)? data_i[1020] : 1'b0;
  assign data_o[479] = (N1)? data_i[479] : 
                       (N0)? data_i[1019] : 1'b0;
  assign data_o[478] = (N1)? data_i[478] : 
                       (N0)? data_i[1018] : 1'b0;
  assign data_o[477] = (N1)? data_i[477] : 
                       (N0)? data_i[1017] : 1'b0;
  assign data_o[476] = (N1)? data_i[476] : 
                       (N0)? data_i[1016] : 1'b0;
  assign data_o[475] = (N1)? data_i[475] : 
                       (N0)? data_i[1015] : 1'b0;
  assign data_o[474] = (N1)? data_i[474] : 
                       (N0)? data_i[1014] : 1'b0;
  assign data_o[473] = (N1)? data_i[473] : 
                       (N0)? data_i[1013] : 1'b0;
  assign data_o[472] = (N1)? data_i[472] : 
                       (N0)? data_i[1012] : 1'b0;
  assign data_o[471] = (N1)? data_i[471] : 
                       (N0)? data_i[1011] : 1'b0;
  assign data_o[470] = (N1)? data_i[470] : 
                       (N0)? data_i[1010] : 1'b0;
  assign data_o[469] = (N1)? data_i[469] : 
                       (N0)? data_i[1009] : 1'b0;
  assign data_o[468] = (N1)? data_i[468] : 
                       (N0)? data_i[1008] : 1'b0;
  assign data_o[467] = (N1)? data_i[467] : 
                       (N0)? data_i[1007] : 1'b0;
  assign data_o[466] = (N1)? data_i[466] : 
                       (N0)? data_i[1006] : 1'b0;
  assign data_o[465] = (N1)? data_i[465] : 
                       (N0)? data_i[1005] : 1'b0;
  assign data_o[464] = (N1)? data_i[464] : 
                       (N0)? data_i[1004] : 1'b0;
  assign data_o[463] = (N1)? data_i[463] : 
                       (N0)? data_i[1003] : 1'b0;
  assign data_o[462] = (N1)? data_i[462] : 
                       (N0)? data_i[1002] : 1'b0;
  assign data_o[461] = (N1)? data_i[461] : 
                       (N0)? data_i[1001] : 1'b0;
  assign data_o[460] = (N1)? data_i[460] : 
                       (N0)? data_i[1000] : 1'b0;
  assign data_o[459] = (N1)? data_i[459] : 
                       (N0)? data_i[999] : 1'b0;
  assign data_o[458] = (N1)? data_i[458] : 
                       (N0)? data_i[998] : 1'b0;
  assign data_o[457] = (N1)? data_i[457] : 
                       (N0)? data_i[997] : 1'b0;
  assign data_o[456] = (N1)? data_i[456] : 
                       (N0)? data_i[996] : 1'b0;
  assign data_o[455] = (N1)? data_i[455] : 
                       (N0)? data_i[995] : 1'b0;
  assign data_o[454] = (N1)? data_i[454] : 
                       (N0)? data_i[994] : 1'b0;
  assign data_o[453] = (N1)? data_i[453] : 
                       (N0)? data_i[993] : 1'b0;
  assign data_o[452] = (N1)? data_i[452] : 
                       (N0)? data_i[992] : 1'b0;
  assign data_o[451] = (N1)? data_i[451] : 
                       (N0)? data_i[991] : 1'b0;
  assign data_o[450] = (N1)? data_i[450] : 
                       (N0)? data_i[990] : 1'b0;
  assign data_o[449] = (N1)? data_i[449] : 
                       (N0)? data_i[989] : 1'b0;
  assign data_o[448] = (N1)? data_i[448] : 
                       (N0)? data_i[988] : 1'b0;
  assign data_o[447] = (N1)? data_i[447] : 
                       (N0)? data_i[987] : 1'b0;
  assign data_o[446] = (N1)? data_i[446] : 
                       (N0)? data_i[986] : 1'b0;
  assign data_o[445] = (N1)? data_i[445] : 
                       (N0)? data_i[985] : 1'b0;
  assign data_o[444] = (N1)? data_i[444] : 
                       (N0)? data_i[984] : 1'b0;
  assign data_o[443] = (N1)? data_i[443] : 
                       (N0)? data_i[983] : 1'b0;
  assign data_o[442] = (N1)? data_i[442] : 
                       (N0)? data_i[982] : 1'b0;
  assign data_o[441] = (N1)? data_i[441] : 
                       (N0)? data_i[981] : 1'b0;
  assign data_o[440] = (N1)? data_i[440] : 
                       (N0)? data_i[980] : 1'b0;
  assign data_o[439] = (N1)? data_i[439] : 
                       (N0)? data_i[979] : 1'b0;
  assign data_o[438] = (N1)? data_i[438] : 
                       (N0)? data_i[978] : 1'b0;
  assign data_o[437] = (N1)? data_i[437] : 
                       (N0)? data_i[977] : 1'b0;
  assign data_o[436] = (N1)? data_i[436] : 
                       (N0)? data_i[976] : 1'b0;
  assign data_o[435] = (N1)? data_i[435] : 
                       (N0)? data_i[975] : 1'b0;
  assign data_o[434] = (N1)? data_i[434] : 
                       (N0)? data_i[974] : 1'b0;
  assign data_o[433] = (N1)? data_i[433] : 
                       (N0)? data_i[973] : 1'b0;
  assign data_o[432] = (N1)? data_i[432] : 
                       (N0)? data_i[972] : 1'b0;
  assign data_o[431] = (N1)? data_i[431] : 
                       (N0)? data_i[971] : 1'b0;
  assign data_o[430] = (N1)? data_i[430] : 
                       (N0)? data_i[970] : 1'b0;
  assign data_o[429] = (N1)? data_i[429] : 
                       (N0)? data_i[969] : 1'b0;
  assign data_o[428] = (N1)? data_i[428] : 
                       (N0)? data_i[968] : 1'b0;
  assign data_o[427] = (N1)? data_i[427] : 
                       (N0)? data_i[967] : 1'b0;
  assign data_o[426] = (N1)? data_i[426] : 
                       (N0)? data_i[966] : 1'b0;
  assign data_o[425] = (N1)? data_i[425] : 
                       (N0)? data_i[965] : 1'b0;
  assign data_o[424] = (N1)? data_i[424] : 
                       (N0)? data_i[964] : 1'b0;
  assign data_o[423] = (N1)? data_i[423] : 
                       (N0)? data_i[963] : 1'b0;
  assign data_o[422] = (N1)? data_i[422] : 
                       (N0)? data_i[962] : 1'b0;
  assign data_o[421] = (N1)? data_i[421] : 
                       (N0)? data_i[961] : 1'b0;
  assign data_o[420] = (N1)? data_i[420] : 
                       (N0)? data_i[960] : 1'b0;
  assign data_o[419] = (N1)? data_i[419] : 
                       (N0)? data_i[959] : 1'b0;
  assign data_o[418] = (N1)? data_i[418] : 
                       (N0)? data_i[958] : 1'b0;
  assign data_o[417] = (N1)? data_i[417] : 
                       (N0)? data_i[957] : 1'b0;
  assign data_o[416] = (N1)? data_i[416] : 
                       (N0)? data_i[956] : 1'b0;
  assign data_o[415] = (N1)? data_i[415] : 
                       (N0)? data_i[955] : 1'b0;
  assign data_o[414] = (N1)? data_i[414] : 
                       (N0)? data_i[954] : 1'b0;
  assign data_o[413] = (N1)? data_i[413] : 
                       (N0)? data_i[953] : 1'b0;
  assign data_o[412] = (N1)? data_i[412] : 
                       (N0)? data_i[952] : 1'b0;
  assign data_o[411] = (N1)? data_i[411] : 
                       (N0)? data_i[951] : 1'b0;
  assign data_o[410] = (N1)? data_i[410] : 
                       (N0)? data_i[950] : 1'b0;
  assign data_o[409] = (N1)? data_i[409] : 
                       (N0)? data_i[949] : 1'b0;
  assign data_o[408] = (N1)? data_i[408] : 
                       (N0)? data_i[948] : 1'b0;
  assign data_o[407] = (N1)? data_i[407] : 
                       (N0)? data_i[947] : 1'b0;
  assign data_o[406] = (N1)? data_i[406] : 
                       (N0)? data_i[946] : 1'b0;
  assign data_o[405] = (N1)? data_i[405] : 
                       (N0)? data_i[945] : 1'b0;
  assign data_o[404] = (N1)? data_i[404] : 
                       (N0)? data_i[944] : 1'b0;
  assign data_o[403] = (N1)? data_i[403] : 
                       (N0)? data_i[943] : 1'b0;
  assign data_o[402] = (N1)? data_i[402] : 
                       (N0)? data_i[942] : 1'b0;
  assign data_o[401] = (N1)? data_i[401] : 
                       (N0)? data_i[941] : 1'b0;
  assign data_o[400] = (N1)? data_i[400] : 
                       (N0)? data_i[940] : 1'b0;
  assign data_o[399] = (N1)? data_i[399] : 
                       (N0)? data_i[939] : 1'b0;
  assign data_o[398] = (N1)? data_i[398] : 
                       (N0)? data_i[938] : 1'b0;
  assign data_o[397] = (N1)? data_i[397] : 
                       (N0)? data_i[937] : 1'b0;
  assign data_o[396] = (N1)? data_i[396] : 
                       (N0)? data_i[936] : 1'b0;
  assign data_o[395] = (N1)? data_i[395] : 
                       (N0)? data_i[935] : 1'b0;
  assign data_o[394] = (N1)? data_i[394] : 
                       (N0)? data_i[934] : 1'b0;
  assign data_o[393] = (N1)? data_i[393] : 
                       (N0)? data_i[933] : 1'b0;
  assign data_o[392] = (N1)? data_i[392] : 
                       (N0)? data_i[932] : 1'b0;
  assign data_o[391] = (N1)? data_i[391] : 
                       (N0)? data_i[931] : 1'b0;
  assign data_o[390] = (N1)? data_i[390] : 
                       (N0)? data_i[930] : 1'b0;
  assign data_o[389] = (N1)? data_i[389] : 
                       (N0)? data_i[929] : 1'b0;
  assign data_o[388] = (N1)? data_i[388] : 
                       (N0)? data_i[928] : 1'b0;
  assign data_o[387] = (N1)? data_i[387] : 
                       (N0)? data_i[927] : 1'b0;
  assign data_o[386] = (N1)? data_i[386] : 
                       (N0)? data_i[926] : 1'b0;
  assign data_o[385] = (N1)? data_i[385] : 
                       (N0)? data_i[925] : 1'b0;
  assign data_o[384] = (N1)? data_i[384] : 
                       (N0)? data_i[924] : 1'b0;
  assign data_o[383] = (N1)? data_i[383] : 
                       (N0)? data_i[923] : 1'b0;
  assign data_o[382] = (N1)? data_i[382] : 
                       (N0)? data_i[922] : 1'b0;
  assign data_o[381] = (N1)? data_i[381] : 
                       (N0)? data_i[921] : 1'b0;
  assign data_o[380] = (N1)? data_i[380] : 
                       (N0)? data_i[920] : 1'b0;
  assign data_o[379] = (N1)? data_i[379] : 
                       (N0)? data_i[919] : 1'b0;
  assign data_o[378] = (N1)? data_i[378] : 
                       (N0)? data_i[918] : 1'b0;
  assign data_o[377] = (N1)? data_i[377] : 
                       (N0)? data_i[917] : 1'b0;
  assign data_o[376] = (N1)? data_i[376] : 
                       (N0)? data_i[916] : 1'b0;
  assign data_o[375] = (N1)? data_i[375] : 
                       (N0)? data_i[915] : 1'b0;
  assign data_o[374] = (N1)? data_i[374] : 
                       (N0)? data_i[914] : 1'b0;
  assign data_o[373] = (N1)? data_i[373] : 
                       (N0)? data_i[913] : 1'b0;
  assign data_o[372] = (N1)? data_i[372] : 
                       (N0)? data_i[912] : 1'b0;
  assign data_o[371] = (N1)? data_i[371] : 
                       (N0)? data_i[911] : 1'b0;
  assign data_o[370] = (N1)? data_i[370] : 
                       (N0)? data_i[910] : 1'b0;
  assign data_o[369] = (N1)? data_i[369] : 
                       (N0)? data_i[909] : 1'b0;
  assign data_o[368] = (N1)? data_i[368] : 
                       (N0)? data_i[908] : 1'b0;
  assign data_o[367] = (N1)? data_i[367] : 
                       (N0)? data_i[907] : 1'b0;
  assign data_o[366] = (N1)? data_i[366] : 
                       (N0)? data_i[906] : 1'b0;
  assign data_o[365] = (N1)? data_i[365] : 
                       (N0)? data_i[905] : 1'b0;
  assign data_o[364] = (N1)? data_i[364] : 
                       (N0)? data_i[904] : 1'b0;
  assign data_o[363] = (N1)? data_i[363] : 
                       (N0)? data_i[903] : 1'b0;
  assign data_o[362] = (N1)? data_i[362] : 
                       (N0)? data_i[902] : 1'b0;
  assign data_o[361] = (N1)? data_i[361] : 
                       (N0)? data_i[901] : 1'b0;
  assign data_o[360] = (N1)? data_i[360] : 
                       (N0)? data_i[900] : 1'b0;
  assign data_o[359] = (N1)? data_i[359] : 
                       (N0)? data_i[899] : 1'b0;
  assign data_o[358] = (N1)? data_i[358] : 
                       (N0)? data_i[898] : 1'b0;
  assign data_o[357] = (N1)? data_i[357] : 
                       (N0)? data_i[897] : 1'b0;
  assign data_o[356] = (N1)? data_i[356] : 
                       (N0)? data_i[896] : 1'b0;
  assign data_o[355] = (N1)? data_i[355] : 
                       (N0)? data_i[895] : 1'b0;
  assign data_o[354] = (N1)? data_i[354] : 
                       (N0)? data_i[894] : 1'b0;
  assign data_o[353] = (N1)? data_i[353] : 
                       (N0)? data_i[893] : 1'b0;
  assign data_o[352] = (N1)? data_i[352] : 
                       (N0)? data_i[892] : 1'b0;
  assign data_o[351] = (N1)? data_i[351] : 
                       (N0)? data_i[891] : 1'b0;
  assign data_o[350] = (N1)? data_i[350] : 
                       (N0)? data_i[890] : 1'b0;
  assign data_o[349] = (N1)? data_i[349] : 
                       (N0)? data_i[889] : 1'b0;
  assign data_o[348] = (N1)? data_i[348] : 
                       (N0)? data_i[888] : 1'b0;
  assign data_o[347] = (N1)? data_i[347] : 
                       (N0)? data_i[887] : 1'b0;
  assign data_o[346] = (N1)? data_i[346] : 
                       (N0)? data_i[886] : 1'b0;
  assign data_o[345] = (N1)? data_i[345] : 
                       (N0)? data_i[885] : 1'b0;
  assign data_o[344] = (N1)? data_i[344] : 
                       (N0)? data_i[884] : 1'b0;
  assign data_o[343] = (N1)? data_i[343] : 
                       (N0)? data_i[883] : 1'b0;
  assign data_o[342] = (N1)? data_i[342] : 
                       (N0)? data_i[882] : 1'b0;
  assign data_o[341] = (N1)? data_i[341] : 
                       (N0)? data_i[881] : 1'b0;
  assign data_o[340] = (N1)? data_i[340] : 
                       (N0)? data_i[880] : 1'b0;
  assign data_o[339] = (N1)? data_i[339] : 
                       (N0)? data_i[879] : 1'b0;
  assign data_o[338] = (N1)? data_i[338] : 
                       (N0)? data_i[878] : 1'b0;
  assign data_o[337] = (N1)? data_i[337] : 
                       (N0)? data_i[877] : 1'b0;
  assign data_o[336] = (N1)? data_i[336] : 
                       (N0)? data_i[876] : 1'b0;
  assign data_o[335] = (N1)? data_i[335] : 
                       (N0)? data_i[875] : 1'b0;
  assign data_o[334] = (N1)? data_i[334] : 
                       (N0)? data_i[874] : 1'b0;
  assign data_o[333] = (N1)? data_i[333] : 
                       (N0)? data_i[873] : 1'b0;
  assign data_o[332] = (N1)? data_i[332] : 
                       (N0)? data_i[872] : 1'b0;
  assign data_o[331] = (N1)? data_i[331] : 
                       (N0)? data_i[871] : 1'b0;
  assign data_o[330] = (N1)? data_i[330] : 
                       (N0)? data_i[870] : 1'b0;
  assign data_o[329] = (N1)? data_i[329] : 
                       (N0)? data_i[869] : 1'b0;
  assign data_o[328] = (N1)? data_i[328] : 
                       (N0)? data_i[868] : 1'b0;
  assign data_o[327] = (N1)? data_i[327] : 
                       (N0)? data_i[867] : 1'b0;
  assign data_o[326] = (N1)? data_i[326] : 
                       (N0)? data_i[866] : 1'b0;
  assign data_o[325] = (N1)? data_i[325] : 
                       (N0)? data_i[865] : 1'b0;
  assign data_o[324] = (N1)? data_i[324] : 
                       (N0)? data_i[864] : 1'b0;
  assign data_o[323] = (N1)? data_i[323] : 
                       (N0)? data_i[863] : 1'b0;
  assign data_o[322] = (N1)? data_i[322] : 
                       (N0)? data_i[862] : 1'b0;
  assign data_o[321] = (N1)? data_i[321] : 
                       (N0)? data_i[861] : 1'b0;
  assign data_o[320] = (N1)? data_i[320] : 
                       (N0)? data_i[860] : 1'b0;
  assign data_o[319] = (N1)? data_i[319] : 
                       (N0)? data_i[859] : 1'b0;
  assign data_o[318] = (N1)? data_i[318] : 
                       (N0)? data_i[858] : 1'b0;
  assign data_o[317] = (N1)? data_i[317] : 
                       (N0)? data_i[857] : 1'b0;
  assign data_o[316] = (N1)? data_i[316] : 
                       (N0)? data_i[856] : 1'b0;
  assign data_o[315] = (N1)? data_i[315] : 
                       (N0)? data_i[855] : 1'b0;
  assign data_o[314] = (N1)? data_i[314] : 
                       (N0)? data_i[854] : 1'b0;
  assign data_o[313] = (N1)? data_i[313] : 
                       (N0)? data_i[853] : 1'b0;
  assign data_o[312] = (N1)? data_i[312] : 
                       (N0)? data_i[852] : 1'b0;
  assign data_o[311] = (N1)? data_i[311] : 
                       (N0)? data_i[851] : 1'b0;
  assign data_o[310] = (N1)? data_i[310] : 
                       (N0)? data_i[850] : 1'b0;
  assign data_o[309] = (N1)? data_i[309] : 
                       (N0)? data_i[849] : 1'b0;
  assign data_o[308] = (N1)? data_i[308] : 
                       (N0)? data_i[848] : 1'b0;
  assign data_o[307] = (N1)? data_i[307] : 
                       (N0)? data_i[847] : 1'b0;
  assign data_o[306] = (N1)? data_i[306] : 
                       (N0)? data_i[846] : 1'b0;
  assign data_o[305] = (N1)? data_i[305] : 
                       (N0)? data_i[845] : 1'b0;
  assign data_o[304] = (N1)? data_i[304] : 
                       (N0)? data_i[844] : 1'b0;
  assign data_o[303] = (N1)? data_i[303] : 
                       (N0)? data_i[843] : 1'b0;
  assign data_o[302] = (N1)? data_i[302] : 
                       (N0)? data_i[842] : 1'b0;
  assign data_o[301] = (N1)? data_i[301] : 
                       (N0)? data_i[841] : 1'b0;
  assign data_o[300] = (N1)? data_i[300] : 
                       (N0)? data_i[840] : 1'b0;
  assign data_o[299] = (N1)? data_i[299] : 
                       (N0)? data_i[839] : 1'b0;
  assign data_o[298] = (N1)? data_i[298] : 
                       (N0)? data_i[838] : 1'b0;
  assign data_o[297] = (N1)? data_i[297] : 
                       (N0)? data_i[837] : 1'b0;
  assign data_o[296] = (N1)? data_i[296] : 
                       (N0)? data_i[836] : 1'b0;
  assign data_o[295] = (N1)? data_i[295] : 
                       (N0)? data_i[835] : 1'b0;
  assign data_o[294] = (N1)? data_i[294] : 
                       (N0)? data_i[834] : 1'b0;
  assign data_o[293] = (N1)? data_i[293] : 
                       (N0)? data_i[833] : 1'b0;
  assign data_o[292] = (N1)? data_i[292] : 
                       (N0)? data_i[832] : 1'b0;
  assign data_o[291] = (N1)? data_i[291] : 
                       (N0)? data_i[831] : 1'b0;
  assign data_o[290] = (N1)? data_i[290] : 
                       (N0)? data_i[830] : 1'b0;
  assign data_o[289] = (N1)? data_i[289] : 
                       (N0)? data_i[829] : 1'b0;
  assign data_o[288] = (N1)? data_i[288] : 
                       (N0)? data_i[828] : 1'b0;
  assign data_o[287] = (N1)? data_i[287] : 
                       (N0)? data_i[827] : 1'b0;
  assign data_o[286] = (N1)? data_i[286] : 
                       (N0)? data_i[826] : 1'b0;
  assign data_o[285] = (N1)? data_i[285] : 
                       (N0)? data_i[825] : 1'b0;
  assign data_o[284] = (N1)? data_i[284] : 
                       (N0)? data_i[824] : 1'b0;
  assign data_o[283] = (N1)? data_i[283] : 
                       (N0)? data_i[823] : 1'b0;
  assign data_o[282] = (N1)? data_i[282] : 
                       (N0)? data_i[822] : 1'b0;
  assign data_o[281] = (N1)? data_i[281] : 
                       (N0)? data_i[821] : 1'b0;
  assign data_o[280] = (N1)? data_i[280] : 
                       (N0)? data_i[820] : 1'b0;
  assign data_o[279] = (N1)? data_i[279] : 
                       (N0)? data_i[819] : 1'b0;
  assign data_o[278] = (N1)? data_i[278] : 
                       (N0)? data_i[818] : 1'b0;
  assign data_o[277] = (N1)? data_i[277] : 
                       (N0)? data_i[817] : 1'b0;
  assign data_o[276] = (N1)? data_i[276] : 
                       (N0)? data_i[816] : 1'b0;
  assign data_o[275] = (N1)? data_i[275] : 
                       (N0)? data_i[815] : 1'b0;
  assign data_o[274] = (N1)? data_i[274] : 
                       (N0)? data_i[814] : 1'b0;
  assign data_o[273] = (N1)? data_i[273] : 
                       (N0)? data_i[813] : 1'b0;
  assign data_o[272] = (N1)? data_i[272] : 
                       (N0)? data_i[812] : 1'b0;
  assign data_o[271] = (N1)? data_i[271] : 
                       (N0)? data_i[811] : 1'b0;
  assign data_o[270] = (N1)? data_i[270] : 
                       (N0)? data_i[810] : 1'b0;
  assign data_o[269] = (N1)? data_i[269] : 
                       (N0)? data_i[809] : 1'b0;
  assign data_o[268] = (N1)? data_i[268] : 
                       (N0)? data_i[808] : 1'b0;
  assign data_o[267] = (N1)? data_i[267] : 
                       (N0)? data_i[807] : 1'b0;
  assign data_o[266] = (N1)? data_i[266] : 
                       (N0)? data_i[806] : 1'b0;
  assign data_o[265] = (N1)? data_i[265] : 
                       (N0)? data_i[805] : 1'b0;
  assign data_o[264] = (N1)? data_i[264] : 
                       (N0)? data_i[804] : 1'b0;
  assign data_o[263] = (N1)? data_i[263] : 
                       (N0)? data_i[803] : 1'b0;
  assign data_o[262] = (N1)? data_i[262] : 
                       (N0)? data_i[802] : 1'b0;
  assign data_o[261] = (N1)? data_i[261] : 
                       (N0)? data_i[801] : 1'b0;
  assign data_o[260] = (N1)? data_i[260] : 
                       (N0)? data_i[800] : 1'b0;
  assign data_o[259] = (N1)? data_i[259] : 
                       (N0)? data_i[799] : 1'b0;
  assign data_o[258] = (N1)? data_i[258] : 
                       (N0)? data_i[798] : 1'b0;
  assign data_o[257] = (N1)? data_i[257] : 
                       (N0)? data_i[797] : 1'b0;
  assign data_o[256] = (N1)? data_i[256] : 
                       (N0)? data_i[796] : 1'b0;
  assign data_o[255] = (N1)? data_i[255] : 
                       (N0)? data_i[795] : 1'b0;
  assign data_o[254] = (N1)? data_i[254] : 
                       (N0)? data_i[794] : 1'b0;
  assign data_o[253] = (N1)? data_i[253] : 
                       (N0)? data_i[793] : 1'b0;
  assign data_o[252] = (N1)? data_i[252] : 
                       (N0)? data_i[792] : 1'b0;
  assign data_o[251] = (N1)? data_i[251] : 
                       (N0)? data_i[791] : 1'b0;
  assign data_o[250] = (N1)? data_i[250] : 
                       (N0)? data_i[790] : 1'b0;
  assign data_o[249] = (N1)? data_i[249] : 
                       (N0)? data_i[789] : 1'b0;
  assign data_o[248] = (N1)? data_i[248] : 
                       (N0)? data_i[788] : 1'b0;
  assign data_o[247] = (N1)? data_i[247] : 
                       (N0)? data_i[787] : 1'b0;
  assign data_o[246] = (N1)? data_i[246] : 
                       (N0)? data_i[786] : 1'b0;
  assign data_o[245] = (N1)? data_i[245] : 
                       (N0)? data_i[785] : 1'b0;
  assign data_o[244] = (N1)? data_i[244] : 
                       (N0)? data_i[784] : 1'b0;
  assign data_o[243] = (N1)? data_i[243] : 
                       (N0)? data_i[783] : 1'b0;
  assign data_o[242] = (N1)? data_i[242] : 
                       (N0)? data_i[782] : 1'b0;
  assign data_o[241] = (N1)? data_i[241] : 
                       (N0)? data_i[781] : 1'b0;
  assign data_o[240] = (N1)? data_i[240] : 
                       (N0)? data_i[780] : 1'b0;
  assign data_o[239] = (N1)? data_i[239] : 
                       (N0)? data_i[779] : 1'b0;
  assign data_o[238] = (N1)? data_i[238] : 
                       (N0)? data_i[778] : 1'b0;
  assign data_o[237] = (N1)? data_i[237] : 
                       (N0)? data_i[777] : 1'b0;
  assign data_o[236] = (N1)? data_i[236] : 
                       (N0)? data_i[776] : 1'b0;
  assign data_o[235] = (N1)? data_i[235] : 
                       (N0)? data_i[775] : 1'b0;
  assign data_o[234] = (N1)? data_i[234] : 
                       (N0)? data_i[774] : 1'b0;
  assign data_o[233] = (N1)? data_i[233] : 
                       (N0)? data_i[773] : 1'b0;
  assign data_o[232] = (N1)? data_i[232] : 
                       (N0)? data_i[772] : 1'b0;
  assign data_o[231] = (N1)? data_i[231] : 
                       (N0)? data_i[771] : 1'b0;
  assign data_o[230] = (N1)? data_i[230] : 
                       (N0)? data_i[770] : 1'b0;
  assign data_o[229] = (N1)? data_i[229] : 
                       (N0)? data_i[769] : 1'b0;
  assign data_o[228] = (N1)? data_i[228] : 
                       (N0)? data_i[768] : 1'b0;
  assign data_o[227] = (N1)? data_i[227] : 
                       (N0)? data_i[767] : 1'b0;
  assign data_o[226] = (N1)? data_i[226] : 
                       (N0)? data_i[766] : 1'b0;
  assign data_o[225] = (N1)? data_i[225] : 
                       (N0)? data_i[765] : 1'b0;
  assign data_o[224] = (N1)? data_i[224] : 
                       (N0)? data_i[764] : 1'b0;
  assign data_o[223] = (N1)? data_i[223] : 
                       (N0)? data_i[763] : 1'b0;
  assign data_o[222] = (N1)? data_i[222] : 
                       (N0)? data_i[762] : 1'b0;
  assign data_o[221] = (N1)? data_i[221] : 
                       (N0)? data_i[761] : 1'b0;
  assign data_o[220] = (N1)? data_i[220] : 
                       (N0)? data_i[760] : 1'b0;
  assign data_o[219] = (N1)? data_i[219] : 
                       (N0)? data_i[759] : 1'b0;
  assign data_o[218] = (N1)? data_i[218] : 
                       (N0)? data_i[758] : 1'b0;
  assign data_o[217] = (N1)? data_i[217] : 
                       (N0)? data_i[757] : 1'b0;
  assign data_o[216] = (N1)? data_i[216] : 
                       (N0)? data_i[756] : 1'b0;
  assign data_o[215] = (N1)? data_i[215] : 
                       (N0)? data_i[755] : 1'b0;
  assign data_o[214] = (N1)? data_i[214] : 
                       (N0)? data_i[754] : 1'b0;
  assign data_o[213] = (N1)? data_i[213] : 
                       (N0)? data_i[753] : 1'b0;
  assign data_o[212] = (N1)? data_i[212] : 
                       (N0)? data_i[752] : 1'b0;
  assign data_o[211] = (N1)? data_i[211] : 
                       (N0)? data_i[751] : 1'b0;
  assign data_o[210] = (N1)? data_i[210] : 
                       (N0)? data_i[750] : 1'b0;
  assign data_o[209] = (N1)? data_i[209] : 
                       (N0)? data_i[749] : 1'b0;
  assign data_o[208] = (N1)? data_i[208] : 
                       (N0)? data_i[748] : 1'b0;
  assign data_o[207] = (N1)? data_i[207] : 
                       (N0)? data_i[747] : 1'b0;
  assign data_o[206] = (N1)? data_i[206] : 
                       (N0)? data_i[746] : 1'b0;
  assign data_o[205] = (N1)? data_i[205] : 
                       (N0)? data_i[745] : 1'b0;
  assign data_o[204] = (N1)? data_i[204] : 
                       (N0)? data_i[744] : 1'b0;
  assign data_o[203] = (N1)? data_i[203] : 
                       (N0)? data_i[743] : 1'b0;
  assign data_o[202] = (N1)? data_i[202] : 
                       (N0)? data_i[742] : 1'b0;
  assign data_o[201] = (N1)? data_i[201] : 
                       (N0)? data_i[741] : 1'b0;
  assign data_o[200] = (N1)? data_i[200] : 
                       (N0)? data_i[740] : 1'b0;
  assign data_o[199] = (N1)? data_i[199] : 
                       (N0)? data_i[739] : 1'b0;
  assign data_o[198] = (N1)? data_i[198] : 
                       (N0)? data_i[738] : 1'b0;
  assign data_o[197] = (N1)? data_i[197] : 
                       (N0)? data_i[737] : 1'b0;
  assign data_o[196] = (N1)? data_i[196] : 
                       (N0)? data_i[736] : 1'b0;
  assign data_o[195] = (N1)? data_i[195] : 
                       (N0)? data_i[735] : 1'b0;
  assign data_o[194] = (N1)? data_i[194] : 
                       (N0)? data_i[734] : 1'b0;
  assign data_o[193] = (N1)? data_i[193] : 
                       (N0)? data_i[733] : 1'b0;
  assign data_o[192] = (N1)? data_i[192] : 
                       (N0)? data_i[732] : 1'b0;
  assign data_o[191] = (N1)? data_i[191] : 
                       (N0)? data_i[731] : 1'b0;
  assign data_o[190] = (N1)? data_i[190] : 
                       (N0)? data_i[730] : 1'b0;
  assign data_o[189] = (N1)? data_i[189] : 
                       (N0)? data_i[729] : 1'b0;
  assign data_o[188] = (N1)? data_i[188] : 
                       (N0)? data_i[728] : 1'b0;
  assign data_o[187] = (N1)? data_i[187] : 
                       (N0)? data_i[727] : 1'b0;
  assign data_o[186] = (N1)? data_i[186] : 
                       (N0)? data_i[726] : 1'b0;
  assign data_o[185] = (N1)? data_i[185] : 
                       (N0)? data_i[725] : 1'b0;
  assign data_o[184] = (N1)? data_i[184] : 
                       (N0)? data_i[724] : 1'b0;
  assign data_o[183] = (N1)? data_i[183] : 
                       (N0)? data_i[723] : 1'b0;
  assign data_o[182] = (N1)? data_i[182] : 
                       (N0)? data_i[722] : 1'b0;
  assign data_o[181] = (N1)? data_i[181] : 
                       (N0)? data_i[721] : 1'b0;
  assign data_o[180] = (N1)? data_i[180] : 
                       (N0)? data_i[720] : 1'b0;
  assign data_o[179] = (N1)? data_i[179] : 
                       (N0)? data_i[719] : 1'b0;
  assign data_o[178] = (N1)? data_i[178] : 
                       (N0)? data_i[718] : 1'b0;
  assign data_o[177] = (N1)? data_i[177] : 
                       (N0)? data_i[717] : 1'b0;
  assign data_o[176] = (N1)? data_i[176] : 
                       (N0)? data_i[716] : 1'b0;
  assign data_o[175] = (N1)? data_i[175] : 
                       (N0)? data_i[715] : 1'b0;
  assign data_o[174] = (N1)? data_i[174] : 
                       (N0)? data_i[714] : 1'b0;
  assign data_o[173] = (N1)? data_i[173] : 
                       (N0)? data_i[713] : 1'b0;
  assign data_o[172] = (N1)? data_i[172] : 
                       (N0)? data_i[712] : 1'b0;
  assign data_o[171] = (N1)? data_i[171] : 
                       (N0)? data_i[711] : 1'b0;
  assign data_o[170] = (N1)? data_i[170] : 
                       (N0)? data_i[710] : 1'b0;
  assign data_o[169] = (N1)? data_i[169] : 
                       (N0)? data_i[709] : 1'b0;
  assign data_o[168] = (N1)? data_i[168] : 
                       (N0)? data_i[708] : 1'b0;
  assign data_o[167] = (N1)? data_i[167] : 
                       (N0)? data_i[707] : 1'b0;
  assign data_o[166] = (N1)? data_i[166] : 
                       (N0)? data_i[706] : 1'b0;
  assign data_o[165] = (N1)? data_i[165] : 
                       (N0)? data_i[705] : 1'b0;
  assign data_o[164] = (N1)? data_i[164] : 
                       (N0)? data_i[704] : 1'b0;
  assign data_o[163] = (N1)? data_i[163] : 
                       (N0)? data_i[703] : 1'b0;
  assign data_o[162] = (N1)? data_i[162] : 
                       (N0)? data_i[702] : 1'b0;
  assign data_o[161] = (N1)? data_i[161] : 
                       (N0)? data_i[701] : 1'b0;
  assign data_o[160] = (N1)? data_i[160] : 
                       (N0)? data_i[700] : 1'b0;
  assign data_o[159] = (N1)? data_i[159] : 
                       (N0)? data_i[699] : 1'b0;
  assign data_o[158] = (N1)? data_i[158] : 
                       (N0)? data_i[698] : 1'b0;
  assign data_o[157] = (N1)? data_i[157] : 
                       (N0)? data_i[697] : 1'b0;
  assign data_o[156] = (N1)? data_i[156] : 
                       (N0)? data_i[696] : 1'b0;
  assign data_o[155] = (N1)? data_i[155] : 
                       (N0)? data_i[695] : 1'b0;
  assign data_o[154] = (N1)? data_i[154] : 
                       (N0)? data_i[694] : 1'b0;
  assign data_o[153] = (N1)? data_i[153] : 
                       (N0)? data_i[693] : 1'b0;
  assign data_o[152] = (N1)? data_i[152] : 
                       (N0)? data_i[692] : 1'b0;
  assign data_o[151] = (N1)? data_i[151] : 
                       (N0)? data_i[691] : 1'b0;
  assign data_o[150] = (N1)? data_i[150] : 
                       (N0)? data_i[690] : 1'b0;
  assign data_o[149] = (N1)? data_i[149] : 
                       (N0)? data_i[689] : 1'b0;
  assign data_o[148] = (N1)? data_i[148] : 
                       (N0)? data_i[688] : 1'b0;
  assign data_o[147] = (N1)? data_i[147] : 
                       (N0)? data_i[687] : 1'b0;
  assign data_o[146] = (N1)? data_i[146] : 
                       (N0)? data_i[686] : 1'b0;
  assign data_o[145] = (N1)? data_i[145] : 
                       (N0)? data_i[685] : 1'b0;
  assign data_o[144] = (N1)? data_i[144] : 
                       (N0)? data_i[684] : 1'b0;
  assign data_o[143] = (N1)? data_i[143] : 
                       (N0)? data_i[683] : 1'b0;
  assign data_o[142] = (N1)? data_i[142] : 
                       (N0)? data_i[682] : 1'b0;
  assign data_o[141] = (N1)? data_i[141] : 
                       (N0)? data_i[681] : 1'b0;
  assign data_o[140] = (N1)? data_i[140] : 
                       (N0)? data_i[680] : 1'b0;
  assign data_o[139] = (N1)? data_i[139] : 
                       (N0)? data_i[679] : 1'b0;
  assign data_o[138] = (N1)? data_i[138] : 
                       (N0)? data_i[678] : 1'b0;
  assign data_o[137] = (N1)? data_i[137] : 
                       (N0)? data_i[677] : 1'b0;
  assign data_o[136] = (N1)? data_i[136] : 
                       (N0)? data_i[676] : 1'b0;
  assign data_o[135] = (N1)? data_i[135] : 
                       (N0)? data_i[675] : 1'b0;
  assign data_o[134] = (N1)? data_i[134] : 
                       (N0)? data_i[674] : 1'b0;
  assign data_o[133] = (N1)? data_i[133] : 
                       (N0)? data_i[673] : 1'b0;
  assign data_o[132] = (N1)? data_i[132] : 
                       (N0)? data_i[672] : 1'b0;
  assign data_o[131] = (N1)? data_i[131] : 
                       (N0)? data_i[671] : 1'b0;
  assign data_o[130] = (N1)? data_i[130] : 
                       (N0)? data_i[670] : 1'b0;
  assign data_o[129] = (N1)? data_i[129] : 
                       (N0)? data_i[669] : 1'b0;
  assign data_o[128] = (N1)? data_i[128] : 
                       (N0)? data_i[668] : 1'b0;
  assign data_o[127] = (N1)? data_i[127] : 
                       (N0)? data_i[667] : 1'b0;
  assign data_o[126] = (N1)? data_i[126] : 
                       (N0)? data_i[666] : 1'b0;
  assign data_o[125] = (N1)? data_i[125] : 
                       (N0)? data_i[665] : 1'b0;
  assign data_o[124] = (N1)? data_i[124] : 
                       (N0)? data_i[664] : 1'b0;
  assign data_o[123] = (N1)? data_i[123] : 
                       (N0)? data_i[663] : 1'b0;
  assign data_o[122] = (N1)? data_i[122] : 
                       (N0)? data_i[662] : 1'b0;
  assign data_o[121] = (N1)? data_i[121] : 
                       (N0)? data_i[661] : 1'b0;
  assign data_o[120] = (N1)? data_i[120] : 
                       (N0)? data_i[660] : 1'b0;
  assign data_o[119] = (N1)? data_i[119] : 
                       (N0)? data_i[659] : 1'b0;
  assign data_o[118] = (N1)? data_i[118] : 
                       (N0)? data_i[658] : 1'b0;
  assign data_o[117] = (N1)? data_i[117] : 
                       (N0)? data_i[657] : 1'b0;
  assign data_o[116] = (N1)? data_i[116] : 
                       (N0)? data_i[656] : 1'b0;
  assign data_o[115] = (N1)? data_i[115] : 
                       (N0)? data_i[655] : 1'b0;
  assign data_o[114] = (N1)? data_i[114] : 
                       (N0)? data_i[654] : 1'b0;
  assign data_o[113] = (N1)? data_i[113] : 
                       (N0)? data_i[653] : 1'b0;
  assign data_o[112] = (N1)? data_i[112] : 
                       (N0)? data_i[652] : 1'b0;
  assign data_o[111] = (N1)? data_i[111] : 
                       (N0)? data_i[651] : 1'b0;
  assign data_o[110] = (N1)? data_i[110] : 
                       (N0)? data_i[650] : 1'b0;
  assign data_o[109] = (N1)? data_i[109] : 
                       (N0)? data_i[649] : 1'b0;
  assign data_o[108] = (N1)? data_i[108] : 
                       (N0)? data_i[648] : 1'b0;
  assign data_o[107] = (N1)? data_i[107] : 
                       (N0)? data_i[647] : 1'b0;
  assign data_o[106] = (N1)? data_i[106] : 
                       (N0)? data_i[646] : 1'b0;
  assign data_o[105] = (N1)? data_i[105] : 
                       (N0)? data_i[645] : 1'b0;
  assign data_o[104] = (N1)? data_i[104] : 
                       (N0)? data_i[644] : 1'b0;
  assign data_o[103] = (N1)? data_i[103] : 
                       (N0)? data_i[643] : 1'b0;
  assign data_o[102] = (N1)? data_i[102] : 
                       (N0)? data_i[642] : 1'b0;
  assign data_o[101] = (N1)? data_i[101] : 
                       (N0)? data_i[641] : 1'b0;
  assign data_o[100] = (N1)? data_i[100] : 
                       (N0)? data_i[640] : 1'b0;
  assign data_o[99] = (N1)? data_i[99] : 
                      (N0)? data_i[639] : 1'b0;
  assign data_o[98] = (N1)? data_i[98] : 
                      (N0)? data_i[638] : 1'b0;
  assign data_o[97] = (N1)? data_i[97] : 
                      (N0)? data_i[637] : 1'b0;
  assign data_o[96] = (N1)? data_i[96] : 
                      (N0)? data_i[636] : 1'b0;
  assign data_o[95] = (N1)? data_i[95] : 
                      (N0)? data_i[635] : 1'b0;
  assign data_o[94] = (N1)? data_i[94] : 
                      (N0)? data_i[634] : 1'b0;
  assign data_o[93] = (N1)? data_i[93] : 
                      (N0)? data_i[633] : 1'b0;
  assign data_o[92] = (N1)? data_i[92] : 
                      (N0)? data_i[632] : 1'b0;
  assign data_o[91] = (N1)? data_i[91] : 
                      (N0)? data_i[631] : 1'b0;
  assign data_o[90] = (N1)? data_i[90] : 
                      (N0)? data_i[630] : 1'b0;
  assign data_o[89] = (N1)? data_i[89] : 
                      (N0)? data_i[629] : 1'b0;
  assign data_o[88] = (N1)? data_i[88] : 
                      (N0)? data_i[628] : 1'b0;
  assign data_o[87] = (N1)? data_i[87] : 
                      (N0)? data_i[627] : 1'b0;
  assign data_o[86] = (N1)? data_i[86] : 
                      (N0)? data_i[626] : 1'b0;
  assign data_o[85] = (N1)? data_i[85] : 
                      (N0)? data_i[625] : 1'b0;
  assign data_o[84] = (N1)? data_i[84] : 
                      (N0)? data_i[624] : 1'b0;
  assign data_o[83] = (N1)? data_i[83] : 
                      (N0)? data_i[623] : 1'b0;
  assign data_o[82] = (N1)? data_i[82] : 
                      (N0)? data_i[622] : 1'b0;
  assign data_o[81] = (N1)? data_i[81] : 
                      (N0)? data_i[621] : 1'b0;
  assign data_o[80] = (N1)? data_i[80] : 
                      (N0)? data_i[620] : 1'b0;
  assign data_o[79] = (N1)? data_i[79] : 
                      (N0)? data_i[619] : 1'b0;
  assign data_o[78] = (N1)? data_i[78] : 
                      (N0)? data_i[618] : 1'b0;
  assign data_o[77] = (N1)? data_i[77] : 
                      (N0)? data_i[617] : 1'b0;
  assign data_o[76] = (N1)? data_i[76] : 
                      (N0)? data_i[616] : 1'b0;
  assign data_o[75] = (N1)? data_i[75] : 
                      (N0)? data_i[615] : 1'b0;
  assign data_o[74] = (N1)? data_i[74] : 
                      (N0)? data_i[614] : 1'b0;
  assign data_o[73] = (N1)? data_i[73] : 
                      (N0)? data_i[613] : 1'b0;
  assign data_o[72] = (N1)? data_i[72] : 
                      (N0)? data_i[612] : 1'b0;
  assign data_o[71] = (N1)? data_i[71] : 
                      (N0)? data_i[611] : 1'b0;
  assign data_o[70] = (N1)? data_i[70] : 
                      (N0)? data_i[610] : 1'b0;
  assign data_o[69] = (N1)? data_i[69] : 
                      (N0)? data_i[609] : 1'b0;
  assign data_o[68] = (N1)? data_i[68] : 
                      (N0)? data_i[608] : 1'b0;
  assign data_o[67] = (N1)? data_i[67] : 
                      (N0)? data_i[607] : 1'b0;
  assign data_o[66] = (N1)? data_i[66] : 
                      (N0)? data_i[606] : 1'b0;
  assign data_o[65] = (N1)? data_i[65] : 
                      (N0)? data_i[605] : 1'b0;
  assign data_o[64] = (N1)? data_i[64] : 
                      (N0)? data_i[604] : 1'b0;
  assign data_o[63] = (N1)? data_i[63] : 
                      (N0)? data_i[603] : 1'b0;
  assign data_o[62] = (N1)? data_i[62] : 
                      (N0)? data_i[602] : 1'b0;
  assign data_o[61] = (N1)? data_i[61] : 
                      (N0)? data_i[601] : 1'b0;
  assign data_o[60] = (N1)? data_i[60] : 
                      (N0)? data_i[600] : 1'b0;
  assign data_o[59] = (N1)? data_i[59] : 
                      (N0)? data_i[599] : 1'b0;
  assign data_o[58] = (N1)? data_i[58] : 
                      (N0)? data_i[598] : 1'b0;
  assign data_o[57] = (N1)? data_i[57] : 
                      (N0)? data_i[597] : 1'b0;
  assign data_o[56] = (N1)? data_i[56] : 
                      (N0)? data_i[596] : 1'b0;
  assign data_o[55] = (N1)? data_i[55] : 
                      (N0)? data_i[595] : 1'b0;
  assign data_o[54] = (N1)? data_i[54] : 
                      (N0)? data_i[594] : 1'b0;
  assign data_o[53] = (N1)? data_i[53] : 
                      (N0)? data_i[593] : 1'b0;
  assign data_o[52] = (N1)? data_i[52] : 
                      (N0)? data_i[592] : 1'b0;
  assign data_o[51] = (N1)? data_i[51] : 
                      (N0)? data_i[591] : 1'b0;
  assign data_o[50] = (N1)? data_i[50] : 
                      (N0)? data_i[590] : 1'b0;
  assign data_o[49] = (N1)? data_i[49] : 
                      (N0)? data_i[589] : 1'b0;
  assign data_o[48] = (N1)? data_i[48] : 
                      (N0)? data_i[588] : 1'b0;
  assign data_o[47] = (N1)? data_i[47] : 
                      (N0)? data_i[587] : 1'b0;
  assign data_o[46] = (N1)? data_i[46] : 
                      (N0)? data_i[586] : 1'b0;
  assign data_o[45] = (N1)? data_i[45] : 
                      (N0)? data_i[585] : 1'b0;
  assign data_o[44] = (N1)? data_i[44] : 
                      (N0)? data_i[584] : 1'b0;
  assign data_o[43] = (N1)? data_i[43] : 
                      (N0)? data_i[583] : 1'b0;
  assign data_o[42] = (N1)? data_i[42] : 
                      (N0)? data_i[582] : 1'b0;
  assign data_o[41] = (N1)? data_i[41] : 
                      (N0)? data_i[581] : 1'b0;
  assign data_o[40] = (N1)? data_i[40] : 
                      (N0)? data_i[580] : 1'b0;
  assign data_o[39] = (N1)? data_i[39] : 
                      (N0)? data_i[579] : 1'b0;
  assign data_o[38] = (N1)? data_i[38] : 
                      (N0)? data_i[578] : 1'b0;
  assign data_o[37] = (N1)? data_i[37] : 
                      (N0)? data_i[577] : 1'b0;
  assign data_o[36] = (N1)? data_i[36] : 
                      (N0)? data_i[576] : 1'b0;
  assign data_o[35] = (N1)? data_i[35] : 
                      (N0)? data_i[575] : 1'b0;
  assign data_o[34] = (N1)? data_i[34] : 
                      (N0)? data_i[574] : 1'b0;
  assign data_o[33] = (N1)? data_i[33] : 
                      (N0)? data_i[573] : 1'b0;
  assign data_o[32] = (N1)? data_i[32] : 
                      (N0)? data_i[572] : 1'b0;
  assign data_o[31] = (N1)? data_i[31] : 
                      (N0)? data_i[571] : 1'b0;
  assign data_o[30] = (N1)? data_i[30] : 
                      (N0)? data_i[570] : 1'b0;
  assign data_o[29] = (N1)? data_i[29] : 
                      (N0)? data_i[569] : 1'b0;
  assign data_o[28] = (N1)? data_i[28] : 
                      (N0)? data_i[568] : 1'b0;
  assign data_o[27] = (N1)? data_i[27] : 
                      (N0)? data_i[567] : 1'b0;
  assign data_o[26] = (N1)? data_i[26] : 
                      (N0)? data_i[566] : 1'b0;
  assign data_o[25] = (N1)? data_i[25] : 
                      (N0)? data_i[565] : 1'b0;
  assign data_o[24] = (N1)? data_i[24] : 
                      (N0)? data_i[564] : 1'b0;
  assign data_o[23] = (N1)? data_i[23] : 
                      (N0)? data_i[563] : 1'b0;
  assign data_o[22] = (N1)? data_i[22] : 
                      (N0)? data_i[562] : 1'b0;
  assign data_o[21] = (N1)? data_i[21] : 
                      (N0)? data_i[561] : 1'b0;
  assign data_o[20] = (N1)? data_i[20] : 
                      (N0)? data_i[560] : 1'b0;
  assign data_o[19] = (N1)? data_i[19] : 
                      (N0)? data_i[559] : 1'b0;
  assign data_o[18] = (N1)? data_i[18] : 
                      (N0)? data_i[558] : 1'b0;
  assign data_o[17] = (N1)? data_i[17] : 
                      (N0)? data_i[557] : 1'b0;
  assign data_o[16] = (N1)? data_i[16] : 
                      (N0)? data_i[556] : 1'b0;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[555] : 1'b0;
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[554] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[553] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[552] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[551] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[550] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[549] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[548] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[547] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[546] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[545] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[544] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[543] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[542] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[541] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[540] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_dff_reset_en_0000021d
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [540:0] data_i;
  output [540:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [540:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7;
  reg data_o_540_sv2v_reg,data_o_539_sv2v_reg,data_o_538_sv2v_reg,data_o_537_sv2v_reg,
  data_o_536_sv2v_reg,data_o_535_sv2v_reg,data_o_534_sv2v_reg,data_o_533_sv2v_reg,
  data_o_532_sv2v_reg,data_o_531_sv2v_reg,data_o_530_sv2v_reg,data_o_529_sv2v_reg,
  data_o_528_sv2v_reg,data_o_527_sv2v_reg,data_o_526_sv2v_reg,data_o_525_sv2v_reg,
  data_o_524_sv2v_reg,data_o_523_sv2v_reg,data_o_522_sv2v_reg,data_o_521_sv2v_reg,
  data_o_520_sv2v_reg,data_o_519_sv2v_reg,data_o_518_sv2v_reg,data_o_517_sv2v_reg,
  data_o_516_sv2v_reg,data_o_515_sv2v_reg,data_o_514_sv2v_reg,data_o_513_sv2v_reg,
  data_o_512_sv2v_reg,data_o_511_sv2v_reg,data_o_510_sv2v_reg,data_o_509_sv2v_reg,
  data_o_508_sv2v_reg,data_o_507_sv2v_reg,data_o_506_sv2v_reg,data_o_505_sv2v_reg,
  data_o_504_sv2v_reg,data_o_503_sv2v_reg,data_o_502_sv2v_reg,data_o_501_sv2v_reg,
  data_o_500_sv2v_reg,data_o_499_sv2v_reg,data_o_498_sv2v_reg,data_o_497_sv2v_reg,
  data_o_496_sv2v_reg,data_o_495_sv2v_reg,data_o_494_sv2v_reg,data_o_493_sv2v_reg,
  data_o_492_sv2v_reg,data_o_491_sv2v_reg,data_o_490_sv2v_reg,data_o_489_sv2v_reg,
  data_o_488_sv2v_reg,data_o_487_sv2v_reg,data_o_486_sv2v_reg,data_o_485_sv2v_reg,
  data_o_484_sv2v_reg,data_o_483_sv2v_reg,data_o_482_sv2v_reg,data_o_481_sv2v_reg,
  data_o_480_sv2v_reg,data_o_479_sv2v_reg,data_o_478_sv2v_reg,data_o_477_sv2v_reg,
  data_o_476_sv2v_reg,data_o_475_sv2v_reg,data_o_474_sv2v_reg,data_o_473_sv2v_reg,
  data_o_472_sv2v_reg,data_o_471_sv2v_reg,data_o_470_sv2v_reg,data_o_469_sv2v_reg,
  data_o_468_sv2v_reg,data_o_467_sv2v_reg,data_o_466_sv2v_reg,data_o_465_sv2v_reg,
  data_o_464_sv2v_reg,data_o_463_sv2v_reg,data_o_462_sv2v_reg,data_o_461_sv2v_reg,
  data_o_460_sv2v_reg,data_o_459_sv2v_reg,data_o_458_sv2v_reg,data_o_457_sv2v_reg,
  data_o_456_sv2v_reg,data_o_455_sv2v_reg,data_o_454_sv2v_reg,data_o_453_sv2v_reg,
  data_o_452_sv2v_reg,data_o_451_sv2v_reg,data_o_450_sv2v_reg,data_o_449_sv2v_reg,
  data_o_448_sv2v_reg,data_o_447_sv2v_reg,data_o_446_sv2v_reg,data_o_445_sv2v_reg,
  data_o_444_sv2v_reg,data_o_443_sv2v_reg,data_o_442_sv2v_reg,data_o_441_sv2v_reg,
  data_o_440_sv2v_reg,data_o_439_sv2v_reg,data_o_438_sv2v_reg,data_o_437_sv2v_reg,
  data_o_436_sv2v_reg,data_o_435_sv2v_reg,data_o_434_sv2v_reg,data_o_433_sv2v_reg,
  data_o_432_sv2v_reg,data_o_431_sv2v_reg,data_o_430_sv2v_reg,data_o_429_sv2v_reg,
  data_o_428_sv2v_reg,data_o_427_sv2v_reg,data_o_426_sv2v_reg,data_o_425_sv2v_reg,
  data_o_424_sv2v_reg,data_o_423_sv2v_reg,data_o_422_sv2v_reg,data_o_421_sv2v_reg,
  data_o_420_sv2v_reg,data_o_419_sv2v_reg,data_o_418_sv2v_reg,data_o_417_sv2v_reg,
  data_o_416_sv2v_reg,data_o_415_sv2v_reg,data_o_414_sv2v_reg,data_o_413_sv2v_reg,
  data_o_412_sv2v_reg,data_o_411_sv2v_reg,data_o_410_sv2v_reg,data_o_409_sv2v_reg,
  data_o_408_sv2v_reg,data_o_407_sv2v_reg,data_o_406_sv2v_reg,data_o_405_sv2v_reg,
  data_o_404_sv2v_reg,data_o_403_sv2v_reg,data_o_402_sv2v_reg,data_o_401_sv2v_reg,
  data_o_400_sv2v_reg,data_o_399_sv2v_reg,data_o_398_sv2v_reg,data_o_397_sv2v_reg,
  data_o_396_sv2v_reg,data_o_395_sv2v_reg,data_o_394_sv2v_reg,data_o_393_sv2v_reg,
  data_o_392_sv2v_reg,data_o_391_sv2v_reg,data_o_390_sv2v_reg,data_o_389_sv2v_reg,
  data_o_388_sv2v_reg,data_o_387_sv2v_reg,data_o_386_sv2v_reg,data_o_385_sv2v_reg,
  data_o_384_sv2v_reg,data_o_383_sv2v_reg,data_o_382_sv2v_reg,data_o_381_sv2v_reg,
  data_o_380_sv2v_reg,data_o_379_sv2v_reg,data_o_378_sv2v_reg,data_o_377_sv2v_reg,
  data_o_376_sv2v_reg,data_o_375_sv2v_reg,data_o_374_sv2v_reg,data_o_373_sv2v_reg,
  data_o_372_sv2v_reg,data_o_371_sv2v_reg,data_o_370_sv2v_reg,data_o_369_sv2v_reg,
  data_o_368_sv2v_reg,data_o_367_sv2v_reg,data_o_366_sv2v_reg,data_o_365_sv2v_reg,
  data_o_364_sv2v_reg,data_o_363_sv2v_reg,data_o_362_sv2v_reg,data_o_361_sv2v_reg,
  data_o_360_sv2v_reg,data_o_359_sv2v_reg,data_o_358_sv2v_reg,data_o_357_sv2v_reg,
  data_o_356_sv2v_reg,data_o_355_sv2v_reg,data_o_354_sv2v_reg,data_o_353_sv2v_reg,
  data_o_352_sv2v_reg,data_o_351_sv2v_reg,data_o_350_sv2v_reg,data_o_349_sv2v_reg,
  data_o_348_sv2v_reg,data_o_347_sv2v_reg,data_o_346_sv2v_reg,data_o_345_sv2v_reg,
  data_o_344_sv2v_reg,data_o_343_sv2v_reg,data_o_342_sv2v_reg,data_o_341_sv2v_reg,
  data_o_340_sv2v_reg,data_o_339_sv2v_reg,data_o_338_sv2v_reg,data_o_337_sv2v_reg,
  data_o_336_sv2v_reg,data_o_335_sv2v_reg,data_o_334_sv2v_reg,data_o_333_sv2v_reg,
  data_o_332_sv2v_reg,data_o_331_sv2v_reg,data_o_330_sv2v_reg,data_o_329_sv2v_reg,
  data_o_328_sv2v_reg,data_o_327_sv2v_reg,data_o_326_sv2v_reg,data_o_325_sv2v_reg,
  data_o_324_sv2v_reg,data_o_323_sv2v_reg,data_o_322_sv2v_reg,data_o_321_sv2v_reg,
  data_o_320_sv2v_reg,data_o_319_sv2v_reg,data_o_318_sv2v_reg,data_o_317_sv2v_reg,
  data_o_316_sv2v_reg,data_o_315_sv2v_reg,data_o_314_sv2v_reg,data_o_313_sv2v_reg,
  data_o_312_sv2v_reg,data_o_311_sv2v_reg,data_o_310_sv2v_reg,data_o_309_sv2v_reg,
  data_o_308_sv2v_reg,data_o_307_sv2v_reg,data_o_306_sv2v_reg,data_o_305_sv2v_reg,
  data_o_304_sv2v_reg,data_o_303_sv2v_reg,data_o_302_sv2v_reg,data_o_301_sv2v_reg,
  data_o_300_sv2v_reg,data_o_299_sv2v_reg,data_o_298_sv2v_reg,data_o_297_sv2v_reg,
  data_o_296_sv2v_reg,data_o_295_sv2v_reg,data_o_294_sv2v_reg,data_o_293_sv2v_reg,
  data_o_292_sv2v_reg,data_o_291_sv2v_reg,data_o_290_sv2v_reg,data_o_289_sv2v_reg,
  data_o_288_sv2v_reg,data_o_287_sv2v_reg,data_o_286_sv2v_reg,data_o_285_sv2v_reg,
  data_o_284_sv2v_reg,data_o_283_sv2v_reg,data_o_282_sv2v_reg,data_o_281_sv2v_reg,
  data_o_280_sv2v_reg,data_o_279_sv2v_reg,data_o_278_sv2v_reg,data_o_277_sv2v_reg,
  data_o_276_sv2v_reg,data_o_275_sv2v_reg,data_o_274_sv2v_reg,data_o_273_sv2v_reg,
  data_o_272_sv2v_reg,data_o_271_sv2v_reg,data_o_270_sv2v_reg,data_o_269_sv2v_reg,
  data_o_268_sv2v_reg,data_o_267_sv2v_reg,data_o_266_sv2v_reg,data_o_265_sv2v_reg,
  data_o_264_sv2v_reg,data_o_263_sv2v_reg,data_o_262_sv2v_reg,data_o_261_sv2v_reg,
  data_o_260_sv2v_reg,data_o_259_sv2v_reg,data_o_258_sv2v_reg,data_o_257_sv2v_reg,
  data_o_256_sv2v_reg,data_o_255_sv2v_reg,data_o_254_sv2v_reg,data_o_253_sv2v_reg,
  data_o_252_sv2v_reg,data_o_251_sv2v_reg,data_o_250_sv2v_reg,data_o_249_sv2v_reg,
  data_o_248_sv2v_reg,data_o_247_sv2v_reg,data_o_246_sv2v_reg,data_o_245_sv2v_reg,
  data_o_244_sv2v_reg,data_o_243_sv2v_reg,data_o_242_sv2v_reg,data_o_241_sv2v_reg,
  data_o_240_sv2v_reg,data_o_239_sv2v_reg,data_o_238_sv2v_reg,data_o_237_sv2v_reg,
  data_o_236_sv2v_reg,data_o_235_sv2v_reg,data_o_234_sv2v_reg,data_o_233_sv2v_reg,
  data_o_232_sv2v_reg,data_o_231_sv2v_reg,data_o_230_sv2v_reg,data_o_229_sv2v_reg,
  data_o_228_sv2v_reg,data_o_227_sv2v_reg,data_o_226_sv2v_reg,data_o_225_sv2v_reg,
  data_o_224_sv2v_reg,data_o_223_sv2v_reg,data_o_222_sv2v_reg,data_o_221_sv2v_reg,
  data_o_220_sv2v_reg,data_o_219_sv2v_reg,data_o_218_sv2v_reg,data_o_217_sv2v_reg,
  data_o_216_sv2v_reg,data_o_215_sv2v_reg,data_o_214_sv2v_reg,data_o_213_sv2v_reg,
  data_o_212_sv2v_reg,data_o_211_sv2v_reg,data_o_210_sv2v_reg,data_o_209_sv2v_reg,
  data_o_208_sv2v_reg,data_o_207_sv2v_reg,data_o_206_sv2v_reg,data_o_205_sv2v_reg,
  data_o_204_sv2v_reg,data_o_203_sv2v_reg,data_o_202_sv2v_reg,data_o_201_sv2v_reg,
  data_o_200_sv2v_reg,data_o_199_sv2v_reg,data_o_198_sv2v_reg,data_o_197_sv2v_reg,
  data_o_196_sv2v_reg,data_o_195_sv2v_reg,data_o_194_sv2v_reg,data_o_193_sv2v_reg,
  data_o_192_sv2v_reg,data_o_191_sv2v_reg,data_o_190_sv2v_reg,data_o_189_sv2v_reg,
  data_o_188_sv2v_reg,data_o_187_sv2v_reg,data_o_186_sv2v_reg,data_o_185_sv2v_reg,
  data_o_184_sv2v_reg,data_o_183_sv2v_reg,data_o_182_sv2v_reg,data_o_181_sv2v_reg,
  data_o_180_sv2v_reg,data_o_179_sv2v_reg,data_o_178_sv2v_reg,data_o_177_sv2v_reg,
  data_o_176_sv2v_reg,data_o_175_sv2v_reg,data_o_174_sv2v_reg,data_o_173_sv2v_reg,
  data_o_172_sv2v_reg,data_o_171_sv2v_reg,data_o_170_sv2v_reg,data_o_169_sv2v_reg,
  data_o_168_sv2v_reg,data_o_167_sv2v_reg,data_o_166_sv2v_reg,data_o_165_sv2v_reg,
  data_o_164_sv2v_reg,data_o_163_sv2v_reg,data_o_162_sv2v_reg,data_o_161_sv2v_reg,
  data_o_160_sv2v_reg,data_o_159_sv2v_reg,data_o_158_sv2v_reg,data_o_157_sv2v_reg,
  data_o_156_sv2v_reg,data_o_155_sv2v_reg,data_o_154_sv2v_reg,data_o_153_sv2v_reg,
  data_o_152_sv2v_reg,data_o_151_sv2v_reg,data_o_150_sv2v_reg,data_o_149_sv2v_reg,
  data_o_148_sv2v_reg,data_o_147_sv2v_reg,data_o_146_sv2v_reg,data_o_145_sv2v_reg,
  data_o_144_sv2v_reg,data_o_143_sv2v_reg,data_o_142_sv2v_reg,data_o_141_sv2v_reg,
  data_o_140_sv2v_reg,data_o_139_sv2v_reg,data_o_138_sv2v_reg,data_o_137_sv2v_reg,
  data_o_136_sv2v_reg,data_o_135_sv2v_reg,data_o_134_sv2v_reg,data_o_133_sv2v_reg,
  data_o_132_sv2v_reg,data_o_131_sv2v_reg,data_o_130_sv2v_reg,data_o_129_sv2v_reg,
  data_o_128_sv2v_reg,data_o_127_sv2v_reg,data_o_126_sv2v_reg,data_o_125_sv2v_reg,
  data_o_124_sv2v_reg,data_o_123_sv2v_reg,data_o_122_sv2v_reg,data_o_121_sv2v_reg,
  data_o_120_sv2v_reg,data_o_119_sv2v_reg,data_o_118_sv2v_reg,data_o_117_sv2v_reg,
  data_o_116_sv2v_reg,data_o_115_sv2v_reg,data_o_114_sv2v_reg,data_o_113_sv2v_reg,
  data_o_112_sv2v_reg,data_o_111_sv2v_reg,data_o_110_sv2v_reg,data_o_109_sv2v_reg,
  data_o_108_sv2v_reg,data_o_107_sv2v_reg,data_o_106_sv2v_reg,data_o_105_sv2v_reg,
  data_o_104_sv2v_reg,data_o_103_sv2v_reg,data_o_102_sv2v_reg,data_o_101_sv2v_reg,
  data_o_100_sv2v_reg,data_o_99_sv2v_reg,data_o_98_sv2v_reg,data_o_97_sv2v_reg,
  data_o_96_sv2v_reg,data_o_95_sv2v_reg,data_o_94_sv2v_reg,data_o_93_sv2v_reg,
  data_o_92_sv2v_reg,data_o_91_sv2v_reg,data_o_90_sv2v_reg,data_o_89_sv2v_reg,
  data_o_88_sv2v_reg,data_o_87_sv2v_reg,data_o_86_sv2v_reg,data_o_85_sv2v_reg,
  data_o_84_sv2v_reg,data_o_83_sv2v_reg,data_o_82_sv2v_reg,data_o_81_sv2v_reg,data_o_80_sv2v_reg,
  data_o_79_sv2v_reg,data_o_78_sv2v_reg,data_o_77_sv2v_reg,data_o_76_sv2v_reg,
  data_o_75_sv2v_reg,data_o_74_sv2v_reg,data_o_73_sv2v_reg,data_o_72_sv2v_reg,
  data_o_71_sv2v_reg,data_o_70_sv2v_reg,data_o_69_sv2v_reg,data_o_68_sv2v_reg,
  data_o_67_sv2v_reg,data_o_66_sv2v_reg,data_o_65_sv2v_reg,data_o_64_sv2v_reg,
  data_o_63_sv2v_reg,data_o_62_sv2v_reg,data_o_61_sv2v_reg,data_o_60_sv2v_reg,data_o_59_sv2v_reg,
  data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,data_o_55_sv2v_reg,
  data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,data_o_51_sv2v_reg,
  data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,data_o_47_sv2v_reg,
  data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,data_o_43_sv2v_reg,
  data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,
  data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,
  data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,
  data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,
  data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,
  data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,
  data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,
  data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,
  data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[540] = data_o_540_sv2v_reg;
  assign data_o[539] = data_o_539_sv2v_reg;
  assign data_o[538] = data_o_538_sv2v_reg;
  assign data_o[537] = data_o_537_sv2v_reg;
  assign data_o[536] = data_o_536_sv2v_reg;
  assign data_o[535] = data_o_535_sv2v_reg;
  assign data_o[534] = data_o_534_sv2v_reg;
  assign data_o[533] = data_o_533_sv2v_reg;
  assign data_o[532] = data_o_532_sv2v_reg;
  assign data_o[531] = data_o_531_sv2v_reg;
  assign data_o[530] = data_o_530_sv2v_reg;
  assign data_o[529] = data_o_529_sv2v_reg;
  assign data_o[528] = data_o_528_sv2v_reg;
  assign data_o[527] = data_o_527_sv2v_reg;
  assign data_o[526] = data_o_526_sv2v_reg;
  assign data_o[525] = data_o_525_sv2v_reg;
  assign data_o[524] = data_o_524_sv2v_reg;
  assign data_o[523] = data_o_523_sv2v_reg;
  assign data_o[522] = data_o_522_sv2v_reg;
  assign data_o[521] = data_o_521_sv2v_reg;
  assign data_o[520] = data_o_520_sv2v_reg;
  assign data_o[519] = data_o_519_sv2v_reg;
  assign data_o[518] = data_o_518_sv2v_reg;
  assign data_o[517] = data_o_517_sv2v_reg;
  assign data_o[516] = data_o_516_sv2v_reg;
  assign data_o[515] = data_o_515_sv2v_reg;
  assign data_o[514] = data_o_514_sv2v_reg;
  assign data_o[513] = data_o_513_sv2v_reg;
  assign data_o[512] = data_o_512_sv2v_reg;
  assign data_o[511] = data_o_511_sv2v_reg;
  assign data_o[510] = data_o_510_sv2v_reg;
  assign data_o[509] = data_o_509_sv2v_reg;
  assign data_o[508] = data_o_508_sv2v_reg;
  assign data_o[507] = data_o_507_sv2v_reg;
  assign data_o[506] = data_o_506_sv2v_reg;
  assign data_o[505] = data_o_505_sv2v_reg;
  assign data_o[504] = data_o_504_sv2v_reg;
  assign data_o[503] = data_o_503_sv2v_reg;
  assign data_o[502] = data_o_502_sv2v_reg;
  assign data_o[501] = data_o_501_sv2v_reg;
  assign data_o[500] = data_o_500_sv2v_reg;
  assign data_o[499] = data_o_499_sv2v_reg;
  assign data_o[498] = data_o_498_sv2v_reg;
  assign data_o[497] = data_o_497_sv2v_reg;
  assign data_o[496] = data_o_496_sv2v_reg;
  assign data_o[495] = data_o_495_sv2v_reg;
  assign data_o[494] = data_o_494_sv2v_reg;
  assign data_o[493] = data_o_493_sv2v_reg;
  assign data_o[492] = data_o_492_sv2v_reg;
  assign data_o[491] = data_o_491_sv2v_reg;
  assign data_o[490] = data_o_490_sv2v_reg;
  assign data_o[489] = data_o_489_sv2v_reg;
  assign data_o[488] = data_o_488_sv2v_reg;
  assign data_o[487] = data_o_487_sv2v_reg;
  assign data_o[486] = data_o_486_sv2v_reg;
  assign data_o[485] = data_o_485_sv2v_reg;
  assign data_o[484] = data_o_484_sv2v_reg;
  assign data_o[483] = data_o_483_sv2v_reg;
  assign data_o[482] = data_o_482_sv2v_reg;
  assign data_o[481] = data_o_481_sv2v_reg;
  assign data_o[480] = data_o_480_sv2v_reg;
  assign data_o[479] = data_o_479_sv2v_reg;
  assign data_o[478] = data_o_478_sv2v_reg;
  assign data_o[477] = data_o_477_sv2v_reg;
  assign data_o[476] = data_o_476_sv2v_reg;
  assign data_o[475] = data_o_475_sv2v_reg;
  assign data_o[474] = data_o_474_sv2v_reg;
  assign data_o[473] = data_o_473_sv2v_reg;
  assign data_o[472] = data_o_472_sv2v_reg;
  assign data_o[471] = data_o_471_sv2v_reg;
  assign data_o[470] = data_o_470_sv2v_reg;
  assign data_o[469] = data_o_469_sv2v_reg;
  assign data_o[468] = data_o_468_sv2v_reg;
  assign data_o[467] = data_o_467_sv2v_reg;
  assign data_o[466] = data_o_466_sv2v_reg;
  assign data_o[465] = data_o_465_sv2v_reg;
  assign data_o[464] = data_o_464_sv2v_reg;
  assign data_o[463] = data_o_463_sv2v_reg;
  assign data_o[462] = data_o_462_sv2v_reg;
  assign data_o[461] = data_o_461_sv2v_reg;
  assign data_o[460] = data_o_460_sv2v_reg;
  assign data_o[459] = data_o_459_sv2v_reg;
  assign data_o[458] = data_o_458_sv2v_reg;
  assign data_o[457] = data_o_457_sv2v_reg;
  assign data_o[456] = data_o_456_sv2v_reg;
  assign data_o[455] = data_o_455_sv2v_reg;
  assign data_o[454] = data_o_454_sv2v_reg;
  assign data_o[453] = data_o_453_sv2v_reg;
  assign data_o[452] = data_o_452_sv2v_reg;
  assign data_o[451] = data_o_451_sv2v_reg;
  assign data_o[450] = data_o_450_sv2v_reg;
  assign data_o[449] = data_o_449_sv2v_reg;
  assign data_o[448] = data_o_448_sv2v_reg;
  assign data_o[447] = data_o_447_sv2v_reg;
  assign data_o[446] = data_o_446_sv2v_reg;
  assign data_o[445] = data_o_445_sv2v_reg;
  assign data_o[444] = data_o_444_sv2v_reg;
  assign data_o[443] = data_o_443_sv2v_reg;
  assign data_o[442] = data_o_442_sv2v_reg;
  assign data_o[441] = data_o_441_sv2v_reg;
  assign data_o[440] = data_o_440_sv2v_reg;
  assign data_o[439] = data_o_439_sv2v_reg;
  assign data_o[438] = data_o_438_sv2v_reg;
  assign data_o[437] = data_o_437_sv2v_reg;
  assign data_o[436] = data_o_436_sv2v_reg;
  assign data_o[435] = data_o_435_sv2v_reg;
  assign data_o[434] = data_o_434_sv2v_reg;
  assign data_o[433] = data_o_433_sv2v_reg;
  assign data_o[432] = data_o_432_sv2v_reg;
  assign data_o[431] = data_o_431_sv2v_reg;
  assign data_o[430] = data_o_430_sv2v_reg;
  assign data_o[429] = data_o_429_sv2v_reg;
  assign data_o[428] = data_o_428_sv2v_reg;
  assign data_o[427] = data_o_427_sv2v_reg;
  assign data_o[426] = data_o_426_sv2v_reg;
  assign data_o[425] = data_o_425_sv2v_reg;
  assign data_o[424] = data_o_424_sv2v_reg;
  assign data_o[423] = data_o_423_sv2v_reg;
  assign data_o[422] = data_o_422_sv2v_reg;
  assign data_o[421] = data_o_421_sv2v_reg;
  assign data_o[420] = data_o_420_sv2v_reg;
  assign data_o[419] = data_o_419_sv2v_reg;
  assign data_o[418] = data_o_418_sv2v_reg;
  assign data_o[417] = data_o_417_sv2v_reg;
  assign data_o[416] = data_o_416_sv2v_reg;
  assign data_o[415] = data_o_415_sv2v_reg;
  assign data_o[414] = data_o_414_sv2v_reg;
  assign data_o[413] = data_o_413_sv2v_reg;
  assign data_o[412] = data_o_412_sv2v_reg;
  assign data_o[411] = data_o_411_sv2v_reg;
  assign data_o[410] = data_o_410_sv2v_reg;
  assign data_o[409] = data_o_409_sv2v_reg;
  assign data_o[408] = data_o_408_sv2v_reg;
  assign data_o[407] = data_o_407_sv2v_reg;
  assign data_o[406] = data_o_406_sv2v_reg;
  assign data_o[405] = data_o_405_sv2v_reg;
  assign data_o[404] = data_o_404_sv2v_reg;
  assign data_o[403] = data_o_403_sv2v_reg;
  assign data_o[402] = data_o_402_sv2v_reg;
  assign data_o[401] = data_o_401_sv2v_reg;
  assign data_o[400] = data_o_400_sv2v_reg;
  assign data_o[399] = data_o_399_sv2v_reg;
  assign data_o[398] = data_o_398_sv2v_reg;
  assign data_o[397] = data_o_397_sv2v_reg;
  assign data_o[396] = data_o_396_sv2v_reg;
  assign data_o[395] = data_o_395_sv2v_reg;
  assign data_o[394] = data_o_394_sv2v_reg;
  assign data_o[393] = data_o_393_sv2v_reg;
  assign data_o[392] = data_o_392_sv2v_reg;
  assign data_o[391] = data_o_391_sv2v_reg;
  assign data_o[390] = data_o_390_sv2v_reg;
  assign data_o[389] = data_o_389_sv2v_reg;
  assign data_o[388] = data_o_388_sv2v_reg;
  assign data_o[387] = data_o_387_sv2v_reg;
  assign data_o[386] = data_o_386_sv2v_reg;
  assign data_o[385] = data_o_385_sv2v_reg;
  assign data_o[384] = data_o_384_sv2v_reg;
  assign data_o[383] = data_o_383_sv2v_reg;
  assign data_o[382] = data_o_382_sv2v_reg;
  assign data_o[381] = data_o_381_sv2v_reg;
  assign data_o[380] = data_o_380_sv2v_reg;
  assign data_o[379] = data_o_379_sv2v_reg;
  assign data_o[378] = data_o_378_sv2v_reg;
  assign data_o[377] = data_o_377_sv2v_reg;
  assign data_o[376] = data_o_376_sv2v_reg;
  assign data_o[375] = data_o_375_sv2v_reg;
  assign data_o[374] = data_o_374_sv2v_reg;
  assign data_o[373] = data_o_373_sv2v_reg;
  assign data_o[372] = data_o_372_sv2v_reg;
  assign data_o[371] = data_o_371_sv2v_reg;
  assign data_o[370] = data_o_370_sv2v_reg;
  assign data_o[369] = data_o_369_sv2v_reg;
  assign data_o[368] = data_o_368_sv2v_reg;
  assign data_o[367] = data_o_367_sv2v_reg;
  assign data_o[366] = data_o_366_sv2v_reg;
  assign data_o[365] = data_o_365_sv2v_reg;
  assign data_o[364] = data_o_364_sv2v_reg;
  assign data_o[363] = data_o_363_sv2v_reg;
  assign data_o[362] = data_o_362_sv2v_reg;
  assign data_o[361] = data_o_361_sv2v_reg;
  assign data_o[360] = data_o_360_sv2v_reg;
  assign data_o[359] = data_o_359_sv2v_reg;
  assign data_o[358] = data_o_358_sv2v_reg;
  assign data_o[357] = data_o_357_sv2v_reg;
  assign data_o[356] = data_o_356_sv2v_reg;
  assign data_o[355] = data_o_355_sv2v_reg;
  assign data_o[354] = data_o_354_sv2v_reg;
  assign data_o[353] = data_o_353_sv2v_reg;
  assign data_o[352] = data_o_352_sv2v_reg;
  assign data_o[351] = data_o_351_sv2v_reg;
  assign data_o[350] = data_o_350_sv2v_reg;
  assign data_o[349] = data_o_349_sv2v_reg;
  assign data_o[348] = data_o_348_sv2v_reg;
  assign data_o[347] = data_o_347_sv2v_reg;
  assign data_o[346] = data_o_346_sv2v_reg;
  assign data_o[345] = data_o_345_sv2v_reg;
  assign data_o[344] = data_o_344_sv2v_reg;
  assign data_o[343] = data_o_343_sv2v_reg;
  assign data_o[342] = data_o_342_sv2v_reg;
  assign data_o[341] = data_o_341_sv2v_reg;
  assign data_o[340] = data_o_340_sv2v_reg;
  assign data_o[339] = data_o_339_sv2v_reg;
  assign data_o[338] = data_o_338_sv2v_reg;
  assign data_o[337] = data_o_337_sv2v_reg;
  assign data_o[336] = data_o_336_sv2v_reg;
  assign data_o[335] = data_o_335_sv2v_reg;
  assign data_o[334] = data_o_334_sv2v_reg;
  assign data_o[333] = data_o_333_sv2v_reg;
  assign data_o[332] = data_o_332_sv2v_reg;
  assign data_o[331] = data_o_331_sv2v_reg;
  assign data_o[330] = data_o_330_sv2v_reg;
  assign data_o[329] = data_o_329_sv2v_reg;
  assign data_o[328] = data_o_328_sv2v_reg;
  assign data_o[327] = data_o_327_sv2v_reg;
  assign data_o[326] = data_o_326_sv2v_reg;
  assign data_o[325] = data_o_325_sv2v_reg;
  assign data_o[324] = data_o_324_sv2v_reg;
  assign data_o[323] = data_o_323_sv2v_reg;
  assign data_o[322] = data_o_322_sv2v_reg;
  assign data_o[321] = data_o_321_sv2v_reg;
  assign data_o[320] = data_o_320_sv2v_reg;
  assign data_o[319] = data_o_319_sv2v_reg;
  assign data_o[318] = data_o_318_sv2v_reg;
  assign data_o[317] = data_o_317_sv2v_reg;
  assign data_o[316] = data_o_316_sv2v_reg;
  assign data_o[315] = data_o_315_sv2v_reg;
  assign data_o[314] = data_o_314_sv2v_reg;
  assign data_o[313] = data_o_313_sv2v_reg;
  assign data_o[312] = data_o_312_sv2v_reg;
  assign data_o[311] = data_o_311_sv2v_reg;
  assign data_o[310] = data_o_310_sv2v_reg;
  assign data_o[309] = data_o_309_sv2v_reg;
  assign data_o[308] = data_o_308_sv2v_reg;
  assign data_o[307] = data_o_307_sv2v_reg;
  assign data_o[306] = data_o_306_sv2v_reg;
  assign data_o[305] = data_o_305_sv2v_reg;
  assign data_o[304] = data_o_304_sv2v_reg;
  assign data_o[303] = data_o_303_sv2v_reg;
  assign data_o[302] = data_o_302_sv2v_reg;
  assign data_o[301] = data_o_301_sv2v_reg;
  assign data_o[300] = data_o_300_sv2v_reg;
  assign data_o[299] = data_o_299_sv2v_reg;
  assign data_o[298] = data_o_298_sv2v_reg;
  assign data_o[297] = data_o_297_sv2v_reg;
  assign data_o[296] = data_o_296_sv2v_reg;
  assign data_o[295] = data_o_295_sv2v_reg;
  assign data_o[294] = data_o_294_sv2v_reg;
  assign data_o[293] = data_o_293_sv2v_reg;
  assign data_o[292] = data_o_292_sv2v_reg;
  assign data_o[291] = data_o_291_sv2v_reg;
  assign data_o[290] = data_o_290_sv2v_reg;
  assign data_o[289] = data_o_289_sv2v_reg;
  assign data_o[288] = data_o_288_sv2v_reg;
  assign data_o[287] = data_o_287_sv2v_reg;
  assign data_o[286] = data_o_286_sv2v_reg;
  assign data_o[285] = data_o_285_sv2v_reg;
  assign data_o[284] = data_o_284_sv2v_reg;
  assign data_o[283] = data_o_283_sv2v_reg;
  assign data_o[282] = data_o_282_sv2v_reg;
  assign data_o[281] = data_o_281_sv2v_reg;
  assign data_o[280] = data_o_280_sv2v_reg;
  assign data_o[279] = data_o_279_sv2v_reg;
  assign data_o[278] = data_o_278_sv2v_reg;
  assign data_o[277] = data_o_277_sv2v_reg;
  assign data_o[276] = data_o_276_sv2v_reg;
  assign data_o[275] = data_o_275_sv2v_reg;
  assign data_o[274] = data_o_274_sv2v_reg;
  assign data_o[273] = data_o_273_sv2v_reg;
  assign data_o[272] = data_o_272_sv2v_reg;
  assign data_o[271] = data_o_271_sv2v_reg;
  assign data_o[270] = data_o_270_sv2v_reg;
  assign data_o[269] = data_o_269_sv2v_reg;
  assign data_o[268] = data_o_268_sv2v_reg;
  assign data_o[267] = data_o_267_sv2v_reg;
  assign data_o[266] = data_o_266_sv2v_reg;
  assign data_o[265] = data_o_265_sv2v_reg;
  assign data_o[264] = data_o_264_sv2v_reg;
  assign data_o[263] = data_o_263_sv2v_reg;
  assign data_o[262] = data_o_262_sv2v_reg;
  assign data_o[261] = data_o_261_sv2v_reg;
  assign data_o[260] = data_o_260_sv2v_reg;
  assign data_o[259] = data_o_259_sv2v_reg;
  assign data_o[258] = data_o_258_sv2v_reg;
  assign data_o[257] = data_o_257_sv2v_reg;
  assign data_o[256] = data_o_256_sv2v_reg;
  assign data_o[255] = data_o_255_sv2v_reg;
  assign data_o[254] = data_o_254_sv2v_reg;
  assign data_o[253] = data_o_253_sv2v_reg;
  assign data_o[252] = data_o_252_sv2v_reg;
  assign data_o[251] = data_o_251_sv2v_reg;
  assign data_o[250] = data_o_250_sv2v_reg;
  assign data_o[249] = data_o_249_sv2v_reg;
  assign data_o[248] = data_o_248_sv2v_reg;
  assign data_o[247] = data_o_247_sv2v_reg;
  assign data_o[246] = data_o_246_sv2v_reg;
  assign data_o[245] = data_o_245_sv2v_reg;
  assign data_o[244] = data_o_244_sv2v_reg;
  assign data_o[243] = data_o_243_sv2v_reg;
  assign data_o[242] = data_o_242_sv2v_reg;
  assign data_o[241] = data_o_241_sv2v_reg;
  assign data_o[240] = data_o_240_sv2v_reg;
  assign data_o[239] = data_o_239_sv2v_reg;
  assign data_o[238] = data_o_238_sv2v_reg;
  assign data_o[237] = data_o_237_sv2v_reg;
  assign data_o[236] = data_o_236_sv2v_reg;
  assign data_o[235] = data_o_235_sv2v_reg;
  assign data_o[234] = data_o_234_sv2v_reg;
  assign data_o[233] = data_o_233_sv2v_reg;
  assign data_o[232] = data_o_232_sv2v_reg;
  assign data_o[231] = data_o_231_sv2v_reg;
  assign data_o[230] = data_o_230_sv2v_reg;
  assign data_o[229] = data_o_229_sv2v_reg;
  assign data_o[228] = data_o_228_sv2v_reg;
  assign data_o[227] = data_o_227_sv2v_reg;
  assign data_o[226] = data_o_226_sv2v_reg;
  assign data_o[225] = data_o_225_sv2v_reg;
  assign data_o[224] = data_o_224_sv2v_reg;
  assign data_o[223] = data_o_223_sv2v_reg;
  assign data_o[222] = data_o_222_sv2v_reg;
  assign data_o[221] = data_o_221_sv2v_reg;
  assign data_o[220] = data_o_220_sv2v_reg;
  assign data_o[219] = data_o_219_sv2v_reg;
  assign data_o[218] = data_o_218_sv2v_reg;
  assign data_o[217] = data_o_217_sv2v_reg;
  assign data_o[216] = data_o_216_sv2v_reg;
  assign data_o[215] = data_o_215_sv2v_reg;
  assign data_o[214] = data_o_214_sv2v_reg;
  assign data_o[213] = data_o_213_sv2v_reg;
  assign data_o[212] = data_o_212_sv2v_reg;
  assign data_o[211] = data_o_211_sv2v_reg;
  assign data_o[210] = data_o_210_sv2v_reg;
  assign data_o[209] = data_o_209_sv2v_reg;
  assign data_o[208] = data_o_208_sv2v_reg;
  assign data_o[207] = data_o_207_sv2v_reg;
  assign data_o[206] = data_o_206_sv2v_reg;
  assign data_o[205] = data_o_205_sv2v_reg;
  assign data_o[204] = data_o_204_sv2v_reg;
  assign data_o[203] = data_o_203_sv2v_reg;
  assign data_o[202] = data_o_202_sv2v_reg;
  assign data_o[201] = data_o_201_sv2v_reg;
  assign data_o[200] = data_o_200_sv2v_reg;
  assign data_o[199] = data_o_199_sv2v_reg;
  assign data_o[198] = data_o_198_sv2v_reg;
  assign data_o[197] = data_o_197_sv2v_reg;
  assign data_o[196] = data_o_196_sv2v_reg;
  assign data_o[195] = data_o_195_sv2v_reg;
  assign data_o[194] = data_o_194_sv2v_reg;
  assign data_o[193] = data_o_193_sv2v_reg;
  assign data_o[192] = data_o_192_sv2v_reg;
  assign data_o[191] = data_o_191_sv2v_reg;
  assign data_o[190] = data_o_190_sv2v_reg;
  assign data_o[189] = data_o_189_sv2v_reg;
  assign data_o[188] = data_o_188_sv2v_reg;
  assign data_o[187] = data_o_187_sv2v_reg;
  assign data_o[186] = data_o_186_sv2v_reg;
  assign data_o[185] = data_o_185_sv2v_reg;
  assign data_o[184] = data_o_184_sv2v_reg;
  assign data_o[183] = data_o_183_sv2v_reg;
  assign data_o[182] = data_o_182_sv2v_reg;
  assign data_o[181] = data_o_181_sv2v_reg;
  assign data_o[180] = data_o_180_sv2v_reg;
  assign data_o[179] = data_o_179_sv2v_reg;
  assign data_o[178] = data_o_178_sv2v_reg;
  assign data_o[177] = data_o_177_sv2v_reg;
  assign data_o[176] = data_o_176_sv2v_reg;
  assign data_o[175] = data_o_175_sv2v_reg;
  assign data_o[174] = data_o_174_sv2v_reg;
  assign data_o[173] = data_o_173_sv2v_reg;
  assign data_o[172] = data_o_172_sv2v_reg;
  assign data_o[171] = data_o_171_sv2v_reg;
  assign data_o[170] = data_o_170_sv2v_reg;
  assign data_o[169] = data_o_169_sv2v_reg;
  assign data_o[168] = data_o_168_sv2v_reg;
  assign data_o[167] = data_o_167_sv2v_reg;
  assign data_o[166] = data_o_166_sv2v_reg;
  assign data_o[165] = data_o_165_sv2v_reg;
  assign data_o[164] = data_o_164_sv2v_reg;
  assign data_o[163] = data_o_163_sv2v_reg;
  assign data_o[162] = data_o_162_sv2v_reg;
  assign data_o[161] = data_o_161_sv2v_reg;
  assign data_o[160] = data_o_160_sv2v_reg;
  assign data_o[159] = data_o_159_sv2v_reg;
  assign data_o[158] = data_o_158_sv2v_reg;
  assign data_o[157] = data_o_157_sv2v_reg;
  assign data_o[156] = data_o_156_sv2v_reg;
  assign data_o[155] = data_o_155_sv2v_reg;
  assign data_o[154] = data_o_154_sv2v_reg;
  assign data_o[153] = data_o_153_sv2v_reg;
  assign data_o[152] = data_o_152_sv2v_reg;
  assign data_o[151] = data_o_151_sv2v_reg;
  assign data_o[150] = data_o_150_sv2v_reg;
  assign data_o[149] = data_o_149_sv2v_reg;
  assign data_o[148] = data_o_148_sv2v_reg;
  assign data_o[147] = data_o_147_sv2v_reg;
  assign data_o[146] = data_o_146_sv2v_reg;
  assign data_o[145] = data_o_145_sv2v_reg;
  assign data_o[144] = data_o_144_sv2v_reg;
  assign data_o[143] = data_o_143_sv2v_reg;
  assign data_o[142] = data_o_142_sv2v_reg;
  assign data_o[141] = data_o_141_sv2v_reg;
  assign data_o[140] = data_o_140_sv2v_reg;
  assign data_o[139] = data_o_139_sv2v_reg;
  assign data_o[138] = data_o_138_sv2v_reg;
  assign data_o[137] = data_o_137_sv2v_reg;
  assign data_o[136] = data_o_136_sv2v_reg;
  assign data_o[135] = data_o_135_sv2v_reg;
  assign data_o[134] = data_o_134_sv2v_reg;
  assign data_o[133] = data_o_133_sv2v_reg;
  assign data_o[132] = data_o_132_sv2v_reg;
  assign data_o[131] = data_o_131_sv2v_reg;
  assign data_o[130] = data_o_130_sv2v_reg;
  assign data_o[129] = data_o_129_sv2v_reg;
  assign data_o[128] = data_o_128_sv2v_reg;
  assign data_o[127] = data_o_127_sv2v_reg;
  assign data_o[126] = data_o_126_sv2v_reg;
  assign data_o[125] = data_o_125_sv2v_reg;
  assign data_o[124] = data_o_124_sv2v_reg;
  assign data_o[123] = data_o_123_sv2v_reg;
  assign data_o[122] = data_o_122_sv2v_reg;
  assign data_o[121] = data_o_121_sv2v_reg;
  assign data_o[120] = data_o_120_sv2v_reg;
  assign data_o[119] = data_o_119_sv2v_reg;
  assign data_o[118] = data_o_118_sv2v_reg;
  assign data_o[117] = data_o_117_sv2v_reg;
  assign data_o[116] = data_o_116_sv2v_reg;
  assign data_o[115] = data_o_115_sv2v_reg;
  assign data_o[114] = data_o_114_sv2v_reg;
  assign data_o[113] = data_o_113_sv2v_reg;
  assign data_o[112] = data_o_112_sv2v_reg;
  assign data_o[111] = data_o_111_sv2v_reg;
  assign data_o[110] = data_o_110_sv2v_reg;
  assign data_o[109] = data_o_109_sv2v_reg;
  assign data_o[108] = data_o_108_sv2v_reg;
  assign data_o[107] = data_o_107_sv2v_reg;
  assign data_o[106] = data_o_106_sv2v_reg;
  assign data_o[105] = data_o_105_sv2v_reg;
  assign data_o[104] = data_o_104_sv2v_reg;
  assign data_o[103] = data_o_103_sv2v_reg;
  assign data_o[102] = data_o_102_sv2v_reg;
  assign data_o[101] = data_o_101_sv2v_reg;
  assign data_o[100] = data_o_100_sv2v_reg;
  assign data_o[99] = data_o_99_sv2v_reg;
  assign data_o[98] = data_o_98_sv2v_reg;
  assign data_o[97] = data_o_97_sv2v_reg;
  assign data_o[96] = data_o_96_sv2v_reg;
  assign data_o[95] = data_o_95_sv2v_reg;
  assign data_o[94] = data_o_94_sv2v_reg;
  assign data_o[93] = data_o_93_sv2v_reg;
  assign data_o[92] = data_o_92_sv2v_reg;
  assign data_o[91] = data_o_91_sv2v_reg;
  assign data_o[90] = data_o_90_sv2v_reg;
  assign data_o[89] = data_o_89_sv2v_reg;
  assign data_o[88] = data_o_88_sv2v_reg;
  assign data_o[87] = data_o_87_sv2v_reg;
  assign data_o[86] = data_o_86_sv2v_reg;
  assign data_o[85] = data_o_85_sv2v_reg;
  assign data_o[84] = data_o_84_sv2v_reg;
  assign data_o[83] = data_o_83_sv2v_reg;
  assign data_o[82] = data_o_82_sv2v_reg;
  assign data_o[81] = data_o_81_sv2v_reg;
  assign data_o[80] = data_o_80_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign { N7, N6, N5, N4, N3, N2 } = (N0)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                      (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_540_sv2v_reg <= 1'b0;
      data_o_539_sv2v_reg <= 1'b0;
      data_o_538_sv2v_reg <= 1'b0;
      data_o_537_sv2v_reg <= 1'b0;
      data_o_536_sv2v_reg <= 1'b0;
      data_o_535_sv2v_reg <= 1'b0;
      data_o_534_sv2v_reg <= 1'b0;
      data_o_533_sv2v_reg <= 1'b0;
      data_o_532_sv2v_reg <= 1'b0;
      data_o_531_sv2v_reg <= 1'b0;
      data_o_530_sv2v_reg <= 1'b0;
      data_o_529_sv2v_reg <= 1'b0;
      data_o_528_sv2v_reg <= 1'b0;
      data_o_527_sv2v_reg <= 1'b0;
      data_o_526_sv2v_reg <= 1'b0;
      data_o_525_sv2v_reg <= 1'b0;
      data_o_524_sv2v_reg <= 1'b0;
      data_o_523_sv2v_reg <= 1'b0;
      data_o_522_sv2v_reg <= 1'b0;
      data_o_521_sv2v_reg <= 1'b0;
      data_o_520_sv2v_reg <= 1'b0;
      data_o_519_sv2v_reg <= 1'b0;
      data_o_518_sv2v_reg <= 1'b0;
      data_o_517_sv2v_reg <= 1'b0;
      data_o_516_sv2v_reg <= 1'b0;
      data_o_515_sv2v_reg <= 1'b0;
      data_o_514_sv2v_reg <= 1'b0;
      data_o_513_sv2v_reg <= 1'b0;
      data_o_512_sv2v_reg <= 1'b0;
      data_o_511_sv2v_reg <= 1'b0;
      data_o_510_sv2v_reg <= 1'b0;
      data_o_509_sv2v_reg <= 1'b0;
      data_o_508_sv2v_reg <= 1'b0;
      data_o_507_sv2v_reg <= 1'b0;
      data_o_506_sv2v_reg <= 1'b0;
      data_o_505_sv2v_reg <= 1'b0;
      data_o_504_sv2v_reg <= 1'b0;
      data_o_503_sv2v_reg <= 1'b0;
      data_o_502_sv2v_reg <= 1'b0;
      data_o_501_sv2v_reg <= 1'b0;
      data_o_500_sv2v_reg <= 1'b0;
      data_o_499_sv2v_reg <= 1'b0;
      data_o_498_sv2v_reg <= 1'b0;
      data_o_497_sv2v_reg <= 1'b0;
      data_o_496_sv2v_reg <= 1'b0;
      data_o_495_sv2v_reg <= 1'b0;
      data_o_494_sv2v_reg <= 1'b0;
      data_o_493_sv2v_reg <= 1'b0;
      data_o_492_sv2v_reg <= 1'b0;
      data_o_491_sv2v_reg <= 1'b0;
      data_o_490_sv2v_reg <= 1'b0;
      data_o_489_sv2v_reg <= 1'b0;
      data_o_488_sv2v_reg <= 1'b0;
      data_o_487_sv2v_reg <= 1'b0;
      data_o_486_sv2v_reg <= 1'b0;
      data_o_485_sv2v_reg <= 1'b0;
      data_o_484_sv2v_reg <= 1'b0;
      data_o_483_sv2v_reg <= 1'b0;
      data_o_482_sv2v_reg <= 1'b0;
      data_o_481_sv2v_reg <= 1'b0;
      data_o_480_sv2v_reg <= 1'b0;
      data_o_479_sv2v_reg <= 1'b0;
      data_o_478_sv2v_reg <= 1'b0;
      data_o_477_sv2v_reg <= 1'b0;
      data_o_476_sv2v_reg <= 1'b0;
      data_o_475_sv2v_reg <= 1'b0;
      data_o_474_sv2v_reg <= 1'b0;
      data_o_473_sv2v_reg <= 1'b0;
      data_o_472_sv2v_reg <= 1'b0;
      data_o_471_sv2v_reg <= 1'b0;
      data_o_470_sv2v_reg <= 1'b0;
      data_o_469_sv2v_reg <= 1'b0;
      data_o_468_sv2v_reg <= 1'b0;
      data_o_467_sv2v_reg <= 1'b0;
      data_o_466_sv2v_reg <= 1'b0;
      data_o_465_sv2v_reg <= 1'b0;
      data_o_464_sv2v_reg <= 1'b0;
      data_o_463_sv2v_reg <= 1'b0;
      data_o_462_sv2v_reg <= 1'b0;
      data_o_461_sv2v_reg <= 1'b0;
      data_o_460_sv2v_reg <= 1'b0;
      data_o_459_sv2v_reg <= 1'b0;
      data_o_458_sv2v_reg <= 1'b0;
      data_o_457_sv2v_reg <= 1'b0;
      data_o_456_sv2v_reg <= 1'b0;
      data_o_455_sv2v_reg <= 1'b0;
      data_o_454_sv2v_reg <= 1'b0;
      data_o_453_sv2v_reg <= 1'b0;
      data_o_452_sv2v_reg <= 1'b0;
      data_o_451_sv2v_reg <= 1'b0;
      data_o_450_sv2v_reg <= 1'b0;
      data_o_449_sv2v_reg <= 1'b0;
      data_o_448_sv2v_reg <= 1'b0;
      data_o_447_sv2v_reg <= 1'b0;
      data_o_446_sv2v_reg <= 1'b0;
      data_o_445_sv2v_reg <= 1'b0;
      data_o_444_sv2v_reg <= 1'b0;
      data_o_443_sv2v_reg <= 1'b0;
      data_o_442_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_540_sv2v_reg <= data_i[540];
      data_o_539_sv2v_reg <= data_i[539];
      data_o_538_sv2v_reg <= data_i[538];
      data_o_537_sv2v_reg <= data_i[537];
      data_o_536_sv2v_reg <= data_i[536];
      data_o_535_sv2v_reg <= data_i[535];
      data_o_534_sv2v_reg <= data_i[534];
      data_o_533_sv2v_reg <= data_i[533];
      data_o_532_sv2v_reg <= data_i[532];
      data_o_531_sv2v_reg <= data_i[531];
      data_o_530_sv2v_reg <= data_i[530];
      data_o_529_sv2v_reg <= data_i[529];
      data_o_528_sv2v_reg <= data_i[528];
      data_o_527_sv2v_reg <= data_i[527];
      data_o_526_sv2v_reg <= data_i[526];
      data_o_525_sv2v_reg <= data_i[525];
      data_o_524_sv2v_reg <= data_i[524];
      data_o_523_sv2v_reg <= data_i[523];
      data_o_522_sv2v_reg <= data_i[522];
      data_o_521_sv2v_reg <= data_i[521];
      data_o_520_sv2v_reg <= data_i[520];
      data_o_519_sv2v_reg <= data_i[519];
      data_o_518_sv2v_reg <= data_i[518];
      data_o_517_sv2v_reg <= data_i[517];
      data_o_516_sv2v_reg <= data_i[516];
      data_o_515_sv2v_reg <= data_i[515];
      data_o_514_sv2v_reg <= data_i[514];
      data_o_513_sv2v_reg <= data_i[513];
      data_o_512_sv2v_reg <= data_i[512];
      data_o_511_sv2v_reg <= data_i[511];
      data_o_510_sv2v_reg <= data_i[510];
      data_o_509_sv2v_reg <= data_i[509];
      data_o_508_sv2v_reg <= data_i[508];
      data_o_507_sv2v_reg <= data_i[507];
      data_o_506_sv2v_reg <= data_i[506];
      data_o_505_sv2v_reg <= data_i[505];
      data_o_504_sv2v_reg <= data_i[504];
      data_o_503_sv2v_reg <= data_i[503];
      data_o_502_sv2v_reg <= data_i[502];
      data_o_501_sv2v_reg <= data_i[501];
      data_o_500_sv2v_reg <= data_i[500];
      data_o_499_sv2v_reg <= data_i[499];
      data_o_498_sv2v_reg <= data_i[498];
      data_o_497_sv2v_reg <= data_i[497];
      data_o_496_sv2v_reg <= data_i[496];
      data_o_495_sv2v_reg <= data_i[495];
      data_o_494_sv2v_reg <= data_i[494];
      data_o_493_sv2v_reg <= data_i[493];
      data_o_492_sv2v_reg <= data_i[492];
      data_o_491_sv2v_reg <= data_i[491];
      data_o_490_sv2v_reg <= data_i[490];
      data_o_489_sv2v_reg <= data_i[489];
      data_o_488_sv2v_reg <= data_i[488];
      data_o_487_sv2v_reg <= data_i[487];
      data_o_486_sv2v_reg <= data_i[486];
      data_o_485_sv2v_reg <= data_i[485];
      data_o_484_sv2v_reg <= data_i[484];
      data_o_483_sv2v_reg <= data_i[483];
      data_o_482_sv2v_reg <= data_i[482];
      data_o_481_sv2v_reg <= data_i[481];
      data_o_480_sv2v_reg <= data_i[480];
      data_o_479_sv2v_reg <= data_i[479];
      data_o_478_sv2v_reg <= data_i[478];
      data_o_477_sv2v_reg <= data_i[477];
      data_o_476_sv2v_reg <= data_i[476];
      data_o_475_sv2v_reg <= data_i[475];
      data_o_474_sv2v_reg <= data_i[474];
      data_o_473_sv2v_reg <= data_i[473];
      data_o_472_sv2v_reg <= data_i[472];
      data_o_471_sv2v_reg <= data_i[471];
      data_o_470_sv2v_reg <= data_i[470];
      data_o_469_sv2v_reg <= data_i[469];
      data_o_468_sv2v_reg <= data_i[468];
      data_o_467_sv2v_reg <= data_i[467];
      data_o_466_sv2v_reg <= data_i[466];
      data_o_465_sv2v_reg <= data_i[465];
      data_o_464_sv2v_reg <= data_i[464];
      data_o_463_sv2v_reg <= data_i[463];
      data_o_462_sv2v_reg <= data_i[462];
      data_o_461_sv2v_reg <= data_i[461];
      data_o_460_sv2v_reg <= data_i[460];
      data_o_459_sv2v_reg <= data_i[459];
      data_o_458_sv2v_reg <= data_i[458];
      data_o_457_sv2v_reg <= data_i[457];
      data_o_456_sv2v_reg <= data_i[456];
      data_o_455_sv2v_reg <= data_i[455];
      data_o_454_sv2v_reg <= data_i[454];
      data_o_453_sv2v_reg <= data_i[453];
      data_o_452_sv2v_reg <= data_i[452];
      data_o_451_sv2v_reg <= data_i[451];
      data_o_450_sv2v_reg <= data_i[450];
      data_o_449_sv2v_reg <= data_i[449];
      data_o_448_sv2v_reg <= data_i[448];
      data_o_447_sv2v_reg <= data_i[447];
      data_o_446_sv2v_reg <= data_i[446];
      data_o_445_sv2v_reg <= data_i[445];
      data_o_444_sv2v_reg <= data_i[444];
      data_o_443_sv2v_reg <= data_i[443];
      data_o_442_sv2v_reg <= data_i[442];
      data_o_0_sv2v_reg <= data_i[0];
    end 
    if(reset_i) begin
      data_o_441_sv2v_reg <= 1'b0;
      data_o_440_sv2v_reg <= 1'b0;
      data_o_439_sv2v_reg <= 1'b0;
      data_o_438_sv2v_reg <= 1'b0;
      data_o_437_sv2v_reg <= 1'b0;
      data_o_436_sv2v_reg <= 1'b0;
      data_o_435_sv2v_reg <= 1'b0;
      data_o_434_sv2v_reg <= 1'b0;
      data_o_433_sv2v_reg <= 1'b0;
      data_o_432_sv2v_reg <= 1'b0;
      data_o_431_sv2v_reg <= 1'b0;
      data_o_430_sv2v_reg <= 1'b0;
      data_o_429_sv2v_reg <= 1'b0;
      data_o_428_sv2v_reg <= 1'b0;
      data_o_427_sv2v_reg <= 1'b0;
      data_o_426_sv2v_reg <= 1'b0;
      data_o_425_sv2v_reg <= 1'b0;
      data_o_424_sv2v_reg <= 1'b0;
      data_o_423_sv2v_reg <= 1'b0;
      data_o_422_sv2v_reg <= 1'b0;
      data_o_421_sv2v_reg <= 1'b0;
      data_o_420_sv2v_reg <= 1'b0;
      data_o_419_sv2v_reg <= 1'b0;
      data_o_418_sv2v_reg <= 1'b0;
      data_o_417_sv2v_reg <= 1'b0;
      data_o_416_sv2v_reg <= 1'b0;
      data_o_415_sv2v_reg <= 1'b0;
      data_o_414_sv2v_reg <= 1'b0;
      data_o_413_sv2v_reg <= 1'b0;
      data_o_412_sv2v_reg <= 1'b0;
      data_o_411_sv2v_reg <= 1'b0;
      data_o_410_sv2v_reg <= 1'b0;
      data_o_409_sv2v_reg <= 1'b0;
      data_o_408_sv2v_reg <= 1'b0;
      data_o_407_sv2v_reg <= 1'b0;
      data_o_406_sv2v_reg <= 1'b0;
      data_o_405_sv2v_reg <= 1'b0;
      data_o_404_sv2v_reg <= 1'b0;
      data_o_403_sv2v_reg <= 1'b0;
      data_o_402_sv2v_reg <= 1'b0;
      data_o_401_sv2v_reg <= 1'b0;
      data_o_400_sv2v_reg <= 1'b0;
      data_o_399_sv2v_reg <= 1'b0;
      data_o_398_sv2v_reg <= 1'b0;
      data_o_397_sv2v_reg <= 1'b0;
      data_o_396_sv2v_reg <= 1'b0;
      data_o_395_sv2v_reg <= 1'b0;
      data_o_394_sv2v_reg <= 1'b0;
      data_o_393_sv2v_reg <= 1'b0;
      data_o_392_sv2v_reg <= 1'b0;
      data_o_391_sv2v_reg <= 1'b0;
      data_o_390_sv2v_reg <= 1'b0;
      data_o_389_sv2v_reg <= 1'b0;
      data_o_388_sv2v_reg <= 1'b0;
      data_o_387_sv2v_reg <= 1'b0;
      data_o_386_sv2v_reg <= 1'b0;
      data_o_385_sv2v_reg <= 1'b0;
      data_o_384_sv2v_reg <= 1'b0;
      data_o_383_sv2v_reg <= 1'b0;
      data_o_382_sv2v_reg <= 1'b0;
      data_o_381_sv2v_reg <= 1'b0;
      data_o_380_sv2v_reg <= 1'b0;
      data_o_379_sv2v_reg <= 1'b0;
      data_o_378_sv2v_reg <= 1'b0;
      data_o_377_sv2v_reg <= 1'b0;
      data_o_376_sv2v_reg <= 1'b0;
      data_o_375_sv2v_reg <= 1'b0;
      data_o_374_sv2v_reg <= 1'b0;
      data_o_373_sv2v_reg <= 1'b0;
      data_o_372_sv2v_reg <= 1'b0;
      data_o_371_sv2v_reg <= 1'b0;
      data_o_370_sv2v_reg <= 1'b0;
      data_o_369_sv2v_reg <= 1'b0;
      data_o_368_sv2v_reg <= 1'b0;
      data_o_367_sv2v_reg <= 1'b0;
      data_o_366_sv2v_reg <= 1'b0;
      data_o_365_sv2v_reg <= 1'b0;
      data_o_364_sv2v_reg <= 1'b0;
      data_o_363_sv2v_reg <= 1'b0;
      data_o_362_sv2v_reg <= 1'b0;
      data_o_361_sv2v_reg <= 1'b0;
      data_o_360_sv2v_reg <= 1'b0;
      data_o_359_sv2v_reg <= 1'b0;
      data_o_358_sv2v_reg <= 1'b0;
      data_o_357_sv2v_reg <= 1'b0;
      data_o_356_sv2v_reg <= 1'b0;
      data_o_355_sv2v_reg <= 1'b0;
      data_o_354_sv2v_reg <= 1'b0;
      data_o_353_sv2v_reg <= 1'b0;
      data_o_352_sv2v_reg <= 1'b0;
      data_o_351_sv2v_reg <= 1'b0;
      data_o_350_sv2v_reg <= 1'b0;
      data_o_349_sv2v_reg <= 1'b0;
      data_o_348_sv2v_reg <= 1'b0;
      data_o_347_sv2v_reg <= 1'b0;
      data_o_346_sv2v_reg <= 1'b0;
      data_o_345_sv2v_reg <= 1'b0;
      data_o_344_sv2v_reg <= 1'b0;
      data_o_343_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
    end else if(N3) begin
      data_o_441_sv2v_reg <= data_i[441];
      data_o_440_sv2v_reg <= data_i[440];
      data_o_439_sv2v_reg <= data_i[439];
      data_o_438_sv2v_reg <= data_i[438];
      data_o_437_sv2v_reg <= data_i[437];
      data_o_436_sv2v_reg <= data_i[436];
      data_o_435_sv2v_reg <= data_i[435];
      data_o_434_sv2v_reg <= data_i[434];
      data_o_433_sv2v_reg <= data_i[433];
      data_o_432_sv2v_reg <= data_i[432];
      data_o_431_sv2v_reg <= data_i[431];
      data_o_430_sv2v_reg <= data_i[430];
      data_o_429_sv2v_reg <= data_i[429];
      data_o_428_sv2v_reg <= data_i[428];
      data_o_427_sv2v_reg <= data_i[427];
      data_o_426_sv2v_reg <= data_i[426];
      data_o_425_sv2v_reg <= data_i[425];
      data_o_424_sv2v_reg <= data_i[424];
      data_o_423_sv2v_reg <= data_i[423];
      data_o_422_sv2v_reg <= data_i[422];
      data_o_421_sv2v_reg <= data_i[421];
      data_o_420_sv2v_reg <= data_i[420];
      data_o_419_sv2v_reg <= data_i[419];
      data_o_418_sv2v_reg <= data_i[418];
      data_o_417_sv2v_reg <= data_i[417];
      data_o_416_sv2v_reg <= data_i[416];
      data_o_415_sv2v_reg <= data_i[415];
      data_o_414_sv2v_reg <= data_i[414];
      data_o_413_sv2v_reg <= data_i[413];
      data_o_412_sv2v_reg <= data_i[412];
      data_o_411_sv2v_reg <= data_i[411];
      data_o_410_sv2v_reg <= data_i[410];
      data_o_409_sv2v_reg <= data_i[409];
      data_o_408_sv2v_reg <= data_i[408];
      data_o_407_sv2v_reg <= data_i[407];
      data_o_406_sv2v_reg <= data_i[406];
      data_o_405_sv2v_reg <= data_i[405];
      data_o_404_sv2v_reg <= data_i[404];
      data_o_403_sv2v_reg <= data_i[403];
      data_o_402_sv2v_reg <= data_i[402];
      data_o_401_sv2v_reg <= data_i[401];
      data_o_400_sv2v_reg <= data_i[400];
      data_o_399_sv2v_reg <= data_i[399];
      data_o_398_sv2v_reg <= data_i[398];
      data_o_397_sv2v_reg <= data_i[397];
      data_o_396_sv2v_reg <= data_i[396];
      data_o_395_sv2v_reg <= data_i[395];
      data_o_394_sv2v_reg <= data_i[394];
      data_o_393_sv2v_reg <= data_i[393];
      data_o_392_sv2v_reg <= data_i[392];
      data_o_391_sv2v_reg <= data_i[391];
      data_o_390_sv2v_reg <= data_i[390];
      data_o_389_sv2v_reg <= data_i[389];
      data_o_388_sv2v_reg <= data_i[388];
      data_o_387_sv2v_reg <= data_i[387];
      data_o_386_sv2v_reg <= data_i[386];
      data_o_385_sv2v_reg <= data_i[385];
      data_o_384_sv2v_reg <= data_i[384];
      data_o_383_sv2v_reg <= data_i[383];
      data_o_382_sv2v_reg <= data_i[382];
      data_o_381_sv2v_reg <= data_i[381];
      data_o_380_sv2v_reg <= data_i[380];
      data_o_379_sv2v_reg <= data_i[379];
      data_o_378_sv2v_reg <= data_i[378];
      data_o_377_sv2v_reg <= data_i[377];
      data_o_376_sv2v_reg <= data_i[376];
      data_o_375_sv2v_reg <= data_i[375];
      data_o_374_sv2v_reg <= data_i[374];
      data_o_373_sv2v_reg <= data_i[373];
      data_o_372_sv2v_reg <= data_i[372];
      data_o_371_sv2v_reg <= data_i[371];
      data_o_370_sv2v_reg <= data_i[370];
      data_o_369_sv2v_reg <= data_i[369];
      data_o_368_sv2v_reg <= data_i[368];
      data_o_367_sv2v_reg <= data_i[367];
      data_o_366_sv2v_reg <= data_i[366];
      data_o_365_sv2v_reg <= data_i[365];
      data_o_364_sv2v_reg <= data_i[364];
      data_o_363_sv2v_reg <= data_i[363];
      data_o_362_sv2v_reg <= data_i[362];
      data_o_361_sv2v_reg <= data_i[361];
      data_o_360_sv2v_reg <= data_i[360];
      data_o_359_sv2v_reg <= data_i[359];
      data_o_358_sv2v_reg <= data_i[358];
      data_o_357_sv2v_reg <= data_i[357];
      data_o_356_sv2v_reg <= data_i[356];
      data_o_355_sv2v_reg <= data_i[355];
      data_o_354_sv2v_reg <= data_i[354];
      data_o_353_sv2v_reg <= data_i[353];
      data_o_352_sv2v_reg <= data_i[352];
      data_o_351_sv2v_reg <= data_i[351];
      data_o_350_sv2v_reg <= data_i[350];
      data_o_349_sv2v_reg <= data_i[349];
      data_o_348_sv2v_reg <= data_i[348];
      data_o_347_sv2v_reg <= data_i[347];
      data_o_346_sv2v_reg <= data_i[346];
      data_o_345_sv2v_reg <= data_i[345];
      data_o_344_sv2v_reg <= data_i[344];
      data_o_343_sv2v_reg <= data_i[343];
      data_o_1_sv2v_reg <= data_i[1];
    end 
    if(reset_i) begin
      data_o_342_sv2v_reg <= 1'b0;
      data_o_341_sv2v_reg <= 1'b0;
      data_o_340_sv2v_reg <= 1'b0;
      data_o_339_sv2v_reg <= 1'b0;
      data_o_338_sv2v_reg <= 1'b0;
      data_o_337_sv2v_reg <= 1'b0;
      data_o_336_sv2v_reg <= 1'b0;
      data_o_335_sv2v_reg <= 1'b0;
      data_o_334_sv2v_reg <= 1'b0;
      data_o_333_sv2v_reg <= 1'b0;
      data_o_332_sv2v_reg <= 1'b0;
      data_o_331_sv2v_reg <= 1'b0;
      data_o_330_sv2v_reg <= 1'b0;
      data_o_329_sv2v_reg <= 1'b0;
      data_o_328_sv2v_reg <= 1'b0;
      data_o_327_sv2v_reg <= 1'b0;
      data_o_326_sv2v_reg <= 1'b0;
      data_o_325_sv2v_reg <= 1'b0;
      data_o_324_sv2v_reg <= 1'b0;
      data_o_323_sv2v_reg <= 1'b0;
      data_o_322_sv2v_reg <= 1'b0;
      data_o_321_sv2v_reg <= 1'b0;
      data_o_320_sv2v_reg <= 1'b0;
      data_o_319_sv2v_reg <= 1'b0;
      data_o_318_sv2v_reg <= 1'b0;
      data_o_317_sv2v_reg <= 1'b0;
      data_o_316_sv2v_reg <= 1'b0;
      data_o_315_sv2v_reg <= 1'b0;
      data_o_314_sv2v_reg <= 1'b0;
      data_o_313_sv2v_reg <= 1'b0;
      data_o_312_sv2v_reg <= 1'b0;
      data_o_311_sv2v_reg <= 1'b0;
      data_o_310_sv2v_reg <= 1'b0;
      data_o_309_sv2v_reg <= 1'b0;
      data_o_308_sv2v_reg <= 1'b0;
      data_o_307_sv2v_reg <= 1'b0;
      data_o_306_sv2v_reg <= 1'b0;
      data_o_305_sv2v_reg <= 1'b0;
      data_o_304_sv2v_reg <= 1'b0;
      data_o_303_sv2v_reg <= 1'b0;
      data_o_302_sv2v_reg <= 1'b0;
      data_o_301_sv2v_reg <= 1'b0;
      data_o_300_sv2v_reg <= 1'b0;
      data_o_299_sv2v_reg <= 1'b0;
      data_o_298_sv2v_reg <= 1'b0;
      data_o_297_sv2v_reg <= 1'b0;
      data_o_296_sv2v_reg <= 1'b0;
      data_o_295_sv2v_reg <= 1'b0;
      data_o_294_sv2v_reg <= 1'b0;
      data_o_293_sv2v_reg <= 1'b0;
      data_o_292_sv2v_reg <= 1'b0;
      data_o_291_sv2v_reg <= 1'b0;
      data_o_290_sv2v_reg <= 1'b0;
      data_o_289_sv2v_reg <= 1'b0;
      data_o_288_sv2v_reg <= 1'b0;
      data_o_287_sv2v_reg <= 1'b0;
      data_o_286_sv2v_reg <= 1'b0;
      data_o_285_sv2v_reg <= 1'b0;
      data_o_284_sv2v_reg <= 1'b0;
      data_o_283_sv2v_reg <= 1'b0;
      data_o_282_sv2v_reg <= 1'b0;
      data_o_281_sv2v_reg <= 1'b0;
      data_o_280_sv2v_reg <= 1'b0;
      data_o_279_sv2v_reg <= 1'b0;
      data_o_278_sv2v_reg <= 1'b0;
      data_o_277_sv2v_reg <= 1'b0;
      data_o_276_sv2v_reg <= 1'b0;
      data_o_275_sv2v_reg <= 1'b0;
      data_o_274_sv2v_reg <= 1'b0;
      data_o_273_sv2v_reg <= 1'b0;
      data_o_272_sv2v_reg <= 1'b0;
      data_o_271_sv2v_reg <= 1'b0;
      data_o_270_sv2v_reg <= 1'b0;
      data_o_269_sv2v_reg <= 1'b0;
      data_o_268_sv2v_reg <= 1'b0;
      data_o_267_sv2v_reg <= 1'b0;
      data_o_266_sv2v_reg <= 1'b0;
      data_o_265_sv2v_reg <= 1'b0;
      data_o_264_sv2v_reg <= 1'b0;
      data_o_263_sv2v_reg <= 1'b0;
      data_o_262_sv2v_reg <= 1'b0;
      data_o_261_sv2v_reg <= 1'b0;
      data_o_260_sv2v_reg <= 1'b0;
      data_o_259_sv2v_reg <= 1'b0;
      data_o_258_sv2v_reg <= 1'b0;
      data_o_257_sv2v_reg <= 1'b0;
      data_o_256_sv2v_reg <= 1'b0;
      data_o_255_sv2v_reg <= 1'b0;
      data_o_254_sv2v_reg <= 1'b0;
      data_o_253_sv2v_reg <= 1'b0;
      data_o_252_sv2v_reg <= 1'b0;
      data_o_251_sv2v_reg <= 1'b0;
      data_o_250_sv2v_reg <= 1'b0;
      data_o_249_sv2v_reg <= 1'b0;
      data_o_248_sv2v_reg <= 1'b0;
      data_o_247_sv2v_reg <= 1'b0;
      data_o_246_sv2v_reg <= 1'b0;
      data_o_245_sv2v_reg <= 1'b0;
      data_o_244_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
    end else if(N4) begin
      data_o_342_sv2v_reg <= data_i[342];
      data_o_341_sv2v_reg <= data_i[341];
      data_o_340_sv2v_reg <= data_i[340];
      data_o_339_sv2v_reg <= data_i[339];
      data_o_338_sv2v_reg <= data_i[338];
      data_o_337_sv2v_reg <= data_i[337];
      data_o_336_sv2v_reg <= data_i[336];
      data_o_335_sv2v_reg <= data_i[335];
      data_o_334_sv2v_reg <= data_i[334];
      data_o_333_sv2v_reg <= data_i[333];
      data_o_332_sv2v_reg <= data_i[332];
      data_o_331_sv2v_reg <= data_i[331];
      data_o_330_sv2v_reg <= data_i[330];
      data_o_329_sv2v_reg <= data_i[329];
      data_o_328_sv2v_reg <= data_i[328];
      data_o_327_sv2v_reg <= data_i[327];
      data_o_326_sv2v_reg <= data_i[326];
      data_o_325_sv2v_reg <= data_i[325];
      data_o_324_sv2v_reg <= data_i[324];
      data_o_323_sv2v_reg <= data_i[323];
      data_o_322_sv2v_reg <= data_i[322];
      data_o_321_sv2v_reg <= data_i[321];
      data_o_320_sv2v_reg <= data_i[320];
      data_o_319_sv2v_reg <= data_i[319];
      data_o_318_sv2v_reg <= data_i[318];
      data_o_317_sv2v_reg <= data_i[317];
      data_o_316_sv2v_reg <= data_i[316];
      data_o_315_sv2v_reg <= data_i[315];
      data_o_314_sv2v_reg <= data_i[314];
      data_o_313_sv2v_reg <= data_i[313];
      data_o_312_sv2v_reg <= data_i[312];
      data_o_311_sv2v_reg <= data_i[311];
      data_o_310_sv2v_reg <= data_i[310];
      data_o_309_sv2v_reg <= data_i[309];
      data_o_308_sv2v_reg <= data_i[308];
      data_o_307_sv2v_reg <= data_i[307];
      data_o_306_sv2v_reg <= data_i[306];
      data_o_305_sv2v_reg <= data_i[305];
      data_o_304_sv2v_reg <= data_i[304];
      data_o_303_sv2v_reg <= data_i[303];
      data_o_302_sv2v_reg <= data_i[302];
      data_o_301_sv2v_reg <= data_i[301];
      data_o_300_sv2v_reg <= data_i[300];
      data_o_299_sv2v_reg <= data_i[299];
      data_o_298_sv2v_reg <= data_i[298];
      data_o_297_sv2v_reg <= data_i[297];
      data_o_296_sv2v_reg <= data_i[296];
      data_o_295_sv2v_reg <= data_i[295];
      data_o_294_sv2v_reg <= data_i[294];
      data_o_293_sv2v_reg <= data_i[293];
      data_o_292_sv2v_reg <= data_i[292];
      data_o_291_sv2v_reg <= data_i[291];
      data_o_290_sv2v_reg <= data_i[290];
      data_o_289_sv2v_reg <= data_i[289];
      data_o_288_sv2v_reg <= data_i[288];
      data_o_287_sv2v_reg <= data_i[287];
      data_o_286_sv2v_reg <= data_i[286];
      data_o_285_sv2v_reg <= data_i[285];
      data_o_284_sv2v_reg <= data_i[284];
      data_o_283_sv2v_reg <= data_i[283];
      data_o_282_sv2v_reg <= data_i[282];
      data_o_281_sv2v_reg <= data_i[281];
      data_o_280_sv2v_reg <= data_i[280];
      data_o_279_sv2v_reg <= data_i[279];
      data_o_278_sv2v_reg <= data_i[278];
      data_o_277_sv2v_reg <= data_i[277];
      data_o_276_sv2v_reg <= data_i[276];
      data_o_275_sv2v_reg <= data_i[275];
      data_o_274_sv2v_reg <= data_i[274];
      data_o_273_sv2v_reg <= data_i[273];
      data_o_272_sv2v_reg <= data_i[272];
      data_o_271_sv2v_reg <= data_i[271];
      data_o_270_sv2v_reg <= data_i[270];
      data_o_269_sv2v_reg <= data_i[269];
      data_o_268_sv2v_reg <= data_i[268];
      data_o_267_sv2v_reg <= data_i[267];
      data_o_266_sv2v_reg <= data_i[266];
      data_o_265_sv2v_reg <= data_i[265];
      data_o_264_sv2v_reg <= data_i[264];
      data_o_263_sv2v_reg <= data_i[263];
      data_o_262_sv2v_reg <= data_i[262];
      data_o_261_sv2v_reg <= data_i[261];
      data_o_260_sv2v_reg <= data_i[260];
      data_o_259_sv2v_reg <= data_i[259];
      data_o_258_sv2v_reg <= data_i[258];
      data_o_257_sv2v_reg <= data_i[257];
      data_o_256_sv2v_reg <= data_i[256];
      data_o_255_sv2v_reg <= data_i[255];
      data_o_254_sv2v_reg <= data_i[254];
      data_o_253_sv2v_reg <= data_i[253];
      data_o_252_sv2v_reg <= data_i[252];
      data_o_251_sv2v_reg <= data_i[251];
      data_o_250_sv2v_reg <= data_i[250];
      data_o_249_sv2v_reg <= data_i[249];
      data_o_248_sv2v_reg <= data_i[248];
      data_o_247_sv2v_reg <= data_i[247];
      data_o_246_sv2v_reg <= data_i[246];
      data_o_245_sv2v_reg <= data_i[245];
      data_o_244_sv2v_reg <= data_i[244];
      data_o_2_sv2v_reg <= data_i[2];
    end 
    if(reset_i) begin
      data_o_243_sv2v_reg <= 1'b0;
      data_o_242_sv2v_reg <= 1'b0;
      data_o_241_sv2v_reg <= 1'b0;
      data_o_240_sv2v_reg <= 1'b0;
      data_o_239_sv2v_reg <= 1'b0;
      data_o_238_sv2v_reg <= 1'b0;
      data_o_237_sv2v_reg <= 1'b0;
      data_o_236_sv2v_reg <= 1'b0;
      data_o_235_sv2v_reg <= 1'b0;
      data_o_234_sv2v_reg <= 1'b0;
      data_o_233_sv2v_reg <= 1'b0;
      data_o_232_sv2v_reg <= 1'b0;
      data_o_231_sv2v_reg <= 1'b0;
      data_o_230_sv2v_reg <= 1'b0;
      data_o_229_sv2v_reg <= 1'b0;
      data_o_228_sv2v_reg <= 1'b0;
      data_o_227_sv2v_reg <= 1'b0;
      data_o_226_sv2v_reg <= 1'b0;
      data_o_225_sv2v_reg <= 1'b0;
      data_o_224_sv2v_reg <= 1'b0;
      data_o_223_sv2v_reg <= 1'b0;
      data_o_222_sv2v_reg <= 1'b0;
      data_o_221_sv2v_reg <= 1'b0;
      data_o_220_sv2v_reg <= 1'b0;
      data_o_219_sv2v_reg <= 1'b0;
      data_o_218_sv2v_reg <= 1'b0;
      data_o_217_sv2v_reg <= 1'b0;
      data_o_216_sv2v_reg <= 1'b0;
      data_o_215_sv2v_reg <= 1'b0;
      data_o_214_sv2v_reg <= 1'b0;
      data_o_213_sv2v_reg <= 1'b0;
      data_o_212_sv2v_reg <= 1'b0;
      data_o_211_sv2v_reg <= 1'b0;
      data_o_210_sv2v_reg <= 1'b0;
      data_o_209_sv2v_reg <= 1'b0;
      data_o_208_sv2v_reg <= 1'b0;
      data_o_207_sv2v_reg <= 1'b0;
      data_o_206_sv2v_reg <= 1'b0;
      data_o_205_sv2v_reg <= 1'b0;
      data_o_204_sv2v_reg <= 1'b0;
      data_o_203_sv2v_reg <= 1'b0;
      data_o_202_sv2v_reg <= 1'b0;
      data_o_201_sv2v_reg <= 1'b0;
      data_o_200_sv2v_reg <= 1'b0;
      data_o_199_sv2v_reg <= 1'b0;
      data_o_198_sv2v_reg <= 1'b0;
      data_o_197_sv2v_reg <= 1'b0;
      data_o_196_sv2v_reg <= 1'b0;
      data_o_195_sv2v_reg <= 1'b0;
      data_o_194_sv2v_reg <= 1'b0;
      data_o_193_sv2v_reg <= 1'b0;
      data_o_192_sv2v_reg <= 1'b0;
      data_o_191_sv2v_reg <= 1'b0;
      data_o_190_sv2v_reg <= 1'b0;
      data_o_189_sv2v_reg <= 1'b0;
      data_o_188_sv2v_reg <= 1'b0;
      data_o_187_sv2v_reg <= 1'b0;
      data_o_186_sv2v_reg <= 1'b0;
      data_o_185_sv2v_reg <= 1'b0;
      data_o_184_sv2v_reg <= 1'b0;
      data_o_183_sv2v_reg <= 1'b0;
      data_o_182_sv2v_reg <= 1'b0;
      data_o_181_sv2v_reg <= 1'b0;
      data_o_180_sv2v_reg <= 1'b0;
      data_o_179_sv2v_reg <= 1'b0;
      data_o_178_sv2v_reg <= 1'b0;
      data_o_177_sv2v_reg <= 1'b0;
      data_o_176_sv2v_reg <= 1'b0;
      data_o_175_sv2v_reg <= 1'b0;
      data_o_174_sv2v_reg <= 1'b0;
      data_o_173_sv2v_reg <= 1'b0;
      data_o_172_sv2v_reg <= 1'b0;
      data_o_171_sv2v_reg <= 1'b0;
      data_o_170_sv2v_reg <= 1'b0;
      data_o_169_sv2v_reg <= 1'b0;
      data_o_168_sv2v_reg <= 1'b0;
      data_o_167_sv2v_reg <= 1'b0;
      data_o_166_sv2v_reg <= 1'b0;
      data_o_165_sv2v_reg <= 1'b0;
      data_o_164_sv2v_reg <= 1'b0;
      data_o_163_sv2v_reg <= 1'b0;
      data_o_162_sv2v_reg <= 1'b0;
      data_o_161_sv2v_reg <= 1'b0;
      data_o_160_sv2v_reg <= 1'b0;
      data_o_159_sv2v_reg <= 1'b0;
      data_o_158_sv2v_reg <= 1'b0;
      data_o_157_sv2v_reg <= 1'b0;
      data_o_156_sv2v_reg <= 1'b0;
      data_o_155_sv2v_reg <= 1'b0;
      data_o_154_sv2v_reg <= 1'b0;
      data_o_153_sv2v_reg <= 1'b0;
      data_o_152_sv2v_reg <= 1'b0;
      data_o_151_sv2v_reg <= 1'b0;
      data_o_150_sv2v_reg <= 1'b0;
      data_o_149_sv2v_reg <= 1'b0;
      data_o_148_sv2v_reg <= 1'b0;
      data_o_147_sv2v_reg <= 1'b0;
      data_o_146_sv2v_reg <= 1'b0;
      data_o_145_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
    end else if(N5) begin
      data_o_243_sv2v_reg <= data_i[243];
      data_o_242_sv2v_reg <= data_i[242];
      data_o_241_sv2v_reg <= data_i[241];
      data_o_240_sv2v_reg <= data_i[240];
      data_o_239_sv2v_reg <= data_i[239];
      data_o_238_sv2v_reg <= data_i[238];
      data_o_237_sv2v_reg <= data_i[237];
      data_o_236_sv2v_reg <= data_i[236];
      data_o_235_sv2v_reg <= data_i[235];
      data_o_234_sv2v_reg <= data_i[234];
      data_o_233_sv2v_reg <= data_i[233];
      data_o_232_sv2v_reg <= data_i[232];
      data_o_231_sv2v_reg <= data_i[231];
      data_o_230_sv2v_reg <= data_i[230];
      data_o_229_sv2v_reg <= data_i[229];
      data_o_228_sv2v_reg <= data_i[228];
      data_o_227_sv2v_reg <= data_i[227];
      data_o_226_sv2v_reg <= data_i[226];
      data_o_225_sv2v_reg <= data_i[225];
      data_o_224_sv2v_reg <= data_i[224];
      data_o_223_sv2v_reg <= data_i[223];
      data_o_222_sv2v_reg <= data_i[222];
      data_o_221_sv2v_reg <= data_i[221];
      data_o_220_sv2v_reg <= data_i[220];
      data_o_219_sv2v_reg <= data_i[219];
      data_o_218_sv2v_reg <= data_i[218];
      data_o_217_sv2v_reg <= data_i[217];
      data_o_216_sv2v_reg <= data_i[216];
      data_o_215_sv2v_reg <= data_i[215];
      data_o_214_sv2v_reg <= data_i[214];
      data_o_213_sv2v_reg <= data_i[213];
      data_o_212_sv2v_reg <= data_i[212];
      data_o_211_sv2v_reg <= data_i[211];
      data_o_210_sv2v_reg <= data_i[210];
      data_o_209_sv2v_reg <= data_i[209];
      data_o_208_sv2v_reg <= data_i[208];
      data_o_207_sv2v_reg <= data_i[207];
      data_o_206_sv2v_reg <= data_i[206];
      data_o_205_sv2v_reg <= data_i[205];
      data_o_204_sv2v_reg <= data_i[204];
      data_o_203_sv2v_reg <= data_i[203];
      data_o_202_sv2v_reg <= data_i[202];
      data_o_201_sv2v_reg <= data_i[201];
      data_o_200_sv2v_reg <= data_i[200];
      data_o_199_sv2v_reg <= data_i[199];
      data_o_198_sv2v_reg <= data_i[198];
      data_o_197_sv2v_reg <= data_i[197];
      data_o_196_sv2v_reg <= data_i[196];
      data_o_195_sv2v_reg <= data_i[195];
      data_o_194_sv2v_reg <= data_i[194];
      data_o_193_sv2v_reg <= data_i[193];
      data_o_192_sv2v_reg <= data_i[192];
      data_o_191_sv2v_reg <= data_i[191];
      data_o_190_sv2v_reg <= data_i[190];
      data_o_189_sv2v_reg <= data_i[189];
      data_o_188_sv2v_reg <= data_i[188];
      data_o_187_sv2v_reg <= data_i[187];
      data_o_186_sv2v_reg <= data_i[186];
      data_o_185_sv2v_reg <= data_i[185];
      data_o_184_sv2v_reg <= data_i[184];
      data_o_183_sv2v_reg <= data_i[183];
      data_o_182_sv2v_reg <= data_i[182];
      data_o_181_sv2v_reg <= data_i[181];
      data_o_180_sv2v_reg <= data_i[180];
      data_o_179_sv2v_reg <= data_i[179];
      data_o_178_sv2v_reg <= data_i[178];
      data_o_177_sv2v_reg <= data_i[177];
      data_o_176_sv2v_reg <= data_i[176];
      data_o_175_sv2v_reg <= data_i[175];
      data_o_174_sv2v_reg <= data_i[174];
      data_o_173_sv2v_reg <= data_i[173];
      data_o_172_sv2v_reg <= data_i[172];
      data_o_171_sv2v_reg <= data_i[171];
      data_o_170_sv2v_reg <= data_i[170];
      data_o_169_sv2v_reg <= data_i[169];
      data_o_168_sv2v_reg <= data_i[168];
      data_o_167_sv2v_reg <= data_i[167];
      data_o_166_sv2v_reg <= data_i[166];
      data_o_165_sv2v_reg <= data_i[165];
      data_o_164_sv2v_reg <= data_i[164];
      data_o_163_sv2v_reg <= data_i[163];
      data_o_162_sv2v_reg <= data_i[162];
      data_o_161_sv2v_reg <= data_i[161];
      data_o_160_sv2v_reg <= data_i[160];
      data_o_159_sv2v_reg <= data_i[159];
      data_o_158_sv2v_reg <= data_i[158];
      data_o_157_sv2v_reg <= data_i[157];
      data_o_156_sv2v_reg <= data_i[156];
      data_o_155_sv2v_reg <= data_i[155];
      data_o_154_sv2v_reg <= data_i[154];
      data_o_153_sv2v_reg <= data_i[153];
      data_o_152_sv2v_reg <= data_i[152];
      data_o_151_sv2v_reg <= data_i[151];
      data_o_150_sv2v_reg <= data_i[150];
      data_o_149_sv2v_reg <= data_i[149];
      data_o_148_sv2v_reg <= data_i[148];
      data_o_147_sv2v_reg <= data_i[147];
      data_o_146_sv2v_reg <= data_i[146];
      data_o_145_sv2v_reg <= data_i[145];
      data_o_3_sv2v_reg <= data_i[3];
    end 
    if(reset_i) begin
      data_o_144_sv2v_reg <= 1'b0;
      data_o_143_sv2v_reg <= 1'b0;
      data_o_142_sv2v_reg <= 1'b0;
      data_o_141_sv2v_reg <= 1'b0;
      data_o_140_sv2v_reg <= 1'b0;
      data_o_139_sv2v_reg <= 1'b0;
      data_o_138_sv2v_reg <= 1'b0;
      data_o_137_sv2v_reg <= 1'b0;
      data_o_136_sv2v_reg <= 1'b0;
      data_o_135_sv2v_reg <= 1'b0;
      data_o_134_sv2v_reg <= 1'b0;
      data_o_133_sv2v_reg <= 1'b0;
      data_o_132_sv2v_reg <= 1'b0;
      data_o_131_sv2v_reg <= 1'b0;
      data_o_130_sv2v_reg <= 1'b0;
      data_o_129_sv2v_reg <= 1'b0;
      data_o_128_sv2v_reg <= 1'b0;
      data_o_127_sv2v_reg <= 1'b0;
      data_o_126_sv2v_reg <= 1'b0;
      data_o_125_sv2v_reg <= 1'b0;
      data_o_124_sv2v_reg <= 1'b0;
      data_o_123_sv2v_reg <= 1'b0;
      data_o_122_sv2v_reg <= 1'b0;
      data_o_121_sv2v_reg <= 1'b0;
      data_o_120_sv2v_reg <= 1'b0;
      data_o_119_sv2v_reg <= 1'b0;
      data_o_118_sv2v_reg <= 1'b0;
      data_o_117_sv2v_reg <= 1'b0;
      data_o_116_sv2v_reg <= 1'b0;
      data_o_115_sv2v_reg <= 1'b0;
      data_o_114_sv2v_reg <= 1'b0;
      data_o_113_sv2v_reg <= 1'b0;
      data_o_112_sv2v_reg <= 1'b0;
      data_o_111_sv2v_reg <= 1'b0;
      data_o_110_sv2v_reg <= 1'b0;
      data_o_109_sv2v_reg <= 1'b0;
      data_o_108_sv2v_reg <= 1'b0;
      data_o_107_sv2v_reg <= 1'b0;
      data_o_106_sv2v_reg <= 1'b0;
      data_o_105_sv2v_reg <= 1'b0;
      data_o_104_sv2v_reg <= 1'b0;
      data_o_103_sv2v_reg <= 1'b0;
      data_o_102_sv2v_reg <= 1'b0;
      data_o_101_sv2v_reg <= 1'b0;
      data_o_100_sv2v_reg <= 1'b0;
      data_o_99_sv2v_reg <= 1'b0;
      data_o_98_sv2v_reg <= 1'b0;
      data_o_97_sv2v_reg <= 1'b0;
      data_o_96_sv2v_reg <= 1'b0;
      data_o_95_sv2v_reg <= 1'b0;
      data_o_94_sv2v_reg <= 1'b0;
      data_o_93_sv2v_reg <= 1'b0;
      data_o_92_sv2v_reg <= 1'b0;
      data_o_91_sv2v_reg <= 1'b0;
      data_o_90_sv2v_reg <= 1'b0;
      data_o_89_sv2v_reg <= 1'b0;
      data_o_88_sv2v_reg <= 1'b0;
      data_o_87_sv2v_reg <= 1'b0;
      data_o_86_sv2v_reg <= 1'b0;
      data_o_85_sv2v_reg <= 1'b0;
      data_o_84_sv2v_reg <= 1'b0;
      data_o_83_sv2v_reg <= 1'b0;
      data_o_82_sv2v_reg <= 1'b0;
      data_o_81_sv2v_reg <= 1'b0;
      data_o_80_sv2v_reg <= 1'b0;
      data_o_79_sv2v_reg <= 1'b0;
      data_o_78_sv2v_reg <= 1'b0;
      data_o_77_sv2v_reg <= 1'b0;
      data_o_76_sv2v_reg <= 1'b0;
      data_o_75_sv2v_reg <= 1'b0;
      data_o_74_sv2v_reg <= 1'b0;
      data_o_73_sv2v_reg <= 1'b0;
      data_o_72_sv2v_reg <= 1'b0;
      data_o_71_sv2v_reg <= 1'b0;
      data_o_70_sv2v_reg <= 1'b0;
      data_o_69_sv2v_reg <= 1'b0;
      data_o_68_sv2v_reg <= 1'b0;
      data_o_67_sv2v_reg <= 1'b0;
      data_o_66_sv2v_reg <= 1'b0;
      data_o_65_sv2v_reg <= 1'b0;
      data_o_64_sv2v_reg <= 1'b0;
      data_o_63_sv2v_reg <= 1'b0;
      data_o_62_sv2v_reg <= 1'b0;
      data_o_61_sv2v_reg <= 1'b0;
      data_o_60_sv2v_reg <= 1'b0;
      data_o_59_sv2v_reg <= 1'b0;
      data_o_58_sv2v_reg <= 1'b0;
      data_o_57_sv2v_reg <= 1'b0;
      data_o_56_sv2v_reg <= 1'b0;
      data_o_55_sv2v_reg <= 1'b0;
      data_o_54_sv2v_reg <= 1'b0;
      data_o_53_sv2v_reg <= 1'b0;
      data_o_52_sv2v_reg <= 1'b0;
      data_o_51_sv2v_reg <= 1'b0;
      data_o_50_sv2v_reg <= 1'b0;
      data_o_49_sv2v_reg <= 1'b0;
      data_o_48_sv2v_reg <= 1'b0;
      data_o_47_sv2v_reg <= 1'b0;
      data_o_46_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
    end else if(N6) begin
      data_o_144_sv2v_reg <= data_i[144];
      data_o_143_sv2v_reg <= data_i[143];
      data_o_142_sv2v_reg <= data_i[142];
      data_o_141_sv2v_reg <= data_i[141];
      data_o_140_sv2v_reg <= data_i[140];
      data_o_139_sv2v_reg <= data_i[139];
      data_o_138_sv2v_reg <= data_i[138];
      data_o_137_sv2v_reg <= data_i[137];
      data_o_136_sv2v_reg <= data_i[136];
      data_o_135_sv2v_reg <= data_i[135];
      data_o_134_sv2v_reg <= data_i[134];
      data_o_133_sv2v_reg <= data_i[133];
      data_o_132_sv2v_reg <= data_i[132];
      data_o_131_sv2v_reg <= data_i[131];
      data_o_130_sv2v_reg <= data_i[130];
      data_o_129_sv2v_reg <= data_i[129];
      data_o_128_sv2v_reg <= data_i[128];
      data_o_127_sv2v_reg <= data_i[127];
      data_o_126_sv2v_reg <= data_i[126];
      data_o_125_sv2v_reg <= data_i[125];
      data_o_124_sv2v_reg <= data_i[124];
      data_o_123_sv2v_reg <= data_i[123];
      data_o_122_sv2v_reg <= data_i[122];
      data_o_121_sv2v_reg <= data_i[121];
      data_o_120_sv2v_reg <= data_i[120];
      data_o_119_sv2v_reg <= data_i[119];
      data_o_118_sv2v_reg <= data_i[118];
      data_o_117_sv2v_reg <= data_i[117];
      data_o_116_sv2v_reg <= data_i[116];
      data_o_115_sv2v_reg <= data_i[115];
      data_o_114_sv2v_reg <= data_i[114];
      data_o_113_sv2v_reg <= data_i[113];
      data_o_112_sv2v_reg <= data_i[112];
      data_o_111_sv2v_reg <= data_i[111];
      data_o_110_sv2v_reg <= data_i[110];
      data_o_109_sv2v_reg <= data_i[109];
      data_o_108_sv2v_reg <= data_i[108];
      data_o_107_sv2v_reg <= data_i[107];
      data_o_106_sv2v_reg <= data_i[106];
      data_o_105_sv2v_reg <= data_i[105];
      data_o_104_sv2v_reg <= data_i[104];
      data_o_103_sv2v_reg <= data_i[103];
      data_o_102_sv2v_reg <= data_i[102];
      data_o_101_sv2v_reg <= data_i[101];
      data_o_100_sv2v_reg <= data_i[100];
      data_o_99_sv2v_reg <= data_i[99];
      data_o_98_sv2v_reg <= data_i[98];
      data_o_97_sv2v_reg <= data_i[97];
      data_o_96_sv2v_reg <= data_i[96];
      data_o_95_sv2v_reg <= data_i[95];
      data_o_94_sv2v_reg <= data_i[94];
      data_o_93_sv2v_reg <= data_i[93];
      data_o_92_sv2v_reg <= data_i[92];
      data_o_91_sv2v_reg <= data_i[91];
      data_o_90_sv2v_reg <= data_i[90];
      data_o_89_sv2v_reg <= data_i[89];
      data_o_88_sv2v_reg <= data_i[88];
      data_o_87_sv2v_reg <= data_i[87];
      data_o_86_sv2v_reg <= data_i[86];
      data_o_85_sv2v_reg <= data_i[85];
      data_o_84_sv2v_reg <= data_i[84];
      data_o_83_sv2v_reg <= data_i[83];
      data_o_82_sv2v_reg <= data_i[82];
      data_o_81_sv2v_reg <= data_i[81];
      data_o_80_sv2v_reg <= data_i[80];
      data_o_79_sv2v_reg <= data_i[79];
      data_o_78_sv2v_reg <= data_i[78];
      data_o_77_sv2v_reg <= data_i[77];
      data_o_76_sv2v_reg <= data_i[76];
      data_o_75_sv2v_reg <= data_i[75];
      data_o_74_sv2v_reg <= data_i[74];
      data_o_73_sv2v_reg <= data_i[73];
      data_o_72_sv2v_reg <= data_i[72];
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_4_sv2v_reg <= data_i[4];
    end 
    if(reset_i) begin
      data_o_45_sv2v_reg <= 1'b0;
      data_o_44_sv2v_reg <= 1'b0;
      data_o_43_sv2v_reg <= 1'b0;
      data_o_42_sv2v_reg <= 1'b0;
      data_o_41_sv2v_reg <= 1'b0;
      data_o_40_sv2v_reg <= 1'b0;
      data_o_39_sv2v_reg <= 1'b0;
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
    end else if(N7) begin
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
    end 
  end


endmodule



module bsg_dff_en_00000028
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [39:0] data_i;
  output [39:0] data_o;
  input clk_i;
  input en_i;
  wire [39:0] data_o;
  reg data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,
  data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,
  data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,
  data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,
  data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_adder_one_hot_00000008
(
  a_i,
  b_i,
  o
);

  input [7:0] a_i;
  input [7:0] b_i;
  output [7:0] o;
  wire [7:0] o,\rof_0_.aggregate ,\rof_1_.aggregate ,\rof_2_.aggregate ,\rof_3_.aggregate ,
  \rof_4_.aggregate ,\rof_5_.aggregate ,\rof_6_.aggregate ,\rof_7_.aggregate ;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47;
  assign \rof_0_.aggregate [0] = a_i[0] & b_i[0];
  assign \rof_0_.aggregate [1] = a_i[1] & b_i[7];
  assign \rof_0_.aggregate [2] = a_i[2] & b_i[6];
  assign \rof_0_.aggregate [3] = a_i[3] & b_i[5];
  assign \rof_0_.aggregate [4] = a_i[4] & b_i[4];
  assign \rof_0_.aggregate [5] = a_i[5] & b_i[3];
  assign \rof_0_.aggregate [6] = a_i[6] & b_i[2];
  assign \rof_0_.aggregate [7] = a_i[7] & b_i[1];
  assign o[0] = N5 | \rof_0_.aggregate [0];
  assign N5 = N4 | \rof_0_.aggregate [1];
  assign N4 = N3 | \rof_0_.aggregate [2];
  assign N3 = N2 | \rof_0_.aggregate [3];
  assign N2 = N1 | \rof_0_.aggregate [4];
  assign N1 = N0 | \rof_0_.aggregate [5];
  assign N0 = \rof_0_.aggregate [7] | \rof_0_.aggregate [6];
  assign \rof_1_.aggregate [0] = a_i[0] & b_i[1];
  assign \rof_1_.aggregate [1] = a_i[1] & b_i[0];
  assign \rof_1_.aggregate [2] = a_i[2] & b_i[7];
  assign \rof_1_.aggregate [3] = a_i[3] & b_i[6];
  assign \rof_1_.aggregate [4] = a_i[4] & b_i[5];
  assign \rof_1_.aggregate [5] = a_i[5] & b_i[4];
  assign \rof_1_.aggregate [6] = a_i[6] & b_i[3];
  assign \rof_1_.aggregate [7] = a_i[7] & b_i[2];
  assign o[1] = N11 | \rof_1_.aggregate [0];
  assign N11 = N10 | \rof_1_.aggregate [1];
  assign N10 = N9 | \rof_1_.aggregate [2];
  assign N9 = N8 | \rof_1_.aggregate [3];
  assign N8 = N7 | \rof_1_.aggregate [4];
  assign N7 = N6 | \rof_1_.aggregate [5];
  assign N6 = \rof_1_.aggregate [7] | \rof_1_.aggregate [6];
  assign \rof_2_.aggregate [0] = a_i[0] & b_i[2];
  assign \rof_2_.aggregate [1] = a_i[1] & b_i[1];
  assign \rof_2_.aggregate [2] = a_i[2] & b_i[0];
  assign \rof_2_.aggregate [3] = a_i[3] & b_i[7];
  assign \rof_2_.aggregate [4] = a_i[4] & b_i[6];
  assign \rof_2_.aggregate [5] = a_i[5] & b_i[5];
  assign \rof_2_.aggregate [6] = a_i[6] & b_i[4];
  assign \rof_2_.aggregate [7] = a_i[7] & b_i[3];
  assign o[2] = N17 | \rof_2_.aggregate [0];
  assign N17 = N16 | \rof_2_.aggregate [1];
  assign N16 = N15 | \rof_2_.aggregate [2];
  assign N15 = N14 | \rof_2_.aggregate [3];
  assign N14 = N13 | \rof_2_.aggregate [4];
  assign N13 = N12 | \rof_2_.aggregate [5];
  assign N12 = \rof_2_.aggregate [7] | \rof_2_.aggregate [6];
  assign \rof_3_.aggregate [0] = a_i[0] & b_i[3];
  assign \rof_3_.aggregate [1] = a_i[1] & b_i[2];
  assign \rof_3_.aggregate [2] = a_i[2] & b_i[1];
  assign \rof_3_.aggregate [3] = a_i[3] & b_i[0];
  assign \rof_3_.aggregate [4] = a_i[4] & b_i[7];
  assign \rof_3_.aggregate [5] = a_i[5] & b_i[6];
  assign \rof_3_.aggregate [6] = a_i[6] & b_i[5];
  assign \rof_3_.aggregate [7] = a_i[7] & b_i[4];
  assign o[3] = N23 | \rof_3_.aggregate [0];
  assign N23 = N22 | \rof_3_.aggregate [1];
  assign N22 = N21 | \rof_3_.aggregate [2];
  assign N21 = N20 | \rof_3_.aggregate [3];
  assign N20 = N19 | \rof_3_.aggregate [4];
  assign N19 = N18 | \rof_3_.aggregate [5];
  assign N18 = \rof_3_.aggregate [7] | \rof_3_.aggregate [6];
  assign \rof_4_.aggregate [0] = a_i[0] & b_i[4];
  assign \rof_4_.aggregate [1] = a_i[1] & b_i[3];
  assign \rof_4_.aggregate [2] = a_i[2] & b_i[2];
  assign \rof_4_.aggregate [3] = a_i[3] & b_i[1];
  assign \rof_4_.aggregate [4] = a_i[4] & b_i[0];
  assign \rof_4_.aggregate [5] = a_i[5] & b_i[7];
  assign \rof_4_.aggregate [6] = a_i[6] & b_i[6];
  assign \rof_4_.aggregate [7] = a_i[7] & b_i[5];
  assign o[4] = N29 | \rof_4_.aggregate [0];
  assign N29 = N28 | \rof_4_.aggregate [1];
  assign N28 = N27 | \rof_4_.aggregate [2];
  assign N27 = N26 | \rof_4_.aggregate [3];
  assign N26 = N25 | \rof_4_.aggregate [4];
  assign N25 = N24 | \rof_4_.aggregate [5];
  assign N24 = \rof_4_.aggregate [7] | \rof_4_.aggregate [6];
  assign \rof_5_.aggregate [0] = a_i[0] & b_i[5];
  assign \rof_5_.aggregate [1] = a_i[1] & b_i[4];
  assign \rof_5_.aggregate [2] = a_i[2] & b_i[3];
  assign \rof_5_.aggregate [3] = a_i[3] & b_i[2];
  assign \rof_5_.aggregate [4] = a_i[4] & b_i[1];
  assign \rof_5_.aggregate [5] = a_i[5] & b_i[0];
  assign \rof_5_.aggregate [6] = a_i[6] & b_i[7];
  assign \rof_5_.aggregate [7] = a_i[7] & b_i[6];
  assign o[5] = N35 | \rof_5_.aggregate [0];
  assign N35 = N34 | \rof_5_.aggregate [1];
  assign N34 = N33 | \rof_5_.aggregate [2];
  assign N33 = N32 | \rof_5_.aggregate [3];
  assign N32 = N31 | \rof_5_.aggregate [4];
  assign N31 = N30 | \rof_5_.aggregate [5];
  assign N30 = \rof_5_.aggregate [7] | \rof_5_.aggregate [6];
  assign \rof_6_.aggregate [0] = a_i[0] & b_i[6];
  assign \rof_6_.aggregate [1] = a_i[1] & b_i[5];
  assign \rof_6_.aggregate [2] = a_i[2] & b_i[4];
  assign \rof_6_.aggregate [3] = a_i[3] & b_i[3];
  assign \rof_6_.aggregate [4] = a_i[4] & b_i[2];
  assign \rof_6_.aggregate [5] = a_i[5] & b_i[1];
  assign \rof_6_.aggregate [6] = a_i[6] & b_i[0];
  assign \rof_6_.aggregate [7] = a_i[7] & b_i[7];
  assign o[6] = N41 | \rof_6_.aggregate [0];
  assign N41 = N40 | \rof_6_.aggregate [1];
  assign N40 = N39 | \rof_6_.aggregate [2];
  assign N39 = N38 | \rof_6_.aggregate [3];
  assign N38 = N37 | \rof_6_.aggregate [4];
  assign N37 = N36 | \rof_6_.aggregate [5];
  assign N36 = \rof_6_.aggregate [7] | \rof_6_.aggregate [6];
  assign \rof_7_.aggregate [0] = a_i[0] & b_i[7];
  assign \rof_7_.aggregate [1] = a_i[1] & b_i[6];
  assign \rof_7_.aggregate [2] = a_i[2] & b_i[5];
  assign \rof_7_.aggregate [3] = a_i[3] & b_i[4];
  assign \rof_7_.aggregate [4] = a_i[4] & b_i[3];
  assign \rof_7_.aggregate [5] = a_i[5] & b_i[2];
  assign \rof_7_.aggregate [6] = a_i[6] & b_i[1];
  assign \rof_7_.aggregate [7] = a_i[7] & b_i[0];
  assign o[7] = N47 | \rof_7_.aggregate [0];
  assign N47 = N46 | \rof_7_.aggregate [1];
  assign N46 = N45 | \rof_7_.aggregate [2];
  assign N45 = N44 | \rof_7_.aggregate [3];
  assign N44 = N43 | \rof_7_.aggregate [4];
  assign N43 = N42 | \rof_7_.aggregate [5];
  assign N42 = \rof_7_.aggregate [7] | \rof_7_.aggregate [6];

endmodule



module bsg_mux_one_hot_00000040_00000008
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [511:0] data_i;
  input [7:0] sel_one_hot_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383;
  wire [511:0] data_masked;
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[1];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[1];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[1];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[2];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[2];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[2];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[2];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[2];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[2];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[2];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[2];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[2];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[2];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[2];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[2];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[2];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[2];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[2];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[2];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[2];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[2];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[2];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[2];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[2];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[2];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[2];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[2];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[2];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[2];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[2];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[2];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[2];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[2];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[2];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[2];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[2];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[2];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[2];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[2];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[2];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[2];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[2];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[2];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[2];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[2];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[2];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[2];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[2];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[2];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[2];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[2];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[2];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[2];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[2];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[2];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[2];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[2];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[2];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[2];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[2];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[2];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[2];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[2];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[2];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[2];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[2];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[2];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[3];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[3];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[3];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[3];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[3];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[3];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[3];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[3];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[3];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[3];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[3];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[3];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[3];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[3];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[3];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[3];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[3];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[3];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[3];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[3];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[3];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[3];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[3];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[3];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[3];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[3];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[3];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[3];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[3];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[3];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[3];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[3];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[3];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[3];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[3];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[3];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[3];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[3];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[3];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[3];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[3];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[3];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[3];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[3];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[3];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[3];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[3];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[3];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[3];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[3];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[3];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[3];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[3];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[3];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[3];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[3];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[3];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[3];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[3];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[3];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[3];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[3];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[3];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[3];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[4];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[4];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[4];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[4];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[4];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[4];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[4];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[4];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[4];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[4];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[4];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[4];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[4];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[4];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[4];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[4];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[4];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[4];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[4];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[4];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[4];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[4];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[4];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[4];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[4];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[4];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[4];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[4];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[4];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[4];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[4];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[4];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[4];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[4];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[4];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[4];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[4];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[4];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[4];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[4];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[4];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[4];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[4];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[4];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[4];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[4];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[4];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[4];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[4];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[4];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[4];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[4];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[4];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[4];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[4];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[4];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[4];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[4];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[4];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[4];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[4];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[4];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[4];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[4];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[5];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[5];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[5];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[5];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[5];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[5];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[5];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[5];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[5];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[5];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[5];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[5];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[5];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[5];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[5];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[5];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[5];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[5];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[5];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[5];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[5];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[5];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[5];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[5];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[5];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[5];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[5];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[5];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[5];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[5];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[5];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[5];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[5];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[5];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[5];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[5];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[5];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[5];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[5];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[5];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[5];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[5];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[5];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[5];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[5];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[5];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[5];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[5];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[5];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[5];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[5];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[5];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[5];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[5];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[5];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[5];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[5];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[5];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[5];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[5];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[5];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[5];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[5];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[5];
  assign data_masked[447] = data_i[447] & sel_one_hot_i[6];
  assign data_masked[446] = data_i[446] & sel_one_hot_i[6];
  assign data_masked[445] = data_i[445] & sel_one_hot_i[6];
  assign data_masked[444] = data_i[444] & sel_one_hot_i[6];
  assign data_masked[443] = data_i[443] & sel_one_hot_i[6];
  assign data_masked[442] = data_i[442] & sel_one_hot_i[6];
  assign data_masked[441] = data_i[441] & sel_one_hot_i[6];
  assign data_masked[440] = data_i[440] & sel_one_hot_i[6];
  assign data_masked[439] = data_i[439] & sel_one_hot_i[6];
  assign data_masked[438] = data_i[438] & sel_one_hot_i[6];
  assign data_masked[437] = data_i[437] & sel_one_hot_i[6];
  assign data_masked[436] = data_i[436] & sel_one_hot_i[6];
  assign data_masked[435] = data_i[435] & sel_one_hot_i[6];
  assign data_masked[434] = data_i[434] & sel_one_hot_i[6];
  assign data_masked[433] = data_i[433] & sel_one_hot_i[6];
  assign data_masked[432] = data_i[432] & sel_one_hot_i[6];
  assign data_masked[431] = data_i[431] & sel_one_hot_i[6];
  assign data_masked[430] = data_i[430] & sel_one_hot_i[6];
  assign data_masked[429] = data_i[429] & sel_one_hot_i[6];
  assign data_masked[428] = data_i[428] & sel_one_hot_i[6];
  assign data_masked[427] = data_i[427] & sel_one_hot_i[6];
  assign data_masked[426] = data_i[426] & sel_one_hot_i[6];
  assign data_masked[425] = data_i[425] & sel_one_hot_i[6];
  assign data_masked[424] = data_i[424] & sel_one_hot_i[6];
  assign data_masked[423] = data_i[423] & sel_one_hot_i[6];
  assign data_masked[422] = data_i[422] & sel_one_hot_i[6];
  assign data_masked[421] = data_i[421] & sel_one_hot_i[6];
  assign data_masked[420] = data_i[420] & sel_one_hot_i[6];
  assign data_masked[419] = data_i[419] & sel_one_hot_i[6];
  assign data_masked[418] = data_i[418] & sel_one_hot_i[6];
  assign data_masked[417] = data_i[417] & sel_one_hot_i[6];
  assign data_masked[416] = data_i[416] & sel_one_hot_i[6];
  assign data_masked[415] = data_i[415] & sel_one_hot_i[6];
  assign data_masked[414] = data_i[414] & sel_one_hot_i[6];
  assign data_masked[413] = data_i[413] & sel_one_hot_i[6];
  assign data_masked[412] = data_i[412] & sel_one_hot_i[6];
  assign data_masked[411] = data_i[411] & sel_one_hot_i[6];
  assign data_masked[410] = data_i[410] & sel_one_hot_i[6];
  assign data_masked[409] = data_i[409] & sel_one_hot_i[6];
  assign data_masked[408] = data_i[408] & sel_one_hot_i[6];
  assign data_masked[407] = data_i[407] & sel_one_hot_i[6];
  assign data_masked[406] = data_i[406] & sel_one_hot_i[6];
  assign data_masked[405] = data_i[405] & sel_one_hot_i[6];
  assign data_masked[404] = data_i[404] & sel_one_hot_i[6];
  assign data_masked[403] = data_i[403] & sel_one_hot_i[6];
  assign data_masked[402] = data_i[402] & sel_one_hot_i[6];
  assign data_masked[401] = data_i[401] & sel_one_hot_i[6];
  assign data_masked[400] = data_i[400] & sel_one_hot_i[6];
  assign data_masked[399] = data_i[399] & sel_one_hot_i[6];
  assign data_masked[398] = data_i[398] & sel_one_hot_i[6];
  assign data_masked[397] = data_i[397] & sel_one_hot_i[6];
  assign data_masked[396] = data_i[396] & sel_one_hot_i[6];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[6];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[6];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[6];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[6];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[6];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[6];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[6];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[6];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[6];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[6];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[6];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[6];
  assign data_masked[511] = data_i[511] & sel_one_hot_i[7];
  assign data_masked[510] = data_i[510] & sel_one_hot_i[7];
  assign data_masked[509] = data_i[509] & sel_one_hot_i[7];
  assign data_masked[508] = data_i[508] & sel_one_hot_i[7];
  assign data_masked[507] = data_i[507] & sel_one_hot_i[7];
  assign data_masked[506] = data_i[506] & sel_one_hot_i[7];
  assign data_masked[505] = data_i[505] & sel_one_hot_i[7];
  assign data_masked[504] = data_i[504] & sel_one_hot_i[7];
  assign data_masked[503] = data_i[503] & sel_one_hot_i[7];
  assign data_masked[502] = data_i[502] & sel_one_hot_i[7];
  assign data_masked[501] = data_i[501] & sel_one_hot_i[7];
  assign data_masked[500] = data_i[500] & sel_one_hot_i[7];
  assign data_masked[499] = data_i[499] & sel_one_hot_i[7];
  assign data_masked[498] = data_i[498] & sel_one_hot_i[7];
  assign data_masked[497] = data_i[497] & sel_one_hot_i[7];
  assign data_masked[496] = data_i[496] & sel_one_hot_i[7];
  assign data_masked[495] = data_i[495] & sel_one_hot_i[7];
  assign data_masked[494] = data_i[494] & sel_one_hot_i[7];
  assign data_masked[493] = data_i[493] & sel_one_hot_i[7];
  assign data_masked[492] = data_i[492] & sel_one_hot_i[7];
  assign data_masked[491] = data_i[491] & sel_one_hot_i[7];
  assign data_masked[490] = data_i[490] & sel_one_hot_i[7];
  assign data_masked[489] = data_i[489] & sel_one_hot_i[7];
  assign data_masked[488] = data_i[488] & sel_one_hot_i[7];
  assign data_masked[487] = data_i[487] & sel_one_hot_i[7];
  assign data_masked[486] = data_i[486] & sel_one_hot_i[7];
  assign data_masked[485] = data_i[485] & sel_one_hot_i[7];
  assign data_masked[484] = data_i[484] & sel_one_hot_i[7];
  assign data_masked[483] = data_i[483] & sel_one_hot_i[7];
  assign data_masked[482] = data_i[482] & sel_one_hot_i[7];
  assign data_masked[481] = data_i[481] & sel_one_hot_i[7];
  assign data_masked[480] = data_i[480] & sel_one_hot_i[7];
  assign data_masked[479] = data_i[479] & sel_one_hot_i[7];
  assign data_masked[478] = data_i[478] & sel_one_hot_i[7];
  assign data_masked[477] = data_i[477] & sel_one_hot_i[7];
  assign data_masked[476] = data_i[476] & sel_one_hot_i[7];
  assign data_masked[475] = data_i[475] & sel_one_hot_i[7];
  assign data_masked[474] = data_i[474] & sel_one_hot_i[7];
  assign data_masked[473] = data_i[473] & sel_one_hot_i[7];
  assign data_masked[472] = data_i[472] & sel_one_hot_i[7];
  assign data_masked[471] = data_i[471] & sel_one_hot_i[7];
  assign data_masked[470] = data_i[470] & sel_one_hot_i[7];
  assign data_masked[469] = data_i[469] & sel_one_hot_i[7];
  assign data_masked[468] = data_i[468] & sel_one_hot_i[7];
  assign data_masked[467] = data_i[467] & sel_one_hot_i[7];
  assign data_masked[466] = data_i[466] & sel_one_hot_i[7];
  assign data_masked[465] = data_i[465] & sel_one_hot_i[7];
  assign data_masked[464] = data_i[464] & sel_one_hot_i[7];
  assign data_masked[463] = data_i[463] & sel_one_hot_i[7];
  assign data_masked[462] = data_i[462] & sel_one_hot_i[7];
  assign data_masked[461] = data_i[461] & sel_one_hot_i[7];
  assign data_masked[460] = data_i[460] & sel_one_hot_i[7];
  assign data_masked[459] = data_i[459] & sel_one_hot_i[7];
  assign data_masked[458] = data_i[458] & sel_one_hot_i[7];
  assign data_masked[457] = data_i[457] & sel_one_hot_i[7];
  assign data_masked[456] = data_i[456] & sel_one_hot_i[7];
  assign data_masked[455] = data_i[455] & sel_one_hot_i[7];
  assign data_masked[454] = data_i[454] & sel_one_hot_i[7];
  assign data_masked[453] = data_i[453] & sel_one_hot_i[7];
  assign data_masked[452] = data_i[452] & sel_one_hot_i[7];
  assign data_masked[451] = data_i[451] & sel_one_hot_i[7];
  assign data_masked[450] = data_i[450] & sel_one_hot_i[7];
  assign data_masked[449] = data_i[449] & sel_one_hot_i[7];
  assign data_masked[448] = data_i[448] & sel_one_hot_i[7];
  assign data_o[0] = N5 | data_masked[0];
  assign N5 = N4 | data_masked[64];
  assign N4 = N3 | data_masked[128];
  assign N3 = N2 | data_masked[192];
  assign N2 = N1 | data_masked[256];
  assign N1 = N0 | data_masked[320];
  assign N0 = data_masked[448] | data_masked[384];
  assign data_o[1] = N11 | data_masked[1];
  assign N11 = N10 | data_masked[65];
  assign N10 = N9 | data_masked[129];
  assign N9 = N8 | data_masked[193];
  assign N8 = N7 | data_masked[257];
  assign N7 = N6 | data_masked[321];
  assign N6 = data_masked[449] | data_masked[385];
  assign data_o[2] = N17 | data_masked[2];
  assign N17 = N16 | data_masked[66];
  assign N16 = N15 | data_masked[130];
  assign N15 = N14 | data_masked[194];
  assign N14 = N13 | data_masked[258];
  assign N13 = N12 | data_masked[322];
  assign N12 = data_masked[450] | data_masked[386];
  assign data_o[3] = N23 | data_masked[3];
  assign N23 = N22 | data_masked[67];
  assign N22 = N21 | data_masked[131];
  assign N21 = N20 | data_masked[195];
  assign N20 = N19 | data_masked[259];
  assign N19 = N18 | data_masked[323];
  assign N18 = data_masked[451] | data_masked[387];
  assign data_o[4] = N29 | data_masked[4];
  assign N29 = N28 | data_masked[68];
  assign N28 = N27 | data_masked[132];
  assign N27 = N26 | data_masked[196];
  assign N26 = N25 | data_masked[260];
  assign N25 = N24 | data_masked[324];
  assign N24 = data_masked[452] | data_masked[388];
  assign data_o[5] = N35 | data_masked[5];
  assign N35 = N34 | data_masked[69];
  assign N34 = N33 | data_masked[133];
  assign N33 = N32 | data_masked[197];
  assign N32 = N31 | data_masked[261];
  assign N31 = N30 | data_masked[325];
  assign N30 = data_masked[453] | data_masked[389];
  assign data_o[6] = N41 | data_masked[6];
  assign N41 = N40 | data_masked[70];
  assign N40 = N39 | data_masked[134];
  assign N39 = N38 | data_masked[198];
  assign N38 = N37 | data_masked[262];
  assign N37 = N36 | data_masked[326];
  assign N36 = data_masked[454] | data_masked[390];
  assign data_o[7] = N47 | data_masked[7];
  assign N47 = N46 | data_masked[71];
  assign N46 = N45 | data_masked[135];
  assign N45 = N44 | data_masked[199];
  assign N44 = N43 | data_masked[263];
  assign N43 = N42 | data_masked[327];
  assign N42 = data_masked[455] | data_masked[391];
  assign data_o[8] = N53 | data_masked[8];
  assign N53 = N52 | data_masked[72];
  assign N52 = N51 | data_masked[136];
  assign N51 = N50 | data_masked[200];
  assign N50 = N49 | data_masked[264];
  assign N49 = N48 | data_masked[328];
  assign N48 = data_masked[456] | data_masked[392];
  assign data_o[9] = N59 | data_masked[9];
  assign N59 = N58 | data_masked[73];
  assign N58 = N57 | data_masked[137];
  assign N57 = N56 | data_masked[201];
  assign N56 = N55 | data_masked[265];
  assign N55 = N54 | data_masked[329];
  assign N54 = data_masked[457] | data_masked[393];
  assign data_o[10] = N65 | data_masked[10];
  assign N65 = N64 | data_masked[74];
  assign N64 = N63 | data_masked[138];
  assign N63 = N62 | data_masked[202];
  assign N62 = N61 | data_masked[266];
  assign N61 = N60 | data_masked[330];
  assign N60 = data_masked[458] | data_masked[394];
  assign data_o[11] = N71 | data_masked[11];
  assign N71 = N70 | data_masked[75];
  assign N70 = N69 | data_masked[139];
  assign N69 = N68 | data_masked[203];
  assign N68 = N67 | data_masked[267];
  assign N67 = N66 | data_masked[331];
  assign N66 = data_masked[459] | data_masked[395];
  assign data_o[12] = N77 | data_masked[12];
  assign N77 = N76 | data_masked[76];
  assign N76 = N75 | data_masked[140];
  assign N75 = N74 | data_masked[204];
  assign N74 = N73 | data_masked[268];
  assign N73 = N72 | data_masked[332];
  assign N72 = data_masked[460] | data_masked[396];
  assign data_o[13] = N83 | data_masked[13];
  assign N83 = N82 | data_masked[77];
  assign N82 = N81 | data_masked[141];
  assign N81 = N80 | data_masked[205];
  assign N80 = N79 | data_masked[269];
  assign N79 = N78 | data_masked[333];
  assign N78 = data_masked[461] | data_masked[397];
  assign data_o[14] = N89 | data_masked[14];
  assign N89 = N88 | data_masked[78];
  assign N88 = N87 | data_masked[142];
  assign N87 = N86 | data_masked[206];
  assign N86 = N85 | data_masked[270];
  assign N85 = N84 | data_masked[334];
  assign N84 = data_masked[462] | data_masked[398];
  assign data_o[15] = N95 | data_masked[15];
  assign N95 = N94 | data_masked[79];
  assign N94 = N93 | data_masked[143];
  assign N93 = N92 | data_masked[207];
  assign N92 = N91 | data_masked[271];
  assign N91 = N90 | data_masked[335];
  assign N90 = data_masked[463] | data_masked[399];
  assign data_o[16] = N101 | data_masked[16];
  assign N101 = N100 | data_masked[80];
  assign N100 = N99 | data_masked[144];
  assign N99 = N98 | data_masked[208];
  assign N98 = N97 | data_masked[272];
  assign N97 = N96 | data_masked[336];
  assign N96 = data_masked[464] | data_masked[400];
  assign data_o[17] = N107 | data_masked[17];
  assign N107 = N106 | data_masked[81];
  assign N106 = N105 | data_masked[145];
  assign N105 = N104 | data_masked[209];
  assign N104 = N103 | data_masked[273];
  assign N103 = N102 | data_masked[337];
  assign N102 = data_masked[465] | data_masked[401];
  assign data_o[18] = N113 | data_masked[18];
  assign N113 = N112 | data_masked[82];
  assign N112 = N111 | data_masked[146];
  assign N111 = N110 | data_masked[210];
  assign N110 = N109 | data_masked[274];
  assign N109 = N108 | data_masked[338];
  assign N108 = data_masked[466] | data_masked[402];
  assign data_o[19] = N119 | data_masked[19];
  assign N119 = N118 | data_masked[83];
  assign N118 = N117 | data_masked[147];
  assign N117 = N116 | data_masked[211];
  assign N116 = N115 | data_masked[275];
  assign N115 = N114 | data_masked[339];
  assign N114 = data_masked[467] | data_masked[403];
  assign data_o[20] = N125 | data_masked[20];
  assign N125 = N124 | data_masked[84];
  assign N124 = N123 | data_masked[148];
  assign N123 = N122 | data_masked[212];
  assign N122 = N121 | data_masked[276];
  assign N121 = N120 | data_masked[340];
  assign N120 = data_masked[468] | data_masked[404];
  assign data_o[21] = N131 | data_masked[21];
  assign N131 = N130 | data_masked[85];
  assign N130 = N129 | data_masked[149];
  assign N129 = N128 | data_masked[213];
  assign N128 = N127 | data_masked[277];
  assign N127 = N126 | data_masked[341];
  assign N126 = data_masked[469] | data_masked[405];
  assign data_o[22] = N137 | data_masked[22];
  assign N137 = N136 | data_masked[86];
  assign N136 = N135 | data_masked[150];
  assign N135 = N134 | data_masked[214];
  assign N134 = N133 | data_masked[278];
  assign N133 = N132 | data_masked[342];
  assign N132 = data_masked[470] | data_masked[406];
  assign data_o[23] = N143 | data_masked[23];
  assign N143 = N142 | data_masked[87];
  assign N142 = N141 | data_masked[151];
  assign N141 = N140 | data_masked[215];
  assign N140 = N139 | data_masked[279];
  assign N139 = N138 | data_masked[343];
  assign N138 = data_masked[471] | data_masked[407];
  assign data_o[24] = N149 | data_masked[24];
  assign N149 = N148 | data_masked[88];
  assign N148 = N147 | data_masked[152];
  assign N147 = N146 | data_masked[216];
  assign N146 = N145 | data_masked[280];
  assign N145 = N144 | data_masked[344];
  assign N144 = data_masked[472] | data_masked[408];
  assign data_o[25] = N155 | data_masked[25];
  assign N155 = N154 | data_masked[89];
  assign N154 = N153 | data_masked[153];
  assign N153 = N152 | data_masked[217];
  assign N152 = N151 | data_masked[281];
  assign N151 = N150 | data_masked[345];
  assign N150 = data_masked[473] | data_masked[409];
  assign data_o[26] = N161 | data_masked[26];
  assign N161 = N160 | data_masked[90];
  assign N160 = N159 | data_masked[154];
  assign N159 = N158 | data_masked[218];
  assign N158 = N157 | data_masked[282];
  assign N157 = N156 | data_masked[346];
  assign N156 = data_masked[474] | data_masked[410];
  assign data_o[27] = N167 | data_masked[27];
  assign N167 = N166 | data_masked[91];
  assign N166 = N165 | data_masked[155];
  assign N165 = N164 | data_masked[219];
  assign N164 = N163 | data_masked[283];
  assign N163 = N162 | data_masked[347];
  assign N162 = data_masked[475] | data_masked[411];
  assign data_o[28] = N173 | data_masked[28];
  assign N173 = N172 | data_masked[92];
  assign N172 = N171 | data_masked[156];
  assign N171 = N170 | data_masked[220];
  assign N170 = N169 | data_masked[284];
  assign N169 = N168 | data_masked[348];
  assign N168 = data_masked[476] | data_masked[412];
  assign data_o[29] = N179 | data_masked[29];
  assign N179 = N178 | data_masked[93];
  assign N178 = N177 | data_masked[157];
  assign N177 = N176 | data_masked[221];
  assign N176 = N175 | data_masked[285];
  assign N175 = N174 | data_masked[349];
  assign N174 = data_masked[477] | data_masked[413];
  assign data_o[30] = N185 | data_masked[30];
  assign N185 = N184 | data_masked[94];
  assign N184 = N183 | data_masked[158];
  assign N183 = N182 | data_masked[222];
  assign N182 = N181 | data_masked[286];
  assign N181 = N180 | data_masked[350];
  assign N180 = data_masked[478] | data_masked[414];
  assign data_o[31] = N191 | data_masked[31];
  assign N191 = N190 | data_masked[95];
  assign N190 = N189 | data_masked[159];
  assign N189 = N188 | data_masked[223];
  assign N188 = N187 | data_masked[287];
  assign N187 = N186 | data_masked[351];
  assign N186 = data_masked[479] | data_masked[415];
  assign data_o[32] = N197 | data_masked[32];
  assign N197 = N196 | data_masked[96];
  assign N196 = N195 | data_masked[160];
  assign N195 = N194 | data_masked[224];
  assign N194 = N193 | data_masked[288];
  assign N193 = N192 | data_masked[352];
  assign N192 = data_masked[480] | data_masked[416];
  assign data_o[33] = N203 | data_masked[33];
  assign N203 = N202 | data_masked[97];
  assign N202 = N201 | data_masked[161];
  assign N201 = N200 | data_masked[225];
  assign N200 = N199 | data_masked[289];
  assign N199 = N198 | data_masked[353];
  assign N198 = data_masked[481] | data_masked[417];
  assign data_o[34] = N209 | data_masked[34];
  assign N209 = N208 | data_masked[98];
  assign N208 = N207 | data_masked[162];
  assign N207 = N206 | data_masked[226];
  assign N206 = N205 | data_masked[290];
  assign N205 = N204 | data_masked[354];
  assign N204 = data_masked[482] | data_masked[418];
  assign data_o[35] = N215 | data_masked[35];
  assign N215 = N214 | data_masked[99];
  assign N214 = N213 | data_masked[163];
  assign N213 = N212 | data_masked[227];
  assign N212 = N211 | data_masked[291];
  assign N211 = N210 | data_masked[355];
  assign N210 = data_masked[483] | data_masked[419];
  assign data_o[36] = N221 | data_masked[36];
  assign N221 = N220 | data_masked[100];
  assign N220 = N219 | data_masked[164];
  assign N219 = N218 | data_masked[228];
  assign N218 = N217 | data_masked[292];
  assign N217 = N216 | data_masked[356];
  assign N216 = data_masked[484] | data_masked[420];
  assign data_o[37] = N227 | data_masked[37];
  assign N227 = N226 | data_masked[101];
  assign N226 = N225 | data_masked[165];
  assign N225 = N224 | data_masked[229];
  assign N224 = N223 | data_masked[293];
  assign N223 = N222 | data_masked[357];
  assign N222 = data_masked[485] | data_masked[421];
  assign data_o[38] = N233 | data_masked[38];
  assign N233 = N232 | data_masked[102];
  assign N232 = N231 | data_masked[166];
  assign N231 = N230 | data_masked[230];
  assign N230 = N229 | data_masked[294];
  assign N229 = N228 | data_masked[358];
  assign N228 = data_masked[486] | data_masked[422];
  assign data_o[39] = N239 | data_masked[39];
  assign N239 = N238 | data_masked[103];
  assign N238 = N237 | data_masked[167];
  assign N237 = N236 | data_masked[231];
  assign N236 = N235 | data_masked[295];
  assign N235 = N234 | data_masked[359];
  assign N234 = data_masked[487] | data_masked[423];
  assign data_o[40] = N245 | data_masked[40];
  assign N245 = N244 | data_masked[104];
  assign N244 = N243 | data_masked[168];
  assign N243 = N242 | data_masked[232];
  assign N242 = N241 | data_masked[296];
  assign N241 = N240 | data_masked[360];
  assign N240 = data_masked[488] | data_masked[424];
  assign data_o[41] = N251 | data_masked[41];
  assign N251 = N250 | data_masked[105];
  assign N250 = N249 | data_masked[169];
  assign N249 = N248 | data_masked[233];
  assign N248 = N247 | data_masked[297];
  assign N247 = N246 | data_masked[361];
  assign N246 = data_masked[489] | data_masked[425];
  assign data_o[42] = N257 | data_masked[42];
  assign N257 = N256 | data_masked[106];
  assign N256 = N255 | data_masked[170];
  assign N255 = N254 | data_masked[234];
  assign N254 = N253 | data_masked[298];
  assign N253 = N252 | data_masked[362];
  assign N252 = data_masked[490] | data_masked[426];
  assign data_o[43] = N263 | data_masked[43];
  assign N263 = N262 | data_masked[107];
  assign N262 = N261 | data_masked[171];
  assign N261 = N260 | data_masked[235];
  assign N260 = N259 | data_masked[299];
  assign N259 = N258 | data_masked[363];
  assign N258 = data_masked[491] | data_masked[427];
  assign data_o[44] = N269 | data_masked[44];
  assign N269 = N268 | data_masked[108];
  assign N268 = N267 | data_masked[172];
  assign N267 = N266 | data_masked[236];
  assign N266 = N265 | data_masked[300];
  assign N265 = N264 | data_masked[364];
  assign N264 = data_masked[492] | data_masked[428];
  assign data_o[45] = N275 | data_masked[45];
  assign N275 = N274 | data_masked[109];
  assign N274 = N273 | data_masked[173];
  assign N273 = N272 | data_masked[237];
  assign N272 = N271 | data_masked[301];
  assign N271 = N270 | data_masked[365];
  assign N270 = data_masked[493] | data_masked[429];
  assign data_o[46] = N281 | data_masked[46];
  assign N281 = N280 | data_masked[110];
  assign N280 = N279 | data_masked[174];
  assign N279 = N278 | data_masked[238];
  assign N278 = N277 | data_masked[302];
  assign N277 = N276 | data_masked[366];
  assign N276 = data_masked[494] | data_masked[430];
  assign data_o[47] = N287 | data_masked[47];
  assign N287 = N286 | data_masked[111];
  assign N286 = N285 | data_masked[175];
  assign N285 = N284 | data_masked[239];
  assign N284 = N283 | data_masked[303];
  assign N283 = N282 | data_masked[367];
  assign N282 = data_masked[495] | data_masked[431];
  assign data_o[48] = N293 | data_masked[48];
  assign N293 = N292 | data_masked[112];
  assign N292 = N291 | data_masked[176];
  assign N291 = N290 | data_masked[240];
  assign N290 = N289 | data_masked[304];
  assign N289 = N288 | data_masked[368];
  assign N288 = data_masked[496] | data_masked[432];
  assign data_o[49] = N299 | data_masked[49];
  assign N299 = N298 | data_masked[113];
  assign N298 = N297 | data_masked[177];
  assign N297 = N296 | data_masked[241];
  assign N296 = N295 | data_masked[305];
  assign N295 = N294 | data_masked[369];
  assign N294 = data_masked[497] | data_masked[433];
  assign data_o[50] = N305 | data_masked[50];
  assign N305 = N304 | data_masked[114];
  assign N304 = N303 | data_masked[178];
  assign N303 = N302 | data_masked[242];
  assign N302 = N301 | data_masked[306];
  assign N301 = N300 | data_masked[370];
  assign N300 = data_masked[498] | data_masked[434];
  assign data_o[51] = N311 | data_masked[51];
  assign N311 = N310 | data_masked[115];
  assign N310 = N309 | data_masked[179];
  assign N309 = N308 | data_masked[243];
  assign N308 = N307 | data_masked[307];
  assign N307 = N306 | data_masked[371];
  assign N306 = data_masked[499] | data_masked[435];
  assign data_o[52] = N317 | data_masked[52];
  assign N317 = N316 | data_masked[116];
  assign N316 = N315 | data_masked[180];
  assign N315 = N314 | data_masked[244];
  assign N314 = N313 | data_masked[308];
  assign N313 = N312 | data_masked[372];
  assign N312 = data_masked[500] | data_masked[436];
  assign data_o[53] = N323 | data_masked[53];
  assign N323 = N322 | data_masked[117];
  assign N322 = N321 | data_masked[181];
  assign N321 = N320 | data_masked[245];
  assign N320 = N319 | data_masked[309];
  assign N319 = N318 | data_masked[373];
  assign N318 = data_masked[501] | data_masked[437];
  assign data_o[54] = N329 | data_masked[54];
  assign N329 = N328 | data_masked[118];
  assign N328 = N327 | data_masked[182];
  assign N327 = N326 | data_masked[246];
  assign N326 = N325 | data_masked[310];
  assign N325 = N324 | data_masked[374];
  assign N324 = data_masked[502] | data_masked[438];
  assign data_o[55] = N335 | data_masked[55];
  assign N335 = N334 | data_masked[119];
  assign N334 = N333 | data_masked[183];
  assign N333 = N332 | data_masked[247];
  assign N332 = N331 | data_masked[311];
  assign N331 = N330 | data_masked[375];
  assign N330 = data_masked[503] | data_masked[439];
  assign data_o[56] = N341 | data_masked[56];
  assign N341 = N340 | data_masked[120];
  assign N340 = N339 | data_masked[184];
  assign N339 = N338 | data_masked[248];
  assign N338 = N337 | data_masked[312];
  assign N337 = N336 | data_masked[376];
  assign N336 = data_masked[504] | data_masked[440];
  assign data_o[57] = N347 | data_masked[57];
  assign N347 = N346 | data_masked[121];
  assign N346 = N345 | data_masked[185];
  assign N345 = N344 | data_masked[249];
  assign N344 = N343 | data_masked[313];
  assign N343 = N342 | data_masked[377];
  assign N342 = data_masked[505] | data_masked[441];
  assign data_o[58] = N353 | data_masked[58];
  assign N353 = N352 | data_masked[122];
  assign N352 = N351 | data_masked[186];
  assign N351 = N350 | data_masked[250];
  assign N350 = N349 | data_masked[314];
  assign N349 = N348 | data_masked[378];
  assign N348 = data_masked[506] | data_masked[442];
  assign data_o[59] = N359 | data_masked[59];
  assign N359 = N358 | data_masked[123];
  assign N358 = N357 | data_masked[187];
  assign N357 = N356 | data_masked[251];
  assign N356 = N355 | data_masked[315];
  assign N355 = N354 | data_masked[379];
  assign N354 = data_masked[507] | data_masked[443];
  assign data_o[60] = N365 | data_masked[60];
  assign N365 = N364 | data_masked[124];
  assign N364 = N363 | data_masked[188];
  assign N363 = N362 | data_masked[252];
  assign N362 = N361 | data_masked[316];
  assign N361 = N360 | data_masked[380];
  assign N360 = data_masked[508] | data_masked[444];
  assign data_o[61] = N371 | data_masked[61];
  assign N371 = N370 | data_masked[125];
  assign N370 = N369 | data_masked[189];
  assign N369 = N368 | data_masked[253];
  assign N368 = N367 | data_masked[317];
  assign N367 = N366 | data_masked[381];
  assign N366 = data_masked[509] | data_masked[445];
  assign data_o[62] = N377 | data_masked[62];
  assign N377 = N376 | data_masked[126];
  assign N376 = N375 | data_masked[190];
  assign N375 = N374 | data_masked[254];
  assign N374 = N373 | data_masked[318];
  assign N373 = N372 | data_masked[382];
  assign N372 = data_masked[510] | data_masked[446];
  assign data_o[63] = N383 | data_masked[63];
  assign N383 = N382 | data_masked[127];
  assign N382 = N381 | data_masked[191];
  assign N381 = N380 | data_masked[255];
  assign N380 = N379 | data_masked[319];
  assign N379 = N378 | data_masked[383];
  assign N378 = data_masked[511] | data_masked[447];

endmodule



module bsg_mux_00000040_00000001
(
  data_i,
  sel_i,
  data_o
);

  input [63:0] data_i;
  input [0:0] sel_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  assign data_o[63] = data_i[63];
  assign data_o[62] = data_i[62];
  assign data_o[61] = data_i[61];
  assign data_o[60] = data_i[60];
  assign data_o[59] = data_i[59];
  assign data_o[58] = data_i[58];
  assign data_o[57] = data_i[57];
  assign data_o[56] = data_i[56];
  assign data_o[55] = data_i[55];
  assign data_o[54] = data_i[54];
  assign data_o[53] = data_i[53];
  assign data_o[52] = data_i[52];
  assign data_o[51] = data_i[51];
  assign data_o[50] = data_i[50];
  assign data_o[49] = data_i[49];
  assign data_o[48] = data_i[48];
  assign data_o[47] = data_i[47];
  assign data_o[46] = data_i[46];
  assign data_o[45] = data_i[45];
  assign data_o[44] = data_i[44];
  assign data_o[43] = data_i[43];
  assign data_o[42] = data_i[42];
  assign data_o[41] = data_i[41];
  assign data_o[40] = data_i[40];
  assign data_o[39] = data_i[39];
  assign data_o[38] = data_i[38];
  assign data_o[37] = data_i[37];
  assign data_o[36] = data_i[36];
  assign data_o[35] = data_i[35];
  assign data_o[34] = data_i[34];
  assign data_o[33] = data_i[33];
  assign data_o[32] = data_i[32];
  assign data_o[31] = data_i[31];
  assign data_o[30] = data_i[30];
  assign data_o[29] = data_i[29];
  assign data_o[28] = data_i[28];
  assign data_o[27] = data_i[27];
  assign data_o[26] = data_i[26];
  assign data_o[25] = data_i[25];
  assign data_o[24] = data_i[24];
  assign data_o[23] = data_i[23];
  assign data_o[22] = data_i[22];
  assign data_o[21] = data_i[21];
  assign data_o[20] = data_i[20];
  assign data_o[19] = data_i[19];
  assign data_o[18] = data_i[18];
  assign data_o[17] = data_i[17];
  assign data_o[16] = data_i[16];
  assign data_o[15] = data_i[15];
  assign data_o[14] = data_i[14];
  assign data_o[13] = data_i[13];
  assign data_o[12] = data_i[12];
  assign data_o[11] = data_i[11];
  assign data_o[10] = data_i[10];
  assign data_o[9] = data_i[9];
  assign data_o[8] = data_i[8];
  assign data_o[7] = data_i[7];
  assign data_o[6] = data_i[6];
  assign data_o[5] = data_i[5];
  assign data_o[4] = data_i[4];
  assign data_o[3] = data_i[3];
  assign data_o[2] = data_i[2];
  assign data_o[1] = data_i[1];
  assign data_o[0] = data_i[0];

endmodule



module bsg_mem_1rw_sync_mask_write_bit_00000007_00000040_1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [6:0] data_i;
  input [5:0] addr_i;
  input [6:0] w_mask_i;
  output [6:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [6:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_dff_reset_width_p1
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  wire [0:0] data_o;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_00000004
(
  clk_i,
  data_i,
  data_o
);

  input [3:0] data_i;
  output [3:0] data_o;
  input clk_i;
  wire [3:0] data_o;
  reg data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_00000003
(
  clk_i,
  data_i,
  data_o
);

  input [2:0] data_i;
  output [2:0] data_o;
  input clk_i;
  wire [2:0] data_o;
  reg data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_rotate_left_00000080
(
  data_i,
  rot_i,
  o
);

  input [127:0] data_i;
  input [6:0] rot_i;
  output [127:0] o;
  wire [127:0] o;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,
  sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,
  sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,sv2v_dc_21,sv2v_dc_22,
  sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,sv2v_dc_27,sv2v_dc_28,sv2v_dc_29,
  sv2v_dc_30,sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,sv2v_dc_34,sv2v_dc_35,sv2v_dc_36,sv2v_dc_37,
  sv2v_dc_38,sv2v_dc_39,sv2v_dc_40,sv2v_dc_41,sv2v_dc_42,sv2v_dc_43,sv2v_dc_44,
  sv2v_dc_45,sv2v_dc_46,sv2v_dc_47,sv2v_dc_48,sv2v_dc_49,sv2v_dc_50,sv2v_dc_51,
  sv2v_dc_52,sv2v_dc_53,sv2v_dc_54,sv2v_dc_55,sv2v_dc_56,sv2v_dc_57,sv2v_dc_58,sv2v_dc_59,
  sv2v_dc_60,sv2v_dc_61,sv2v_dc_62,sv2v_dc_63,sv2v_dc_64,sv2v_dc_65,sv2v_dc_66,
  sv2v_dc_67,sv2v_dc_68,sv2v_dc_69,sv2v_dc_70,sv2v_dc_71,sv2v_dc_72,sv2v_dc_73,
  sv2v_dc_74,sv2v_dc_75,sv2v_dc_76,sv2v_dc_77,sv2v_dc_78,sv2v_dc_79,sv2v_dc_80,
  sv2v_dc_81,sv2v_dc_82,sv2v_dc_83,sv2v_dc_84,sv2v_dc_85,sv2v_dc_86,sv2v_dc_87,sv2v_dc_88,
  sv2v_dc_89,sv2v_dc_90,sv2v_dc_91,sv2v_dc_92,sv2v_dc_93,sv2v_dc_94,sv2v_dc_95,
  sv2v_dc_96,sv2v_dc_97,sv2v_dc_98,sv2v_dc_99,sv2v_dc_100,sv2v_dc_101,sv2v_dc_102,
  sv2v_dc_103,sv2v_dc_104,sv2v_dc_105,sv2v_dc_106,sv2v_dc_107,sv2v_dc_108,sv2v_dc_109,
  sv2v_dc_110,sv2v_dc_111,sv2v_dc_112,sv2v_dc_113,sv2v_dc_114,sv2v_dc_115,
  sv2v_dc_116,sv2v_dc_117,sv2v_dc_118,sv2v_dc_119,sv2v_dc_120,sv2v_dc_121,sv2v_dc_122,
  sv2v_dc_123,sv2v_dc_124,sv2v_dc_125,sv2v_dc_126,sv2v_dc_127;
  assign { o, sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36, sv2v_dc_37, sv2v_dc_38, sv2v_dc_39, sv2v_dc_40, sv2v_dc_41, sv2v_dc_42, sv2v_dc_43, sv2v_dc_44, sv2v_dc_45, sv2v_dc_46, sv2v_dc_47, sv2v_dc_48, sv2v_dc_49, sv2v_dc_50, sv2v_dc_51, sv2v_dc_52, sv2v_dc_53, sv2v_dc_54, sv2v_dc_55, sv2v_dc_56, sv2v_dc_57, sv2v_dc_58, sv2v_dc_59, sv2v_dc_60, sv2v_dc_61, sv2v_dc_62, sv2v_dc_63, sv2v_dc_64, sv2v_dc_65, sv2v_dc_66, sv2v_dc_67, sv2v_dc_68, sv2v_dc_69, sv2v_dc_70, sv2v_dc_71, sv2v_dc_72, sv2v_dc_73, sv2v_dc_74, sv2v_dc_75, sv2v_dc_76, sv2v_dc_77, sv2v_dc_78, sv2v_dc_79, sv2v_dc_80, sv2v_dc_81, sv2v_dc_82, sv2v_dc_83, sv2v_dc_84, sv2v_dc_85, sv2v_dc_86, sv2v_dc_87, sv2v_dc_88, sv2v_dc_89, sv2v_dc_90, sv2v_dc_91, sv2v_dc_92, sv2v_dc_93, sv2v_dc_94, sv2v_dc_95, sv2v_dc_96, sv2v_dc_97, sv2v_dc_98, sv2v_dc_99, sv2v_dc_100, sv2v_dc_101, sv2v_dc_102, sv2v_dc_103, sv2v_dc_104, sv2v_dc_105, sv2v_dc_106, sv2v_dc_107, sv2v_dc_108, sv2v_dc_109, sv2v_dc_110, sv2v_dc_111, sv2v_dc_112, sv2v_dc_113, sv2v_dc_114, sv2v_dc_115, sv2v_dc_116, sv2v_dc_117, sv2v_dc_118, sv2v_dc_119, sv2v_dc_120, sv2v_dc_121, sv2v_dc_122, sv2v_dc_123, sv2v_dc_124, sv2v_dc_125, sv2v_dc_126, sv2v_dc_127 } = { data_i, data_i[127:1] } << rot_i;

endmodule



module bsg_expand_bitmask_00000004_00000002
(
  i,
  o
);

  input [3:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire o_7_,o_5_,o_3_,o_1_;
  assign o_7_ = i[3];
  assign o[6] = o_7_;
  assign o[7] = o_7_;
  assign o_5_ = i[2];
  assign o[4] = o_5_;
  assign o[5] = o_5_;
  assign o_3_ = i[1];
  assign o[2] = o_3_;
  assign o[3] = o_3_;
  assign o_1_ = i[0];
  assign o[0] = o_1_;
  assign o[1] = o_1_;

endmodule



module bsg_rotate_left_00000008
(
  data_i,
  rot_i,
  o
);

  input [7:0] data_i;
  input [2:0] rot_i;
  output [7:0] o;
  wire [7:0] o;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7;
  assign { o, sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7 } = { data_i, data_i[7:1] } << rot_i;

endmodule



module bsg_rotate_right_00000200
(
  data_i,
  rot_i,
  o
);

  input [511:0] data_i;
  input [8:0] rot_i;
  output [511:0] o;
  wire [511:0] o;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,
  sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,
  sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,sv2v_dc_21,sv2v_dc_22,
  sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,sv2v_dc_27,sv2v_dc_28,sv2v_dc_29,
  sv2v_dc_30,sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,sv2v_dc_34,sv2v_dc_35,sv2v_dc_36,sv2v_dc_37,
  sv2v_dc_38,sv2v_dc_39,sv2v_dc_40,sv2v_dc_41,sv2v_dc_42,sv2v_dc_43,sv2v_dc_44,
  sv2v_dc_45,sv2v_dc_46,sv2v_dc_47,sv2v_dc_48,sv2v_dc_49,sv2v_dc_50,sv2v_dc_51,
  sv2v_dc_52,sv2v_dc_53,sv2v_dc_54,sv2v_dc_55,sv2v_dc_56,sv2v_dc_57,sv2v_dc_58,sv2v_dc_59,
  sv2v_dc_60,sv2v_dc_61,sv2v_dc_62,sv2v_dc_63,sv2v_dc_64,sv2v_dc_65,sv2v_dc_66,
  sv2v_dc_67,sv2v_dc_68,sv2v_dc_69,sv2v_dc_70,sv2v_dc_71,sv2v_dc_72,sv2v_dc_73,
  sv2v_dc_74,sv2v_dc_75,sv2v_dc_76,sv2v_dc_77,sv2v_dc_78,sv2v_dc_79,sv2v_dc_80,
  sv2v_dc_81,sv2v_dc_82,sv2v_dc_83,sv2v_dc_84,sv2v_dc_85,sv2v_dc_86,sv2v_dc_87,sv2v_dc_88,
  sv2v_dc_89,sv2v_dc_90,sv2v_dc_91,sv2v_dc_92,sv2v_dc_93,sv2v_dc_94,sv2v_dc_95,
  sv2v_dc_96,sv2v_dc_97,sv2v_dc_98,sv2v_dc_99,sv2v_dc_100,sv2v_dc_101,sv2v_dc_102,
  sv2v_dc_103,sv2v_dc_104,sv2v_dc_105,sv2v_dc_106,sv2v_dc_107,sv2v_dc_108,sv2v_dc_109,
  sv2v_dc_110,sv2v_dc_111,sv2v_dc_112,sv2v_dc_113,sv2v_dc_114,sv2v_dc_115,
  sv2v_dc_116,sv2v_dc_117,sv2v_dc_118,sv2v_dc_119,sv2v_dc_120,sv2v_dc_121,sv2v_dc_122,
  sv2v_dc_123,sv2v_dc_124,sv2v_dc_125,sv2v_dc_126,sv2v_dc_127,sv2v_dc_128,sv2v_dc_129,
  sv2v_dc_130,sv2v_dc_131,sv2v_dc_132,sv2v_dc_133,sv2v_dc_134,sv2v_dc_135,
  sv2v_dc_136,sv2v_dc_137,sv2v_dc_138,sv2v_dc_139,sv2v_dc_140,sv2v_dc_141,sv2v_dc_142,
  sv2v_dc_143,sv2v_dc_144,sv2v_dc_145,sv2v_dc_146,sv2v_dc_147,sv2v_dc_148,sv2v_dc_149,
  sv2v_dc_150,sv2v_dc_151,sv2v_dc_152,sv2v_dc_153,sv2v_dc_154,sv2v_dc_155,
  sv2v_dc_156,sv2v_dc_157,sv2v_dc_158,sv2v_dc_159,sv2v_dc_160,sv2v_dc_161,sv2v_dc_162,
  sv2v_dc_163,sv2v_dc_164,sv2v_dc_165,sv2v_dc_166,sv2v_dc_167,sv2v_dc_168,sv2v_dc_169,
  sv2v_dc_170,sv2v_dc_171,sv2v_dc_172,sv2v_dc_173,sv2v_dc_174,sv2v_dc_175,
  sv2v_dc_176,sv2v_dc_177,sv2v_dc_178,sv2v_dc_179,sv2v_dc_180,sv2v_dc_181,sv2v_dc_182,
  sv2v_dc_183,sv2v_dc_184,sv2v_dc_185,sv2v_dc_186,sv2v_dc_187,sv2v_dc_188,sv2v_dc_189,
  sv2v_dc_190,sv2v_dc_191,sv2v_dc_192,sv2v_dc_193,sv2v_dc_194,sv2v_dc_195,
  sv2v_dc_196,sv2v_dc_197,sv2v_dc_198,sv2v_dc_199,sv2v_dc_200,sv2v_dc_201,sv2v_dc_202,
  sv2v_dc_203,sv2v_dc_204,sv2v_dc_205,sv2v_dc_206,sv2v_dc_207,sv2v_dc_208,sv2v_dc_209,
  sv2v_dc_210,sv2v_dc_211,sv2v_dc_212,sv2v_dc_213,sv2v_dc_214,sv2v_dc_215,
  sv2v_dc_216,sv2v_dc_217,sv2v_dc_218,sv2v_dc_219,sv2v_dc_220,sv2v_dc_221,sv2v_dc_222,
  sv2v_dc_223,sv2v_dc_224,sv2v_dc_225,sv2v_dc_226,sv2v_dc_227,sv2v_dc_228,sv2v_dc_229,
  sv2v_dc_230,sv2v_dc_231,sv2v_dc_232,sv2v_dc_233,sv2v_dc_234,sv2v_dc_235,
  sv2v_dc_236,sv2v_dc_237,sv2v_dc_238,sv2v_dc_239,sv2v_dc_240,sv2v_dc_241,sv2v_dc_242,
  sv2v_dc_243,sv2v_dc_244,sv2v_dc_245,sv2v_dc_246,sv2v_dc_247,sv2v_dc_248,sv2v_dc_249,
  sv2v_dc_250,sv2v_dc_251,sv2v_dc_252,sv2v_dc_253,sv2v_dc_254,sv2v_dc_255,
  sv2v_dc_256,sv2v_dc_257,sv2v_dc_258,sv2v_dc_259,sv2v_dc_260,sv2v_dc_261,sv2v_dc_262,
  sv2v_dc_263,sv2v_dc_264,sv2v_dc_265,sv2v_dc_266,sv2v_dc_267,sv2v_dc_268,sv2v_dc_269,
  sv2v_dc_270,sv2v_dc_271,sv2v_dc_272,sv2v_dc_273,sv2v_dc_274,sv2v_dc_275,
  sv2v_dc_276,sv2v_dc_277,sv2v_dc_278,sv2v_dc_279,sv2v_dc_280,sv2v_dc_281,sv2v_dc_282,
  sv2v_dc_283,sv2v_dc_284,sv2v_dc_285,sv2v_dc_286,sv2v_dc_287,sv2v_dc_288,sv2v_dc_289,
  sv2v_dc_290,sv2v_dc_291,sv2v_dc_292,sv2v_dc_293,sv2v_dc_294,sv2v_dc_295,
  sv2v_dc_296,sv2v_dc_297,sv2v_dc_298,sv2v_dc_299,sv2v_dc_300,sv2v_dc_301,sv2v_dc_302,
  sv2v_dc_303,sv2v_dc_304,sv2v_dc_305,sv2v_dc_306,sv2v_dc_307,sv2v_dc_308,sv2v_dc_309,
  sv2v_dc_310,sv2v_dc_311,sv2v_dc_312,sv2v_dc_313,sv2v_dc_314,sv2v_dc_315,
  sv2v_dc_316,sv2v_dc_317,sv2v_dc_318,sv2v_dc_319,sv2v_dc_320,sv2v_dc_321,sv2v_dc_322,
  sv2v_dc_323,sv2v_dc_324,sv2v_dc_325,sv2v_dc_326,sv2v_dc_327,sv2v_dc_328,sv2v_dc_329,
  sv2v_dc_330,sv2v_dc_331,sv2v_dc_332,sv2v_dc_333,sv2v_dc_334,sv2v_dc_335,
  sv2v_dc_336,sv2v_dc_337,sv2v_dc_338,sv2v_dc_339,sv2v_dc_340,sv2v_dc_341,sv2v_dc_342,
  sv2v_dc_343,sv2v_dc_344,sv2v_dc_345,sv2v_dc_346,sv2v_dc_347,sv2v_dc_348,sv2v_dc_349,
  sv2v_dc_350,sv2v_dc_351,sv2v_dc_352,sv2v_dc_353,sv2v_dc_354,sv2v_dc_355,
  sv2v_dc_356,sv2v_dc_357,sv2v_dc_358,sv2v_dc_359,sv2v_dc_360,sv2v_dc_361,sv2v_dc_362,
  sv2v_dc_363,sv2v_dc_364,sv2v_dc_365,sv2v_dc_366,sv2v_dc_367,sv2v_dc_368,sv2v_dc_369,
  sv2v_dc_370,sv2v_dc_371,sv2v_dc_372,sv2v_dc_373,sv2v_dc_374,sv2v_dc_375,
  sv2v_dc_376,sv2v_dc_377,sv2v_dc_378,sv2v_dc_379,sv2v_dc_380,sv2v_dc_381,sv2v_dc_382,
  sv2v_dc_383,sv2v_dc_384,sv2v_dc_385,sv2v_dc_386,sv2v_dc_387,sv2v_dc_388,sv2v_dc_389,
  sv2v_dc_390,sv2v_dc_391,sv2v_dc_392,sv2v_dc_393,sv2v_dc_394,sv2v_dc_395,
  sv2v_dc_396,sv2v_dc_397,sv2v_dc_398,sv2v_dc_399,sv2v_dc_400,sv2v_dc_401,sv2v_dc_402,
  sv2v_dc_403,sv2v_dc_404,sv2v_dc_405,sv2v_dc_406,sv2v_dc_407,sv2v_dc_408,sv2v_dc_409,
  sv2v_dc_410,sv2v_dc_411,sv2v_dc_412,sv2v_dc_413,sv2v_dc_414,sv2v_dc_415,
  sv2v_dc_416,sv2v_dc_417,sv2v_dc_418,sv2v_dc_419,sv2v_dc_420,sv2v_dc_421,sv2v_dc_422,
  sv2v_dc_423,sv2v_dc_424,sv2v_dc_425,sv2v_dc_426,sv2v_dc_427,sv2v_dc_428,sv2v_dc_429,
  sv2v_dc_430,sv2v_dc_431,sv2v_dc_432,sv2v_dc_433,sv2v_dc_434,sv2v_dc_435,
  sv2v_dc_436,sv2v_dc_437,sv2v_dc_438,sv2v_dc_439,sv2v_dc_440,sv2v_dc_441,sv2v_dc_442,
  sv2v_dc_443,sv2v_dc_444,sv2v_dc_445,sv2v_dc_446,sv2v_dc_447,sv2v_dc_448,sv2v_dc_449,
  sv2v_dc_450,sv2v_dc_451,sv2v_dc_452,sv2v_dc_453,sv2v_dc_454,sv2v_dc_455,
  sv2v_dc_456,sv2v_dc_457,sv2v_dc_458,sv2v_dc_459,sv2v_dc_460,sv2v_dc_461,sv2v_dc_462,
  sv2v_dc_463,sv2v_dc_464,sv2v_dc_465,sv2v_dc_466,sv2v_dc_467,sv2v_dc_468,sv2v_dc_469,
  sv2v_dc_470,sv2v_dc_471,sv2v_dc_472,sv2v_dc_473,sv2v_dc_474,sv2v_dc_475,
  sv2v_dc_476,sv2v_dc_477,sv2v_dc_478,sv2v_dc_479,sv2v_dc_480,sv2v_dc_481,sv2v_dc_482,
  sv2v_dc_483,sv2v_dc_484,sv2v_dc_485,sv2v_dc_486,sv2v_dc_487,sv2v_dc_488,sv2v_dc_489,
  sv2v_dc_490,sv2v_dc_491,sv2v_dc_492,sv2v_dc_493,sv2v_dc_494,sv2v_dc_495,
  sv2v_dc_496,sv2v_dc_497,sv2v_dc_498,sv2v_dc_499,sv2v_dc_500,sv2v_dc_501,sv2v_dc_502,
  sv2v_dc_503,sv2v_dc_504,sv2v_dc_505,sv2v_dc_506,sv2v_dc_507,sv2v_dc_508,sv2v_dc_509,
  sv2v_dc_510,sv2v_dc_511;
  assign { sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36, sv2v_dc_37, sv2v_dc_38, sv2v_dc_39, sv2v_dc_40, sv2v_dc_41, sv2v_dc_42, sv2v_dc_43, sv2v_dc_44, sv2v_dc_45, sv2v_dc_46, sv2v_dc_47, sv2v_dc_48, sv2v_dc_49, sv2v_dc_50, sv2v_dc_51, sv2v_dc_52, sv2v_dc_53, sv2v_dc_54, sv2v_dc_55, sv2v_dc_56, sv2v_dc_57, sv2v_dc_58, sv2v_dc_59, sv2v_dc_60, sv2v_dc_61, sv2v_dc_62, sv2v_dc_63, sv2v_dc_64, sv2v_dc_65, sv2v_dc_66, sv2v_dc_67, sv2v_dc_68, sv2v_dc_69, sv2v_dc_70, sv2v_dc_71, sv2v_dc_72, sv2v_dc_73, sv2v_dc_74, sv2v_dc_75, sv2v_dc_76, sv2v_dc_77, sv2v_dc_78, sv2v_dc_79, sv2v_dc_80, sv2v_dc_81, sv2v_dc_82, sv2v_dc_83, sv2v_dc_84, sv2v_dc_85, sv2v_dc_86, sv2v_dc_87, sv2v_dc_88, sv2v_dc_89, sv2v_dc_90, sv2v_dc_91, sv2v_dc_92, sv2v_dc_93, sv2v_dc_94, sv2v_dc_95, sv2v_dc_96, sv2v_dc_97, sv2v_dc_98, sv2v_dc_99, sv2v_dc_100, sv2v_dc_101, sv2v_dc_102, sv2v_dc_103, sv2v_dc_104, sv2v_dc_105, sv2v_dc_106, sv2v_dc_107, sv2v_dc_108, sv2v_dc_109, sv2v_dc_110, sv2v_dc_111, sv2v_dc_112, sv2v_dc_113, sv2v_dc_114, sv2v_dc_115, sv2v_dc_116, sv2v_dc_117, sv2v_dc_118, sv2v_dc_119, sv2v_dc_120, sv2v_dc_121, sv2v_dc_122, sv2v_dc_123, sv2v_dc_124, sv2v_dc_125, sv2v_dc_126, sv2v_dc_127, sv2v_dc_128, sv2v_dc_129, sv2v_dc_130, sv2v_dc_131, sv2v_dc_132, sv2v_dc_133, sv2v_dc_134, sv2v_dc_135, sv2v_dc_136, sv2v_dc_137, sv2v_dc_138, sv2v_dc_139, sv2v_dc_140, sv2v_dc_141, sv2v_dc_142, sv2v_dc_143, sv2v_dc_144, sv2v_dc_145, sv2v_dc_146, sv2v_dc_147, sv2v_dc_148, sv2v_dc_149, sv2v_dc_150, sv2v_dc_151, sv2v_dc_152, sv2v_dc_153, sv2v_dc_154, sv2v_dc_155, sv2v_dc_156, sv2v_dc_157, sv2v_dc_158, sv2v_dc_159, sv2v_dc_160, sv2v_dc_161, sv2v_dc_162, sv2v_dc_163, sv2v_dc_164, sv2v_dc_165, sv2v_dc_166, sv2v_dc_167, sv2v_dc_168, sv2v_dc_169, sv2v_dc_170, sv2v_dc_171, sv2v_dc_172, sv2v_dc_173, sv2v_dc_174, sv2v_dc_175, sv2v_dc_176, sv2v_dc_177, sv2v_dc_178, sv2v_dc_179, sv2v_dc_180, sv2v_dc_181, sv2v_dc_182, sv2v_dc_183, sv2v_dc_184, sv2v_dc_185, sv2v_dc_186, sv2v_dc_187, sv2v_dc_188, sv2v_dc_189, sv2v_dc_190, sv2v_dc_191, sv2v_dc_192, sv2v_dc_193, sv2v_dc_194, sv2v_dc_195, sv2v_dc_196, sv2v_dc_197, sv2v_dc_198, sv2v_dc_199, sv2v_dc_200, sv2v_dc_201, sv2v_dc_202, sv2v_dc_203, sv2v_dc_204, sv2v_dc_205, sv2v_dc_206, sv2v_dc_207, sv2v_dc_208, sv2v_dc_209, sv2v_dc_210, sv2v_dc_211, sv2v_dc_212, sv2v_dc_213, sv2v_dc_214, sv2v_dc_215, sv2v_dc_216, sv2v_dc_217, sv2v_dc_218, sv2v_dc_219, sv2v_dc_220, sv2v_dc_221, sv2v_dc_222, sv2v_dc_223, sv2v_dc_224, sv2v_dc_225, sv2v_dc_226, sv2v_dc_227, sv2v_dc_228, sv2v_dc_229, sv2v_dc_230, sv2v_dc_231, sv2v_dc_232, sv2v_dc_233, sv2v_dc_234, sv2v_dc_235, sv2v_dc_236, sv2v_dc_237, sv2v_dc_238, sv2v_dc_239, sv2v_dc_240, sv2v_dc_241, sv2v_dc_242, sv2v_dc_243, sv2v_dc_244, sv2v_dc_245, sv2v_dc_246, sv2v_dc_247, sv2v_dc_248, sv2v_dc_249, sv2v_dc_250, sv2v_dc_251, sv2v_dc_252, sv2v_dc_253, sv2v_dc_254, sv2v_dc_255, sv2v_dc_256, sv2v_dc_257, sv2v_dc_258, sv2v_dc_259, sv2v_dc_260, sv2v_dc_261, sv2v_dc_262, sv2v_dc_263, sv2v_dc_264, sv2v_dc_265, sv2v_dc_266, sv2v_dc_267, sv2v_dc_268, sv2v_dc_269, sv2v_dc_270, sv2v_dc_271, sv2v_dc_272, sv2v_dc_273, sv2v_dc_274, sv2v_dc_275, sv2v_dc_276, sv2v_dc_277, sv2v_dc_278, sv2v_dc_279, sv2v_dc_280, sv2v_dc_281, sv2v_dc_282, sv2v_dc_283, sv2v_dc_284, sv2v_dc_285, sv2v_dc_286, sv2v_dc_287, sv2v_dc_288, sv2v_dc_289, sv2v_dc_290, sv2v_dc_291, sv2v_dc_292, sv2v_dc_293, sv2v_dc_294, sv2v_dc_295, sv2v_dc_296, sv2v_dc_297, sv2v_dc_298, sv2v_dc_299, sv2v_dc_300, sv2v_dc_301, sv2v_dc_302, sv2v_dc_303, sv2v_dc_304, sv2v_dc_305, sv2v_dc_306, sv2v_dc_307, sv2v_dc_308, sv2v_dc_309, sv2v_dc_310, sv2v_dc_311, sv2v_dc_312, sv2v_dc_313, sv2v_dc_314, sv2v_dc_315, sv2v_dc_316, sv2v_dc_317, sv2v_dc_318, sv2v_dc_319, sv2v_dc_320, sv2v_dc_321, sv2v_dc_322, sv2v_dc_323, sv2v_dc_324, sv2v_dc_325, sv2v_dc_326, sv2v_dc_327, sv2v_dc_328, sv2v_dc_329, sv2v_dc_330, sv2v_dc_331, sv2v_dc_332, sv2v_dc_333, sv2v_dc_334, sv2v_dc_335, sv2v_dc_336, sv2v_dc_337, sv2v_dc_338, sv2v_dc_339, sv2v_dc_340, sv2v_dc_341, sv2v_dc_342, sv2v_dc_343, sv2v_dc_344, sv2v_dc_345, sv2v_dc_346, sv2v_dc_347, sv2v_dc_348, sv2v_dc_349, sv2v_dc_350, sv2v_dc_351, sv2v_dc_352, sv2v_dc_353, sv2v_dc_354, sv2v_dc_355, sv2v_dc_356, sv2v_dc_357, sv2v_dc_358, sv2v_dc_359, sv2v_dc_360, sv2v_dc_361, sv2v_dc_362, sv2v_dc_363, sv2v_dc_364, sv2v_dc_365, sv2v_dc_366, sv2v_dc_367, sv2v_dc_368, sv2v_dc_369, sv2v_dc_370, sv2v_dc_371, sv2v_dc_372, sv2v_dc_373, sv2v_dc_374, sv2v_dc_375, sv2v_dc_376, sv2v_dc_377, sv2v_dc_378, sv2v_dc_379, sv2v_dc_380, sv2v_dc_381, sv2v_dc_382, sv2v_dc_383, sv2v_dc_384, sv2v_dc_385, sv2v_dc_386, sv2v_dc_387, sv2v_dc_388, sv2v_dc_389, sv2v_dc_390, sv2v_dc_391, sv2v_dc_392, sv2v_dc_393, sv2v_dc_394, sv2v_dc_395, sv2v_dc_396, sv2v_dc_397, sv2v_dc_398, sv2v_dc_399, sv2v_dc_400, sv2v_dc_401, sv2v_dc_402, sv2v_dc_403, sv2v_dc_404, sv2v_dc_405, sv2v_dc_406, sv2v_dc_407, sv2v_dc_408, sv2v_dc_409, sv2v_dc_410, sv2v_dc_411, sv2v_dc_412, sv2v_dc_413, sv2v_dc_414, sv2v_dc_415, sv2v_dc_416, sv2v_dc_417, sv2v_dc_418, sv2v_dc_419, sv2v_dc_420, sv2v_dc_421, sv2v_dc_422, sv2v_dc_423, sv2v_dc_424, sv2v_dc_425, sv2v_dc_426, sv2v_dc_427, sv2v_dc_428, sv2v_dc_429, sv2v_dc_430, sv2v_dc_431, sv2v_dc_432, sv2v_dc_433, sv2v_dc_434, sv2v_dc_435, sv2v_dc_436, sv2v_dc_437, sv2v_dc_438, sv2v_dc_439, sv2v_dc_440, sv2v_dc_441, sv2v_dc_442, sv2v_dc_443, sv2v_dc_444, sv2v_dc_445, sv2v_dc_446, sv2v_dc_447, sv2v_dc_448, sv2v_dc_449, sv2v_dc_450, sv2v_dc_451, sv2v_dc_452, sv2v_dc_453, sv2v_dc_454, sv2v_dc_455, sv2v_dc_456, sv2v_dc_457, sv2v_dc_458, sv2v_dc_459, sv2v_dc_460, sv2v_dc_461, sv2v_dc_462, sv2v_dc_463, sv2v_dc_464, sv2v_dc_465, sv2v_dc_466, sv2v_dc_467, sv2v_dc_468, sv2v_dc_469, sv2v_dc_470, sv2v_dc_471, sv2v_dc_472, sv2v_dc_473, sv2v_dc_474, sv2v_dc_475, sv2v_dc_476, sv2v_dc_477, sv2v_dc_478, sv2v_dc_479, sv2v_dc_480, sv2v_dc_481, sv2v_dc_482, sv2v_dc_483, sv2v_dc_484, sv2v_dc_485, sv2v_dc_486, sv2v_dc_487, sv2v_dc_488, sv2v_dc_489, sv2v_dc_490, sv2v_dc_491, sv2v_dc_492, sv2v_dc_493, sv2v_dc_494, sv2v_dc_495, sv2v_dc_496, sv2v_dc_497, sv2v_dc_498, sv2v_dc_499, sv2v_dc_500, sv2v_dc_501, sv2v_dc_502, sv2v_dc_503, sv2v_dc_504, sv2v_dc_505, sv2v_dc_506, sv2v_dc_507, sv2v_dc_508, sv2v_dc_509, sv2v_dc_510, sv2v_dc_511, o } = { data_i[510:0], data_i } >> rot_i;

endmodule



module bp_fe_icache_00
(
  clk_i,
  reset_i,
  cfg_bus_i,
  icache_pkt_i,
  v_i,
  force_i,
  yumi_o,
  tl_flush_i,
  ptag_i,
  ptag_v_i,
  ptag_uncached_i,
  ptag_nonidem_i,
  ptag_dram_i,
  tv_flush_i,
  tv_we_o,
  data_o,
  hit_v_o,
  miss_v_o,
  fence_v_o,
  yumi_i,
  cache_req_o,
  cache_req_v_o,
  cache_req_yumi_i,
  cache_req_lock_i,
  cache_req_metadata_o,
  cache_req_metadata_v_o,
  cache_req_id_i,
  cache_req_critical_i,
  cache_req_last_i,
  cache_req_credits_full_i,
  cache_req_credits_empty_i,
  data_mem_pkt_v_i,
  data_mem_pkt_i,
  data_mem_pkt_yumi_o,
  data_mem_o,
  tag_mem_pkt_v_i,
  tag_mem_pkt_i,
  tag_mem_pkt_yumi_o,
  tag_mem_o,
  stat_mem_pkt_v_i,
  stat_mem_pkt_i,
  stat_mem_pkt_yumi_o,
  stat_mem_o
);

  input [60:0] cfg_bus_i;
  input [71:0] icache_pkt_i;
  input [27:0] ptag_i;
  output [63:0] data_o;
  output [116:0] cache_req_o;
  output [3:0] cache_req_metadata_o;
  input [0:0] cache_req_id_i;
  input [142:0] data_mem_pkt_i;
  output [511:0] data_mem_o;
  input [34:0] tag_mem_pkt_i;
  output [22:0] tag_mem_o;
  input [10:0] stat_mem_pkt_i;
  output [14:0] stat_mem_o;
  input clk_i;
  input reset_i;
  input v_i;
  input force_i;
  input tl_flush_i;
  input ptag_v_i;
  input ptag_uncached_i;
  input ptag_nonidem_i;
  input ptag_dram_i;
  input tv_flush_i;
  input yumi_i;
  input cache_req_yumi_i;
  input cache_req_lock_i;
  input cache_req_critical_i;
  input cache_req_last_i;
  input cache_req_credits_full_i;
  input cache_req_credits_empty_i;
  input data_mem_pkt_v_i;
  input tag_mem_pkt_v_i;
  input stat_mem_pkt_v_i;
  output yumi_o;
  output tv_we_o;
  output hit_v_o;
  output miss_v_o;
  output fence_v_o;
  output cache_req_v_o;
  output cache_req_metadata_v_o;
  output data_mem_pkt_yumi_o;
  output tag_mem_pkt_yumi_o;
  output stat_mem_pkt_yumi_o;
  wire [63:0] data_o,ld_data_way_picked;
  wire [116:0] cache_req_o;
  wire [3:0] cache_req_metadata_o;
  wire [511:0] data_mem_o,data_mem_data_lo,ld_data_tv_n,ld_data_tv_r;
  wire [22:0] tag_mem_o;
  wire [14:0] stat_mem_o;
  wire yumi_o,tv_we_o,hit_v_o,miss_v_o,fence_v_o,cache_req_v_o,cache_req_metadata_v_o,
  data_mem_pkt_yumi_o,tag_mem_pkt_yumi_o,stat_mem_pkt_yumi_o,N0,N1,N2,N3,N4,N5,N6,
  N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,
  N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,
  N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,
  critical_recv,complete_recv,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  decode_lo_fetch_op_,decode_lo_inval_op_,tl_we,tag_mem_v_li,tag_mem_w_li,v_tl_r,N99,N100,
  N101,N102,_0_net_,decode_tl_r_fetch_op_,decode_tl_r_inval_op_,spec_tl_r,N103,
  \tag_comp_tl_0_.tag_match_tl ,N104,N105,\tag_comp_tl_1_.tag_match_tl ,N106,N107,
  \tag_comp_tl_2_.tag_match_tl ,N108,N109,\tag_comp_tl_3_.tag_match_tl ,N110,N111,
  \tag_comp_tl_4_.tag_match_tl ,N112,N113,\tag_comp_tl_5_.tag_match_tl ,N114,N115,
  \tag_comp_tl_6_.tag_match_tl ,N116,N117,\tag_comp_tl_7_.tag_match_tl ,N118,
  fetch_uncached_tl,spec_tl,v_tv_r,N119,_3_net_,decode_tv_n_fetch_op_,
  decode_tv_n_inval_op_,spec_tv_n,uncached_tv_n,snoop_decode_fetch_op_,snoop_decode_inval_op_,
  snoop_spec,snoop_uncached,_6_net_,snoop_tv_r,N120,N121,_9_net_,_10_net__7_,_10_net__6_,
  _10_net__5_,_10_net__4_,_10_net__3_,_10_net__2_,_10_net__1_,_10_net__0_,
  invalid_exist_tv,N122,stat_mem_v_li,stat_mem_w_li,stat_mem_mask_li_lru__6_,
  stat_mem_mask_li_lru__5_,stat_mem_mask_li_lru__4_,stat_mem_mask_li_lru__3_,
  stat_mem_mask_li_lru__2_,stat_mem_mask_li_lru__1_,stat_mem_mask_li_lru__0_,
  stat_mem_data_li_lru__6_,stat_mem_data_li_lru__5_,stat_mem_data_li_lru__4_,stat_mem_data_li_lru__3_,
  stat_mem_data_li_lru__2_,stat_mem_data_li_lru__1_,stat_mem_data_li_lru__0_,
  cached_req,uncached_req,inval_req,N123,N124,N125,N126,N127,metadata_hit_r,N128,N129,N130,
  N131,N132,N133,N134,do_recover,N135,tag_mem_bypass,tag_mem_fast_read,
  tag_mem_slow_read,tag_mem_slow_write,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,
  N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,
  N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,
  N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
  N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,
  N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,
  N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,
  N242,N243,N244,N245,N246,N247,N248,N249,N250,data_mem_bypass,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,
  N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,
  N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,
  stat_mem_fast_read,stat_mem_fast_write,stat_mem_slow_write,N332,N333,N334,N335,N336,N337,N338,
  N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,
  N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,
  N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,
  N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,
  N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,
  N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,
  N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,
  N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,
  N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,
  N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,
  N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,
  N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,
  N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,
  N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,
  N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,
  N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,
  N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,
  N611;
  wire [1:0] state_r,state_n;
  wire [183:0] tag_mem_data_li,tag_mem_w_mask_li,tag_mem_data_lo;
  wire [5:0] tag_mem_addr_li,stat_mem_addr_li;
  wire [71:0] data_mem_addr_li;
  wire [7:0] data_mem_v_li,hit_v_tl,bank_sel_one_hot_tl,bank_sel_one_hot_tv_n,way_v_tv_n,
  hit_v_tv_n,bank_sel_one_hot_tv_r,way_v_tv_r,hit_v_tv_r,ld_data_way_select_tv,
  tag_mem_way_one_hot,vaddr_bank_dec,data_mem_bypass_select,
  data_mem_pkt_fill_mask_expanded,data_mem_write_bank_mask,data_mem_slow_read,data_mem_slow_write,
  data_mem_fast_read,pseudo_hit;
  wire [11:0] paddr_tl;
  wire [26:0] vaddr_vtag_tl;
  wire [39:0] paddr_tv_n;
  wire [2:0] invalid_way_tv,lru_way_li,lru_encode,hit_index_tv,metadata_hit_index_r,
  tag_mem_pkt_way_r,\data_mem_lines_0_.data_mem_pkt_offset ,
  \data_mem_lines_1_.data_mem_pkt_offset ,\data_mem_lines_2_.data_mem_pkt_offset ,
  \data_mem_lines_3_.data_mem_pkt_offset ,\data_mem_lines_4_.data_mem_pkt_offset ,
  \data_mem_lines_5_.data_mem_pkt_offset ,\data_mem_lines_6_.data_mem_pkt_offset ,
  \data_mem_lines_7_.data_mem_pkt_offset ,data_mem_pkt_way_r;
  wire [127:0] data_mem_pkt_fill_data_li;
  wire [6:0] lru_decode_data_lo,lru_decode_mask_lo;
  reg state_r_1_sv2v_reg,state_r_0_sv2v_reg;
  assign state_r[1] = state_r_1_sv2v_reg;
  assign state_r[0] = state_r_0_sv2v_reg;
  assign cache_req_o[0] = 1'b1;
  assign cache_req_o[1] = 1'b1;
  assign cache_req_o[49] = 1'b1;
  assign stat_mem_o[0] = 1'b0;
  assign stat_mem_o[1] = 1'b0;
  assign stat_mem_o[2] = 1'b0;
  assign stat_mem_o[3] = 1'b0;
  assign stat_mem_o[4] = 1'b0;
  assign stat_mem_o[5] = 1'b0;
  assign stat_mem_o[6] = 1'b0;
  assign stat_mem_o[7] = 1'b0;
  assign cache_req_metadata_o[0] = 1'b0;
  assign cache_req_o[2] = 1'b0;
  assign cache_req_o[3] = 1'b0;
  assign cache_req_o[7] = 1'b0;
  assign cache_req_o[51] = 1'b0;
  assign cache_req_o[52] = 1'b0;
  assign cache_req_o[53] = 1'b0;
  assign cache_req_o[54] = 1'b0;
  assign cache_req_o[55] = 1'b0;
  assign cache_req_o[56] = 1'b0;
  assign cache_req_o[57] = 1'b0;
  assign cache_req_o[58] = 1'b0;
  assign cache_req_o[59] = 1'b0;
  assign cache_req_o[60] = 1'b0;
  assign cache_req_o[61] = 1'b0;
  assign cache_req_o[62] = 1'b0;
  assign cache_req_o[63] = 1'b0;
  assign cache_req_o[64] = 1'b0;
  assign cache_req_o[65] = 1'b0;
  assign cache_req_o[66] = 1'b0;
  assign cache_req_o[67] = 1'b0;
  assign cache_req_o[68] = 1'b0;
  assign cache_req_o[69] = 1'b0;
  assign cache_req_o[70] = 1'b0;
  assign cache_req_o[71] = 1'b0;
  assign cache_req_o[72] = 1'b0;
  assign cache_req_o[73] = 1'b0;
  assign cache_req_o[74] = 1'b0;
  assign cache_req_o[75] = 1'b0;
  assign cache_req_o[76] = 1'b0;
  assign cache_req_o[77] = 1'b0;
  assign cache_req_o[78] = 1'b0;
  assign cache_req_o[79] = 1'b0;
  assign cache_req_o[80] = 1'b0;
  assign cache_req_o[81] = 1'b0;
  assign cache_req_o[82] = 1'b0;
  assign cache_req_o[83] = 1'b0;
  assign cache_req_o[84] = 1'b0;
  assign cache_req_o[85] = 1'b0;
  assign cache_req_o[86] = 1'b0;
  assign cache_req_o[87] = 1'b0;
  assign cache_req_o[88] = 1'b0;
  assign cache_req_o[89] = 1'b0;
  assign cache_req_o[90] = 1'b0;
  assign cache_req_o[91] = 1'b0;
  assign cache_req_o[92] = 1'b0;
  assign cache_req_o[93] = 1'b0;
  assign cache_req_o[94] = 1'b0;
  assign cache_req_o[95] = 1'b0;
  assign cache_req_o[96] = 1'b0;
  assign cache_req_o[97] = 1'b0;
  assign cache_req_o[98] = 1'b0;
  assign cache_req_o[99] = 1'b0;
  assign cache_req_o[100] = 1'b0;
  assign cache_req_o[101] = 1'b0;
  assign cache_req_o[102] = 1'b0;
  assign cache_req_o[103] = 1'b0;
  assign cache_req_o[104] = 1'b0;
  assign cache_req_o[105] = 1'b0;
  assign cache_req_o[106] = 1'b0;
  assign cache_req_o[107] = 1'b0;
  assign cache_req_o[108] = 1'b0;
  assign cache_req_o[109] = 1'b0;
  assign cache_req_o[110] = 1'b0;
  assign cache_req_o[111] = 1'b0;
  assign cache_req_o[112] = 1'b0;
  assign cache_req_o[113] = 1'b0;
  assign cache_req_o[114] = 1'b0;
  assign cache_req_o[116] = 1'b0;
  assign N66 = icache_pkt_i[31] | icache_pkt_i[32];
  assign N67 = icache_pkt_i[30] | N66;
  assign N68 = icache_pkt_i[29] | N67;
  assign N69 = icache_pkt_i[28] | N68;
  assign N70 = icache_pkt_i[27] | N69;
  assign N71 = icache_pkt_i[26] | N70;
  assign N72 = icache_pkt_i[25] | N71;
  assign N73 = icache_pkt_i[24] | N72;
  assign N74 = icache_pkt_i[23] | N73;
  assign N75 = icache_pkt_i[22] | N74;
  assign N76 = icache_pkt_i[21] | N75;
  assign N77 = icache_pkt_i[20] | N76;
  assign N78 = icache_pkt_i[19] | N77;
  assign N79 = icache_pkt_i[18] | N78;
  assign N80 = icache_pkt_i[17] | N79;
  assign N81 = icache_pkt_i[16] | N80;
  assign N82 = icache_pkt_i[15] | N81;
  assign N83 = icache_pkt_i[14] | N82;
  assign N84 = icache_pkt_i[13] | N83;
  assign N85 = icache_pkt_i[12] | N84;
  assign N86 = icache_pkt_i[11] | N85;
  assign N87 = icache_pkt_i[10] | N86;
  assign N88 = icache_pkt_i[9] | N87;
  assign N89 = icache_pkt_i[8] | N88;
  assign N90 = icache_pkt_i[7] | N89;
  assign N91 = icache_pkt_i[6] | N90;
  assign N92 = icache_pkt_i[5] | N91;
  assign N93 = icache_pkt_i[4] | N92;
  assign N94 = icache_pkt_i[3] | N93;
  assign N95 = icache_pkt_i[2] | N94;
  assign N96 = icache_pkt_i[1] | N95;
  assign decode_lo_fetch_op_ = ~N96;
  assign N97 = ~icache_pkt_i[1];
  assign N98 = N97 | N95;
  assign decode_lo_inval_op_ = ~N98;

  bsg_mem_1rw_sync_mask_write_bit_000000b8_00000040_1
  tag_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(tag_mem_data_li),
    .addr_i(tag_mem_addr_li),
    .v_i(tag_mem_v_li),
    .w_mask_i(tag_mem_w_mask_li),
    .w_i(tag_mem_w_li),
    .data_o(tag_mem_data_lo)
  );


  bsg_mem_1rw_sync_00000040_00000200_1
  \data_mems_0_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_mem_pkt_fill_data_li[63:0]),
    .addr_i(data_mem_addr_li[8:0]),
    .v_i(data_mem_v_li[0]),
    .w_i(data_mem_slow_write[0]),
    .data_o(data_mem_data_lo[63:0])
  );


  bsg_mem_1rw_sync_00000040_00000200_1
  \data_mems_1_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_mem_pkt_fill_data_li[127:64]),
    .addr_i(data_mem_addr_li[17:9]),
    .v_i(data_mem_v_li[1]),
    .w_i(data_mem_slow_write[1]),
    .data_o(data_mem_data_lo[127:64])
  );


  bsg_mem_1rw_sync_00000040_00000200_1
  \data_mems_2_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_mem_pkt_fill_data_li[63:0]),
    .addr_i(data_mem_addr_li[26:18]),
    .v_i(data_mem_v_li[2]),
    .w_i(data_mem_slow_write[2]),
    .data_o(data_mem_data_lo[191:128])
  );


  bsg_mem_1rw_sync_00000040_00000200_1
  \data_mems_3_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_mem_pkt_fill_data_li[127:64]),
    .addr_i(data_mem_addr_li[35:27]),
    .v_i(data_mem_v_li[3]),
    .w_i(data_mem_slow_write[3]),
    .data_o(data_mem_data_lo[255:192])
  );


  bsg_mem_1rw_sync_00000040_00000200_1
  \data_mems_4_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_mem_pkt_fill_data_li[63:0]),
    .addr_i(data_mem_addr_li[44:36]),
    .v_i(data_mem_v_li[4]),
    .w_i(data_mem_slow_write[4]),
    .data_o(data_mem_data_lo[319:256])
  );


  bsg_mem_1rw_sync_00000040_00000200_1
  \data_mems_5_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_mem_pkt_fill_data_li[127:64]),
    .addr_i(data_mem_addr_li[53:45]),
    .v_i(data_mem_v_li[5]),
    .w_i(data_mem_slow_write[5]),
    .data_o(data_mem_data_lo[383:320])
  );


  bsg_mem_1rw_sync_00000040_00000200_1
  \data_mems_6_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_mem_pkt_fill_data_li[63:0]),
    .addr_i(data_mem_addr_li[62:54]),
    .v_i(data_mem_v_li[6]),
    .w_i(data_mem_slow_write[6]),
    .data_o(data_mem_data_lo[447:384])
  );


  bsg_mem_1rw_sync_00000040_00000200_1
  \data_mems_7_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_mem_pkt_fill_data_li[127:64]),
    .addr_i(data_mem_addr_li[71:63]),
    .v_i(data_mem_v_li[7]),
    .w_i(data_mem_slow_write[7]),
    .data_o(data_mem_data_lo[511:448])
  );


  bsg_dff_reset_en_width_p1
  v_tl_reg
  (
    .clk_i(clk_i),
    .reset_i(_0_net_),
    .en_i(tl_we),
    .data_i(yumi_o),
    .data_o(v_tl_r)
  );


  bsg_dff_reset_en_0000002a
  tl_stage_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(tl_we),
    .data_i({ icache_pkt_i[71:33], icache_pkt_i[0:0], decode_lo_fetch_op_, decode_lo_inval_op_ }),
    .data_o({ vaddr_vtag_tl, paddr_tl, spec_tl_r, decode_tl_r_fetch_op_, decode_tl_r_inval_op_ })
  );

  assign N103 = ptag_i[19:0] == tag_mem_data_lo[19:0];
  assign N104 = tag_mem_data_lo[19:0] == ptag_i[19:0];
  assign N105 = ptag_i[19:0] == tag_mem_data_lo[42:23];
  assign N106 = tag_mem_data_lo[42:23] == ptag_i[19:0];
  assign N107 = ptag_i[19:0] == tag_mem_data_lo[65:46];
  assign N108 = tag_mem_data_lo[65:46] == ptag_i[19:0];
  assign N109 = ptag_i[19:0] == tag_mem_data_lo[88:69];
  assign N110 = tag_mem_data_lo[88:69] == ptag_i[19:0];
  assign N111 = ptag_i[19:0] == tag_mem_data_lo[111:92];
  assign N112 = tag_mem_data_lo[111:92] == ptag_i[19:0];
  assign N113 = ptag_i[19:0] == tag_mem_data_lo[134:115];
  assign N114 = tag_mem_data_lo[134:115] == ptag_i[19:0];
  assign N115 = ptag_i[19:0] == tag_mem_data_lo[157:138];
  assign N116 = tag_mem_data_lo[157:138] == ptag_i[19:0];
  assign N117 = ptag_i[19:0] == tag_mem_data_lo[180:161];
  assign N118 = tag_mem_data_lo[180:161] == ptag_i[19:0];

  bsg_decode_00000008
  offset_decode
  (
    .i(paddr_tl[5:3]),
    .o(bank_sel_one_hot_tl)
  );


  bsg_dff_reset_en_width_p1
  v_tv_reg
  (
    .clk_i(clk_i),
    .reset_i(_3_net_),
    .en_i(tv_we_o),
    .data_i(v_tl_r),
    .data_o(v_tv_r)
  );


  bsg_mux_0000021c_2
  hit_mux
  (
    .data_i({ bank_sel_one_hot_tv_r, pseudo_hit, pseudo_hit, data_mem_pkt_fill_data_li, data_mem_pkt_fill_data_li, data_mem_pkt_fill_data_li, data_mem_pkt_fill_data_li, snoop_spec, snoop_uncached, snoop_decode_fetch_op_, snoop_decode_inval_op_, bank_sel_one_hot_tl, N354, N356, N358, N360, N362, N364, N366, N368, hit_v_tl, data_mem_data_lo, spec_tl, fetch_uncached_tl, decode_tl_r_fetch_op_, decode_tl_r_inval_op_ }),
    .sel_i(critical_recv),
    .data_o({ bank_sel_one_hot_tv_n, way_v_tv_n, hit_v_tv_n, ld_data_tv_n, spec_tv_n, uncached_tv_n, decode_tv_n_fetch_op_, decode_tv_n_inval_op_ })
  );


  bsg_dff_reset_en_0000021d
  tv_stage_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(_6_net_),
    .data_i({ ld_data_tv_n, critical_recv, bank_sel_one_hot_tv_n, way_v_tv_n, hit_v_tv_n, spec_tv_n, uncached_tv_n, decode_tv_n_fetch_op_, decode_tv_n_inval_op_ }),
    .data_o({ ld_data_tv_r, snoop_tv_r, bank_sel_one_hot_tv_r, way_v_tv_r, hit_v_tv_r, snoop_spec, snoop_uncached, snoop_decode_fetch_op_, snoop_decode_inval_op_ })
  );


  bsg_dff_en_00000028
  paddr_reg
  (
    .clk_i(clk_i),
    .data_i(paddr_tv_n),
    .en_i(_9_net_),
    .data_o(cache_req_o[47:8])
  );


  bsg_priority_encode_00000008_1
  pe_invalid
  (
    .i({ _10_net__7_, _10_net__6_, _10_net__5_, _10_net__4_, _10_net__3_, _10_net__2_, _10_net__1_, _10_net__0_ }),
    .addr_o(invalid_way_tv),
    .v_o(invalid_exist_tv)
  );


  bsg_encode_one_hot_00000008_1
  hit_index_encoder
  (
    .i(hit_v_tv_r),
    .addr_o(hit_index_tv),
    .v_o(cache_req_o[115])
  );


  bsg_adder_one_hot_00000008
  select_adder
  (
    .a_i(hit_v_tv_r),
    .b_i(bank_sel_one_hot_tv_r),
    .o(ld_data_way_select_tv)
  );


  bsg_mux_one_hot_00000040_00000008
  data_set_select_mux
  (
    .data_i(ld_data_tv_r),
    .sel_one_hot_i(ld_data_way_select_tv),
    .data_o(ld_data_way_picked)
  );


  bsg_mux_00000040_00000001
  data_select_mux
  (
    .data_i(ld_data_way_picked),
    .sel_i(cache_req_o[10]),
    .data_o(data_o)
  );


  bsg_mem_1rw_sync_mask_write_bit_00000007_00000040_1
  stat_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ stat_mem_data_li_lru__6_, stat_mem_data_li_lru__5_, stat_mem_data_li_lru__4_, stat_mem_data_li_lru__3_, stat_mem_data_li_lru__2_, stat_mem_data_li_lru__1_, stat_mem_data_li_lru__0_ }),
    .addr_i(stat_mem_addr_li),
    .v_i(stat_mem_v_li),
    .w_mask_i({ stat_mem_mask_li_lru__6_, stat_mem_mask_li_lru__5_, stat_mem_mask_li_lru__4_, stat_mem_mask_li_lru__3_, stat_mem_mask_li_lru__2_, stat_mem_mask_li_lru__1_, stat_mem_mask_li_lru__0_ }),
    .w_i(stat_mem_w_li),
    .data_o(stat_mem_o[14:8])
  );


  bsg_lru_pseudo_tree_encode_00000008
  lru_encoder
  (
    .lru_i(stat_mem_o[14:8]),
    .way_id_o(lru_encode)
  );


  bsg_dff_reset_width_p1
  cache_req_v_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(cache_req_yumi_i),
    .data_o(cache_req_metadata_v_o)
  );


  bsg_dff_00000004
  hit_reg
  (
    .clk_i(clk_i),
    .data_i({ cache_req_o[115:115], hit_index_tv }),
    .data_o({ metadata_hit_r, metadata_hit_index_r })
  );

  assign N135 = icache_pkt_i[44:39] == paddr_tl[11:6];

  bsg_decode_00000008
  tag_mem_way_decode
  (
    .i(tag_mem_pkt_i[28:26]),
    .o(tag_mem_way_one_hot)
  );

  assign N145 = tag_mem_pkt_i[2] | tag_mem_pkt_i[1];
  assign N146 = N145 | N144;
  assign N149 = tag_mem_pkt_i[2] | N148;
  assign N150 = N149 | tag_mem_pkt_i[0];
  assign N152 = tag_mem_pkt_i[2] | N148;
  assign N153 = N152 | N144;
  assign N155 = N148 & N144;
  assign N157 = tag_mem_pkt_i[2] | tag_mem_pkt_i[1];
  assign N158 = N157 | N144;
  assign N160 = tag_mem_pkt_i[2] | N148;
  assign N161 = N160 | tag_mem_pkt_i[0];
  assign N163 = tag_mem_pkt_i[2] | N148;
  assign N164 = N163 | N144;
  assign N166 = N148 & N144;
  assign N168 = tag_mem_pkt_i[2] | tag_mem_pkt_i[1];
  assign N169 = N168 | N144;
  assign N171 = tag_mem_pkt_i[2] | N148;
  assign N172 = N171 | tag_mem_pkt_i[0];
  assign N174 = tag_mem_pkt_i[2] | N148;
  assign N175 = N174 | N144;
  assign N177 = N148 & N144;
  assign N179 = tag_mem_pkt_i[2] | tag_mem_pkt_i[1];
  assign N180 = N179 | N144;
  assign N182 = tag_mem_pkt_i[2] | N148;
  assign N183 = N182 | tag_mem_pkt_i[0];
  assign N185 = tag_mem_pkt_i[2] | N148;
  assign N186 = N185 | N144;
  assign N188 = N148 & N144;
  assign N190 = tag_mem_pkt_i[2] | tag_mem_pkt_i[1];
  assign N191 = N190 | N144;
  assign N193 = tag_mem_pkt_i[2] | N148;
  assign N194 = N193 | tag_mem_pkt_i[0];
  assign N196 = tag_mem_pkt_i[2] | N148;
  assign N197 = N196 | N144;
  assign N199 = N148 & N144;
  assign N201 = tag_mem_pkt_i[2] | tag_mem_pkt_i[1];
  assign N202 = N201 | N144;
  assign N204 = tag_mem_pkt_i[2] | N148;
  assign N205 = N204 | tag_mem_pkt_i[0];
  assign N207 = tag_mem_pkt_i[2] | N148;
  assign N208 = N207 | N144;
  assign N210 = N148 & N144;
  assign N212 = tag_mem_pkt_i[2] | tag_mem_pkt_i[1];
  assign N213 = N212 | N144;
  assign N215 = tag_mem_pkt_i[2] | N148;
  assign N216 = N215 | tag_mem_pkt_i[0];
  assign N218 = tag_mem_pkt_i[2] | N148;
  assign N219 = N218 | N144;
  assign N221 = N148 & N144;
  assign N223 = tag_mem_pkt_i[2] | tag_mem_pkt_i[1];
  assign N224 = N223 | N144;
  assign N226 = tag_mem_pkt_i[2] | N148;
  assign N227 = N226 | tag_mem_pkt_i[0];
  assign N229 = tag_mem_pkt_i[2] | N148;
  assign N230 = N229 | N144;
  assign N232 = N148 & N144;

  bsg_dff_00000003
  tag_mem_pkt_way_reg
  (
    .clk_i(clk_i),
    .data_i(tag_mem_pkt_i[28:26]),
    .data_o(tag_mem_pkt_way_r)
  );

  assign tag_mem_o[22] = (N241)? tag_mem_data_lo[22] : 
                         (N243)? tag_mem_data_lo[45] : 
                         (N245)? tag_mem_data_lo[68] : 
                         (N247)? tag_mem_data_lo[91] : 
                         (N242)? tag_mem_data_lo[114] : 
                         (N244)? tag_mem_data_lo[137] : 
                         (N246)? tag_mem_data_lo[160] : 
                         (N248)? tag_mem_data_lo[183] : 1'b0;
  assign tag_mem_o[21] = (N241)? tag_mem_data_lo[21] : 
                         (N243)? tag_mem_data_lo[44] : 
                         (N245)? tag_mem_data_lo[67] : 
                         (N247)? tag_mem_data_lo[90] : 
                         (N242)? tag_mem_data_lo[113] : 
                         (N244)? tag_mem_data_lo[136] : 
                         (N246)? tag_mem_data_lo[159] : 
                         (N248)? tag_mem_data_lo[182] : 1'b0;
  assign tag_mem_o[20] = (N241)? tag_mem_data_lo[20] : 
                         (N243)? tag_mem_data_lo[43] : 
                         (N245)? tag_mem_data_lo[66] : 
                         (N247)? tag_mem_data_lo[89] : 
                         (N242)? tag_mem_data_lo[112] : 
                         (N244)? tag_mem_data_lo[135] : 
                         (N246)? tag_mem_data_lo[158] : 
                         (N248)? tag_mem_data_lo[181] : 1'b0;
  assign tag_mem_o[19] = (N241)? tag_mem_data_lo[19] : 
                         (N243)? tag_mem_data_lo[42] : 
                         (N245)? tag_mem_data_lo[65] : 
                         (N247)? tag_mem_data_lo[88] : 
                         (N242)? tag_mem_data_lo[111] : 
                         (N244)? tag_mem_data_lo[134] : 
                         (N246)? tag_mem_data_lo[157] : 
                         (N248)? tag_mem_data_lo[180] : 1'b0;
  assign tag_mem_o[18] = (N241)? tag_mem_data_lo[18] : 
                         (N243)? tag_mem_data_lo[41] : 
                         (N245)? tag_mem_data_lo[64] : 
                         (N247)? tag_mem_data_lo[87] : 
                         (N242)? tag_mem_data_lo[110] : 
                         (N244)? tag_mem_data_lo[133] : 
                         (N246)? tag_mem_data_lo[156] : 
                         (N248)? tag_mem_data_lo[179] : 1'b0;
  assign tag_mem_o[17] = (N241)? tag_mem_data_lo[17] : 
                         (N243)? tag_mem_data_lo[40] : 
                         (N245)? tag_mem_data_lo[63] : 
                         (N247)? tag_mem_data_lo[86] : 
                         (N242)? tag_mem_data_lo[109] : 
                         (N244)? tag_mem_data_lo[132] : 
                         (N246)? tag_mem_data_lo[155] : 
                         (N248)? tag_mem_data_lo[178] : 1'b0;
  assign tag_mem_o[16] = (N241)? tag_mem_data_lo[16] : 
                         (N243)? tag_mem_data_lo[39] : 
                         (N245)? tag_mem_data_lo[62] : 
                         (N247)? tag_mem_data_lo[85] : 
                         (N242)? tag_mem_data_lo[108] : 
                         (N244)? tag_mem_data_lo[131] : 
                         (N246)? tag_mem_data_lo[154] : 
                         (N248)? tag_mem_data_lo[177] : 1'b0;
  assign tag_mem_o[15] = (N241)? tag_mem_data_lo[15] : 
                         (N243)? tag_mem_data_lo[38] : 
                         (N245)? tag_mem_data_lo[61] : 
                         (N247)? tag_mem_data_lo[84] : 
                         (N242)? tag_mem_data_lo[107] : 
                         (N244)? tag_mem_data_lo[130] : 
                         (N246)? tag_mem_data_lo[153] : 
                         (N248)? tag_mem_data_lo[176] : 1'b0;
  assign tag_mem_o[14] = (N241)? tag_mem_data_lo[14] : 
                         (N243)? tag_mem_data_lo[37] : 
                         (N245)? tag_mem_data_lo[60] : 
                         (N247)? tag_mem_data_lo[83] : 
                         (N242)? tag_mem_data_lo[106] : 
                         (N244)? tag_mem_data_lo[129] : 
                         (N246)? tag_mem_data_lo[152] : 
                         (N248)? tag_mem_data_lo[175] : 1'b0;
  assign tag_mem_o[13] = (N241)? tag_mem_data_lo[13] : 
                         (N243)? tag_mem_data_lo[36] : 
                         (N245)? tag_mem_data_lo[59] : 
                         (N247)? tag_mem_data_lo[82] : 
                         (N242)? tag_mem_data_lo[105] : 
                         (N244)? tag_mem_data_lo[128] : 
                         (N246)? tag_mem_data_lo[151] : 
                         (N248)? tag_mem_data_lo[174] : 1'b0;
  assign tag_mem_o[12] = (N241)? tag_mem_data_lo[12] : 
                         (N243)? tag_mem_data_lo[35] : 
                         (N245)? tag_mem_data_lo[58] : 
                         (N247)? tag_mem_data_lo[81] : 
                         (N242)? tag_mem_data_lo[104] : 
                         (N244)? tag_mem_data_lo[127] : 
                         (N246)? tag_mem_data_lo[150] : 
                         (N248)? tag_mem_data_lo[173] : 1'b0;
  assign tag_mem_o[11] = (N241)? tag_mem_data_lo[11] : 
                         (N243)? tag_mem_data_lo[34] : 
                         (N245)? tag_mem_data_lo[57] : 
                         (N247)? tag_mem_data_lo[80] : 
                         (N242)? tag_mem_data_lo[103] : 
                         (N244)? tag_mem_data_lo[126] : 
                         (N246)? tag_mem_data_lo[149] : 
                         (N248)? tag_mem_data_lo[172] : 1'b0;
  assign tag_mem_o[10] = (N241)? tag_mem_data_lo[10] : 
                         (N243)? tag_mem_data_lo[33] : 
                         (N245)? tag_mem_data_lo[56] : 
                         (N247)? tag_mem_data_lo[79] : 
                         (N242)? tag_mem_data_lo[102] : 
                         (N244)? tag_mem_data_lo[125] : 
                         (N246)? tag_mem_data_lo[148] : 
                         (N248)? tag_mem_data_lo[171] : 1'b0;
  assign tag_mem_o[9] = (N241)? tag_mem_data_lo[9] : 
                        (N243)? tag_mem_data_lo[32] : 
                        (N245)? tag_mem_data_lo[55] : 
                        (N247)? tag_mem_data_lo[78] : 
                        (N242)? tag_mem_data_lo[101] : 
                        (N244)? tag_mem_data_lo[124] : 
                        (N246)? tag_mem_data_lo[147] : 
                        (N248)? tag_mem_data_lo[170] : 1'b0;
  assign tag_mem_o[8] = (N241)? tag_mem_data_lo[8] : 
                        (N243)? tag_mem_data_lo[31] : 
                        (N245)? tag_mem_data_lo[54] : 
                        (N247)? tag_mem_data_lo[77] : 
                        (N242)? tag_mem_data_lo[100] : 
                        (N244)? tag_mem_data_lo[123] : 
                        (N246)? tag_mem_data_lo[146] : 
                        (N248)? tag_mem_data_lo[169] : 1'b0;
  assign tag_mem_o[7] = (N241)? tag_mem_data_lo[7] : 
                        (N243)? tag_mem_data_lo[30] : 
                        (N245)? tag_mem_data_lo[53] : 
                        (N247)? tag_mem_data_lo[76] : 
                        (N242)? tag_mem_data_lo[99] : 
                        (N244)? tag_mem_data_lo[122] : 
                        (N246)? tag_mem_data_lo[145] : 
                        (N248)? tag_mem_data_lo[168] : 1'b0;
  assign tag_mem_o[6] = (N241)? tag_mem_data_lo[6] : 
                        (N243)? tag_mem_data_lo[29] : 
                        (N245)? tag_mem_data_lo[52] : 
                        (N247)? tag_mem_data_lo[75] : 
                        (N242)? tag_mem_data_lo[98] : 
                        (N244)? tag_mem_data_lo[121] : 
                        (N246)? tag_mem_data_lo[144] : 
                        (N248)? tag_mem_data_lo[167] : 1'b0;
  assign tag_mem_o[5] = (N241)? tag_mem_data_lo[5] : 
                        (N243)? tag_mem_data_lo[28] : 
                        (N245)? tag_mem_data_lo[51] : 
                        (N247)? tag_mem_data_lo[74] : 
                        (N242)? tag_mem_data_lo[97] : 
                        (N244)? tag_mem_data_lo[120] : 
                        (N246)? tag_mem_data_lo[143] : 
                        (N248)? tag_mem_data_lo[166] : 1'b0;
  assign tag_mem_o[4] = (N241)? tag_mem_data_lo[4] : 
                        (N243)? tag_mem_data_lo[27] : 
                        (N245)? tag_mem_data_lo[50] : 
                        (N247)? tag_mem_data_lo[73] : 
                        (N242)? tag_mem_data_lo[96] : 
                        (N244)? tag_mem_data_lo[119] : 
                        (N246)? tag_mem_data_lo[142] : 
                        (N248)? tag_mem_data_lo[165] : 1'b0;
  assign tag_mem_o[3] = (N241)? tag_mem_data_lo[3] : 
                        (N243)? tag_mem_data_lo[26] : 
                        (N245)? tag_mem_data_lo[49] : 
                        (N247)? tag_mem_data_lo[72] : 
                        (N242)? tag_mem_data_lo[95] : 
                        (N244)? tag_mem_data_lo[118] : 
                        (N246)? tag_mem_data_lo[141] : 
                        (N248)? tag_mem_data_lo[164] : 1'b0;
  assign tag_mem_o[2] = (N241)? tag_mem_data_lo[2] : 
                        (N243)? tag_mem_data_lo[25] : 
                        (N245)? tag_mem_data_lo[48] : 
                        (N247)? tag_mem_data_lo[71] : 
                        (N242)? tag_mem_data_lo[94] : 
                        (N244)? tag_mem_data_lo[117] : 
                        (N246)? tag_mem_data_lo[140] : 
                        (N248)? tag_mem_data_lo[163] : 1'b0;
  assign tag_mem_o[1] = (N241)? tag_mem_data_lo[1] : 
                        (N243)? tag_mem_data_lo[24] : 
                        (N245)? tag_mem_data_lo[47] : 
                        (N247)? tag_mem_data_lo[70] : 
                        (N242)? tag_mem_data_lo[93] : 
                        (N244)? tag_mem_data_lo[116] : 
                        (N246)? tag_mem_data_lo[139] : 
                        (N248)? tag_mem_data_lo[162] : 1'b0;
  assign tag_mem_o[0] = (N241)? tag_mem_data_lo[0] : 
                        (N243)? tag_mem_data_lo[23] : 
                        (N245)? tag_mem_data_lo[46] : 
                        (N247)? tag_mem_data_lo[69] : 
                        (N242)? tag_mem_data_lo[92] : 
                        (N244)? tag_mem_data_lo[115] : 
                        (N246)? tag_mem_data_lo[138] : 
                        (N248)? tag_mem_data_lo[161] : 1'b0;

  bsg_decode_00000008
  bypass_bank_decode
  (
    .i(icache_pkt_i[38:36]),
    .o(vaddr_bank_dec)
  );


  bsg_adder_one_hot_00000008
  data_mem_bank_select_adder
  (
    .a_i(hit_v_tl),
    .b_i(vaddr_bank_dec),
    .o(data_mem_bypass_select)
  );


  bsg_rotate_left_00000080
  write_data_rotate
  (
    .data_i(data_mem_pkt_i[133:6]),
    .rot_i({ data_mem_pkt_i[134:134], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .o(data_mem_pkt_fill_data_li)
  );


  bsg_expand_bitmask_00000004_00000002
  fill_mask_expand
  (
    .i(data_mem_pkt_i[5:2]),
    .o(data_mem_pkt_fill_mask_expanded)
  );


  bsg_rotate_left_00000008
  write_mask_rotate
  (
    .data_i(data_mem_pkt_fill_mask_expanded),
    .rot_i(data_mem_pkt_i[136:134]),
    .o(data_mem_write_bank_mask)
  );

  assign N249 = icache_pkt_i[44:39] == paddr_tl[11:6];
  assign N250 = icache_pkt_i[71:45] == vaddr_vtag_tl;

  bsg_dff_00000003
  data_mem_pkt_way_reg
  (
    .clk_i(clk_i),
    .data_i(data_mem_pkt_i[136:134]),
    .data_o(data_mem_pkt_way_r)
  );


  bsg_rotate_right_00000200
  read_data_rotate
  (
    .data_i(data_mem_data_lo),
    .rot_i({ data_mem_pkt_way_r, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .o(data_mem_o)
  );


  bsg_lru_pseudo_tree_decode_00000008
  lru_decode
  (
    .way_id_i(hit_index_tv),
    .data_o(lru_decode_data_lo),
    .mask_o(lru_decode_mask_lo)
  );

  assign { N341, N340, N339, N338, N337, N336, N335, N334 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, data_mem_pkt_v_i } << data_mem_pkt_i[136:134];
  assign { N349, N348, N347, N346, N345, N344, N343, N342 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tag_mem_pkt_v_i } << tag_mem_pkt_i[28:26];
  assign N353 = tag_mem_data_lo[182] | tag_mem_data_lo[183];
  assign N354 = tag_mem_data_lo[181] | N353;
  assign N355 = tag_mem_data_lo[159] | tag_mem_data_lo[160];
  assign N356 = tag_mem_data_lo[158] | N355;
  assign N357 = tag_mem_data_lo[136] | tag_mem_data_lo[137];
  assign N358 = tag_mem_data_lo[135] | N357;
  assign N359 = tag_mem_data_lo[113] | tag_mem_data_lo[114];
  assign N360 = tag_mem_data_lo[112] | N359;
  assign N361 = tag_mem_data_lo[90] | tag_mem_data_lo[91];
  assign N362 = tag_mem_data_lo[89] | N361;
  assign N363 = tag_mem_data_lo[67] | tag_mem_data_lo[68];
  assign N364 = tag_mem_data_lo[66] | N363;
  assign N365 = tag_mem_data_lo[44] | tag_mem_data_lo[45];
  assign N366 = tag_mem_data_lo[43] | N365;
  assign N367 = tag_mem_data_lo[21] | tag_mem_data_lo[22];
  assign N368 = tag_mem_data_lo[20] | N367;
  assign N369 = ~tag_mem_pkt_i[2];
  assign N370 = tag_mem_pkt_i[1] | N369;
  assign N371 = tag_mem_pkt_i[0] | N370;
  assign N372 = ~N371;
  assign N373 = tag_mem_pkt_i[1] | N369;
  assign N374 = tag_mem_pkt_i[0] | N373;
  assign N375 = ~data_mem_pkt_i[0];
  assign N376 = N375 | data_mem_pkt_i[1];
  assign N377 = ~N376;
  assign N378 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N379 = ~N378;
  assign N380 = N375 | data_mem_pkt_i[1];
  assign N381 = ~N380;
  assign N382 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N383 = ~N382;
  assign N384 = N375 | data_mem_pkt_i[1];
  assign N385 = ~N384;
  assign N386 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N387 = ~N386;
  assign N388 = N375 | data_mem_pkt_i[1];
  assign N389 = ~N388;
  assign N390 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N391 = ~N390;
  assign N392 = N375 | data_mem_pkt_i[1];
  assign N393 = ~N392;
  assign N394 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N395 = ~N394;
  assign N396 = N375 | data_mem_pkt_i[1];
  assign N397 = ~N396;
  assign N398 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N399 = ~N398;
  assign N400 = N375 | data_mem_pkt_i[1];
  assign N401 = ~N400;
  assign N402 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N403 = ~N402;
  assign N404 = N375 | data_mem_pkt_i[1];
  assign N405 = ~N404;
  assign N406 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N407 = ~N406;
  assign N408 = ~stat_mem_pkt_i[0];
  assign N409 = N408 | stat_mem_pkt_i[1];
  assign N410 = ~state_r[0];
  assign N411 = N410 | state_r[1];
  assign N412 = ~N411;
  assign N413 = ~data_mem_pkt_i[1];
  assign N414 = data_mem_pkt_i[0] | N413;
  assign N415 = ~N414;
  assign N416 = ~state_r[1];
  assign N417 = state_r[0] | N416;
  assign N418 = ~N417;
  assign N419 = state_r[0] | state_r[1];
  assign N420 = ~N419;
  assign \data_mem_lines_1_.data_mem_pkt_offset  = 1'b1 - data_mem_pkt_i[136:134];
  assign \data_mem_lines_3_.data_mem_pkt_offset  = { 1'b1, 1'b1 } - data_mem_pkt_i[136:134];
  assign \data_mem_lines_7_.data_mem_pkt_offset  = { 1'b1, 1'b1, 1'b1 } - data_mem_pkt_i[136:134];
  assign \data_mem_lines_0_.data_mem_pkt_offset  = 1'b0 - data_mem_pkt_i[136:134];
  assign \data_mem_lines_2_.data_mem_pkt_offset  = { 1'b1, 1'b0 } - data_mem_pkt_i[136:134];
  assign \data_mem_lines_4_.data_mem_pkt_offset  = { 1'b1, 1'b0, 1'b0 } - data_mem_pkt_i[136:134];
  assign \data_mem_lines_5_.data_mem_pkt_offset  = { 1'b1, 1'b0, 1'b1 } - data_mem_pkt_i[136:134];
  assign \data_mem_lines_6_.data_mem_pkt_offset  = { 1'b1, 1'b1, 1'b0 } - data_mem_pkt_i[136:134];
  assign tl_we = (N0)? N101 : 
                 (N1)? N102 : 1'b0;
  assign N0 = N100;
  assign N1 = N99;
  assign tv_we_o = (N2)? yumi_i : 
                   (N3)? N420 : 1'b0;
  assign N2 = v_tv_r;
  assign N3 = N119;
  assign paddr_tv_n = (N4)? cache_req_o[47:8] : 
                      (N5)? { ptag_i, paddr_tl } : 1'b0;
  assign N4 = N121;
  assign N5 = N120;
  assign lru_way_li = (N6)? invalid_way_tv : 
                      (N7)? lru_encode : 1'b0;
  assign N6 = invalid_exist_tv;
  assign N7 = N122;
  assign cache_req_o[6:4] = (N8)? { 1'b0, 1'b0, 1'b0 } : 
                            (N127)? { 1'b0, 1'b1, 1'b1 } : 
                            (N125)? { 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N8 = cached_req;
  assign cache_req_metadata_o[3:1] = (N9)? metadata_hit_index_r : 
                                     (N10)? lru_way_li : 1'b0;
  assign N9 = metadata_hit_r;
  assign N10 = N128;
  assign { N132, N131 } = (N11)? { 1'b1, 1'b0 } : 
                          (N12)? state_r : 1'b0;
  assign N11 = complete_recv;
  assign N12 = N130;
  assign { N134, N133 } = (N13)? { 1'b0, 1'b1 } : 
                          (N14)? { N132, N131 } : 1'b0;
  assign N13 = N410;
  assign N14 = state_r[0];
  assign state_n = (N15)? { N134, N133 } : 
                   (N16)? { 1'b0, 1'b0 } : 1'b0;
  assign N15 = N416;
  assign N16 = state_r[1];
  assign { N143, N142, N141, N140, N139, N138 } = (N17)? paddr_tl[11:6] : 
                                                  (N18)? icache_pkt_i[44:39] : 1'b0;
  assign N17 = do_recover;
  assign N18 = N137;
  assign tag_mem_addr_li = (N19)? { N143, N142, N141, N140, N139, N138 } : 
                           (N20)? tag_mem_pkt_i[34:29] : 1'b0;
  assign N19 = tag_mem_fast_read;
  assign N20 = N136;
  assign tag_mem_data_li[22:0] = (N21)? tag_mem_pkt_i[25:3] : 
                                 (N22)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N23)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N21 = N147;
  assign N22 = N151;
  assign N23 = N154;
  assign N24 = N156;
  assign tag_mem_w_mask_li[22:0] = (N21)? { tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0] } : 
                                   (N22)? { tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N23)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N24)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[45:23] = (N25)? tag_mem_pkt_i[25:3] : 
                                  (N26)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N27)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N28)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N25 = N159;
  assign N26 = N162;
  assign N27 = N165;
  assign N28 = N167;
  assign tag_mem_w_mask_li[45:23] = (N25)? { tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1] } : 
                                    (N26)? { tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N27)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N28)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[68:46] = (N29)? tag_mem_pkt_i[25:3] : 
                                  (N30)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N31)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N32)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N29 = N170;
  assign N30 = N173;
  assign N31 = N176;
  assign N32 = N178;
  assign tag_mem_w_mask_li[68:46] = (N29)? { tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2] } : 
                                    (N30)? { tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N31)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N32)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[91:69] = (N33)? tag_mem_pkt_i[25:3] : 
                                  (N34)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N36)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N33 = N181;
  assign N34 = N184;
  assign N35 = N187;
  assign N36 = N189;
  assign tag_mem_w_mask_li[91:69] = (N33)? { tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3] } : 
                                    (N34)? { tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N35)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N36)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[114:92] = (N37)? tag_mem_pkt_i[25:3] : 
                                   (N38)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N39)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N40)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N37 = N192;
  assign N38 = N195;
  assign N39 = N198;
  assign N40 = N200;
  assign tag_mem_w_mask_li[114:92] = (N37)? { tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4] } : 
                                     (N38)? { tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                     (N39)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                     (N40)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[137:115] = (N41)? tag_mem_pkt_i[25:3] : 
                                    (N42)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N43)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N44)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N41 = N203;
  assign N42 = N206;
  assign N43 = N209;
  assign N44 = N211;
  assign tag_mem_w_mask_li[137:115] = (N41)? { tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5] } : 
                                      (N42)? { tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N43)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N44)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[160:138] = (N45)? tag_mem_pkt_i[25:3] : 
                                    (N46)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N47)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N48)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N45 = N214;
  assign N46 = N217;
  assign N47 = N220;
  assign N48 = N222;
  assign tag_mem_w_mask_li[160:138] = (N45)? { tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6] } : 
                                      (N46)? { tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N47)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N48)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[183:161] = (N49)? tag_mem_pkt_i[25:3] : 
                                    (N50)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N51)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N52)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N49 = N225;
  assign N50 = N228;
  assign N51 = N231;
  assign N52 = N233;
  assign tag_mem_w_mask_li[183:161] = (N49)? { tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7] } : 
                                      (N50)? { tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N51)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N52)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign { N260, N259, N258, N257, N256, N255, N254, N253, N252 } = (N17)? paddr_tl[11:3] : 
                                                                    (N18)? icache_pkt_i[44:36] : 1'b0;
  assign data_mem_addr_li[8:0] = (N53)? { N260, N259, N258, N257, N256, N255, N254, N253, N252 } : 
                                 (N251)? { data_mem_pkt_i[142:137], \data_mem_lines_0_.data_mem_pkt_offset  } : 1'b0;
  assign N53 = data_mem_fast_read[0];
  assign { N270, N269, N268, N267, N266, N265, N264, N263, N262 } = (N17)? paddr_tl[11:3] : 
                                                                    (N18)? icache_pkt_i[44:36] : 1'b0;
  assign data_mem_addr_li[17:9] = (N54)? { N270, N269, N268, N267, N266, N265, N264, N263, N262 } : 
                                  (N261)? { data_mem_pkt_i[142:137], \data_mem_lines_1_.data_mem_pkt_offset  } : 1'b0;
  assign N54 = data_mem_fast_read[1];
  assign { N280, N279, N278, N277, N276, N275, N274, N273, N272 } = (N17)? paddr_tl[11:3] : 
                                                                    (N18)? icache_pkt_i[44:36] : 1'b0;
  assign data_mem_addr_li[26:18] = (N55)? { N280, N279, N278, N277, N276, N275, N274, N273, N272 } : 
                                   (N271)? { data_mem_pkt_i[142:137], \data_mem_lines_2_.data_mem_pkt_offset  } : 1'b0;
  assign N55 = data_mem_fast_read[2];
  assign { N290, N289, N288, N287, N286, N285, N284, N283, N282 } = (N17)? paddr_tl[11:3] : 
                                                                    (N18)? icache_pkt_i[44:36] : 1'b0;
  assign data_mem_addr_li[35:27] = (N56)? { N290, N289, N288, N287, N286, N285, N284, N283, N282 } : 
                                   (N281)? { data_mem_pkt_i[142:137], \data_mem_lines_3_.data_mem_pkt_offset  } : 1'b0;
  assign N56 = data_mem_fast_read[3];
  assign { N300, N299, N298, N297, N296, N295, N294, N293, N292 } = (N17)? paddr_tl[11:3] : 
                                                                    (N18)? icache_pkt_i[44:36] : 1'b0;
  assign data_mem_addr_li[44:36] = (N57)? { N300, N299, N298, N297, N296, N295, N294, N293, N292 } : 
                                   (N291)? { data_mem_pkt_i[142:137], \data_mem_lines_4_.data_mem_pkt_offset  } : 1'b0;
  assign N57 = data_mem_fast_read[4];
  assign { N310, N309, N308, N307, N306, N305, N304, N303, N302 } = (N17)? paddr_tl[11:3] : 
                                                                    (N18)? icache_pkt_i[44:36] : 1'b0;
  assign data_mem_addr_li[53:45] = (N58)? { N310, N309, N308, N307, N306, N305, N304, N303, N302 } : 
                                   (N301)? { data_mem_pkt_i[142:137], \data_mem_lines_5_.data_mem_pkt_offset  } : 1'b0;
  assign N58 = data_mem_fast_read[5];
  assign { N320, N319, N318, N317, N316, N315, N314, N313, N312 } = (N17)? paddr_tl[11:3] : 
                                                                    (N18)? icache_pkt_i[44:36] : 1'b0;
  assign data_mem_addr_li[62:54] = (N59)? { N320, N319, N318, N317, N316, N315, N314, N313, N312 } : 
                                   (N311)? { data_mem_pkt_i[142:137], \data_mem_lines_6_.data_mem_pkt_offset  } : 1'b0;
  assign N59 = data_mem_fast_read[6];
  assign { N330, N329, N328, N327, N326, N325, N324, N323, N322 } = (N17)? paddr_tl[11:3] : 
                                                                    (N18)? icache_pkt_i[44:36] : 1'b0;
  assign data_mem_addr_li[71:63] = (N60)? { N330, N329, N328, N327, N326, N325, N324, N323, N322 } : 
                                   (N321)? { data_mem_pkt_i[142:137], \data_mem_lines_7_.data_mem_pkt_offset  } : 1'b0;
  assign N60 = data_mem_fast_read[7];
  assign data_mem_pkt_yumi_o = (N61)? data_mem_pkt_v_i : 
                               (N62)? N331 : 1'b0;
  assign N61 = N415;
  assign N62 = N414;
  assign stat_mem_addr_li = (N63)? cache_req_o[19:14] : 
                            (N333)? stat_mem_pkt_i[10:5] : 1'b0;
  assign N63 = N332;
  assign { stat_mem_data_li_lru__6_, stat_mem_data_li_lru__5_, stat_mem_data_li_lru__4_, stat_mem_data_li_lru__3_, stat_mem_data_li_lru__2_, stat_mem_data_li_lru__1_, stat_mem_data_li_lru__0_ } = (N64)? lru_decode_data_lo : 
                                                                                                                                                                                                    (N65)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N64 = stat_mem_fast_write;
  assign N65 = N607;
  assign { stat_mem_mask_li_lru__6_, stat_mem_mask_li_lru__5_, stat_mem_mask_li_lru__4_, stat_mem_mask_li_lru__3_, stat_mem_mask_li_lru__2_, stat_mem_mask_li_lru__1_, stat_mem_mask_li_lru__0_ } = (N64)? lru_decode_mask_lo : 
                                                                                                                                                                                                    (N65)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign critical_recv = N427 & N429;
  assign N427 = N424 & N426;
  assign N424 = N421 & N423;
  assign N421 = N412 & cache_req_critical_i;
  assign N423 = N422 | stat_mem_pkt_yumi_o;
  assign N422 = ~stat_mem_pkt_v_i;
  assign N426 = N425 | tag_mem_pkt_yumi_o;
  assign N425 = ~tag_mem_pkt_v_i;
  assign N429 = N428 | data_mem_pkt_yumi_o;
  assign N428 = ~data_mem_pkt_v_i;
  assign complete_recv = N434 & N435;
  assign N434 = N432 & N433;
  assign N432 = N430 & N431;
  assign N430 = N412 & cache_req_last_i;
  assign N431 = N422 | stat_mem_pkt_yumi_o;
  assign N433 = N425 | tag_mem_pkt_yumi_o;
  assign N435 = N428 | data_mem_pkt_yumi_o;
  assign yumi_o = v_i & tl_we;
  assign N99 = ~v_tl_r;
  assign N100 = v_tl_r;
  assign N101 = tv_we_o | force_i;
  assign N102 = ~cache_req_lock_i;
  assign _0_net_ = reset_i | tl_flush_i;
  assign \tag_comp_tl_0_.tag_match_tl  = N444 & N103;
  assign N444 = ptag_v_i & N443;
  assign N443 = ~N442;
  assign N442 = N441 | ptag_i[20];
  assign N441 = N440 | ptag_i[21];
  assign N440 = N439 | ptag_i[22];
  assign N439 = N438 | ptag_i[23];
  assign N438 = N437 | ptag_i[24];
  assign N437 = N436 | ptag_i[25];
  assign N436 = ptag_i[27] | ptag_i[26];
  assign hit_v_tl[0] = \tag_comp_tl_0_.tag_match_tl  & N445;
  assign N445 = N104 & N368;
  assign \tag_comp_tl_1_.tag_match_tl  = N454 & N105;
  assign N454 = ptag_v_i & N453;
  assign N453 = ~N452;
  assign N452 = N451 | ptag_i[20];
  assign N451 = N450 | ptag_i[21];
  assign N450 = N449 | ptag_i[22];
  assign N449 = N448 | ptag_i[23];
  assign N448 = N447 | ptag_i[24];
  assign N447 = N446 | ptag_i[25];
  assign N446 = ptag_i[27] | ptag_i[26];
  assign hit_v_tl[1] = \tag_comp_tl_1_.tag_match_tl  & N455;
  assign N455 = N106 & N366;
  assign \tag_comp_tl_2_.tag_match_tl  = N464 & N107;
  assign N464 = ptag_v_i & N463;
  assign N463 = ~N462;
  assign N462 = N461 | ptag_i[20];
  assign N461 = N460 | ptag_i[21];
  assign N460 = N459 | ptag_i[22];
  assign N459 = N458 | ptag_i[23];
  assign N458 = N457 | ptag_i[24];
  assign N457 = N456 | ptag_i[25];
  assign N456 = ptag_i[27] | ptag_i[26];
  assign hit_v_tl[2] = \tag_comp_tl_2_.tag_match_tl  & N465;
  assign N465 = N108 & N364;
  assign \tag_comp_tl_3_.tag_match_tl  = N474 & N109;
  assign N474 = ptag_v_i & N473;
  assign N473 = ~N472;
  assign N472 = N471 | ptag_i[20];
  assign N471 = N470 | ptag_i[21];
  assign N470 = N469 | ptag_i[22];
  assign N469 = N468 | ptag_i[23];
  assign N468 = N467 | ptag_i[24];
  assign N467 = N466 | ptag_i[25];
  assign N466 = ptag_i[27] | ptag_i[26];
  assign hit_v_tl[3] = \tag_comp_tl_3_.tag_match_tl  & N475;
  assign N475 = N110 & N362;
  assign \tag_comp_tl_4_.tag_match_tl  = N484 & N111;
  assign N484 = ptag_v_i & N483;
  assign N483 = ~N482;
  assign N482 = N481 | ptag_i[20];
  assign N481 = N480 | ptag_i[21];
  assign N480 = N479 | ptag_i[22];
  assign N479 = N478 | ptag_i[23];
  assign N478 = N477 | ptag_i[24];
  assign N477 = N476 | ptag_i[25];
  assign N476 = ptag_i[27] | ptag_i[26];
  assign hit_v_tl[4] = \tag_comp_tl_4_.tag_match_tl  & N485;
  assign N485 = N112 & N360;
  assign \tag_comp_tl_5_.tag_match_tl  = N494 & N113;
  assign N494 = ptag_v_i & N493;
  assign N493 = ~N492;
  assign N492 = N491 | ptag_i[20];
  assign N491 = N490 | ptag_i[21];
  assign N490 = N489 | ptag_i[22];
  assign N489 = N488 | ptag_i[23];
  assign N488 = N487 | ptag_i[24];
  assign N487 = N486 | ptag_i[25];
  assign N486 = ptag_i[27] | ptag_i[26];
  assign hit_v_tl[5] = \tag_comp_tl_5_.tag_match_tl  & N495;
  assign N495 = N114 & N358;
  assign \tag_comp_tl_6_.tag_match_tl  = N504 & N115;
  assign N504 = ptag_v_i & N503;
  assign N503 = ~N502;
  assign N502 = N501 | ptag_i[20];
  assign N501 = N500 | ptag_i[21];
  assign N500 = N499 | ptag_i[22];
  assign N499 = N498 | ptag_i[23];
  assign N498 = N497 | ptag_i[24];
  assign N497 = N496 | ptag_i[25];
  assign N496 = ptag_i[27] | ptag_i[26];
  assign hit_v_tl[6] = \tag_comp_tl_6_.tag_match_tl  & N505;
  assign N505 = N116 & N356;
  assign \tag_comp_tl_7_.tag_match_tl  = N514 & N117;
  assign N514 = ptag_v_i & N513;
  assign N513 = ~N512;
  assign N512 = N511 | ptag_i[20];
  assign N511 = N510 | ptag_i[21];
  assign N510 = N509 | ptag_i[22];
  assign N509 = N508 | ptag_i[23];
  assign N508 = N507 | ptag_i[24];
  assign N507 = N506 | ptag_i[25];
  assign N506 = ptag_i[27] | ptag_i[26];
  assign hit_v_tl[7] = \tag_comp_tl_7_.tag_match_tl  & N515;
  assign N515 = N118 & N354;
  assign fetch_uncached_tl = decode_tl_r_fetch_op_ & ptag_uncached_i;
  assign spec_tl = N517 | N519;
  assign N517 = decode_tl_r_fetch_op_ & N516;
  assign N516 = ~ptag_v_i;
  assign N519 = N518 & ptag_nonidem_i;
  assign N518 = decode_tl_r_fetch_op_ & spec_tl_r;
  assign N119 = ~v_tv_r;
  assign _3_net_ = reset_i | tv_flush_i;
  assign _6_net_ = tv_we_o | critical_recv;
  assign N120 = ~critical_recv;
  assign N121 = critical_recv;
  assign _9_net_ = tv_we_o | critical_recv;
  assign _10_net__7_ = ~way_v_tv_r[7];
  assign _10_net__6_ = ~way_v_tv_r[6];
  assign _10_net__5_ = ~way_v_tv_r[5];
  assign _10_net__4_ = ~way_v_tv_r[4];
  assign _10_net__3_ = ~way_v_tv_r[3];
  assign _10_net__2_ = ~way_v_tv_r[2];
  assign _10_net__1_ = ~way_v_tv_r[1];
  assign _10_net__0_ = ~way_v_tv_r[0];
  assign N122 = ~invalid_exist_tv;
  assign hit_v_o = N523 & cache_req_o[115];
  assign N523 = N521 & N522;
  assign N521 = N520 & snoop_decode_fetch_op_;
  assign N520 = N420 & v_tv_r;
  assign N522 = ~snoop_spec;
  assign miss_v_o = N526 & N527;
  assign N526 = N525 & snoop_spec;
  assign N525 = N524 & snoop_decode_fetch_op_;
  assign N524 = N420 & v_tv_r;
  assign N527 = ~cache_req_o[115];
  assign fence_v_o = N529 & snoop_tv_r;
  assign N529 = N528 & snoop_decode_inval_op_;
  assign N528 = N420 & v_tv_r;
  assign cached_req = N535 & N536;
  assign N535 = N533 & N534;
  assign N533 = N531 & N532;
  assign N531 = snoop_decode_fetch_op_ & N530;
  assign N530 = ~snoop_tv_r;
  assign N532 = ~cache_req_o[115];
  assign N534 = ~snoop_uncached;
  assign N536 = ~snoop_spec;
  assign uncached_req = N540 & N541;
  assign N540 = N539 & snoop_uncached;
  assign N539 = N537 & N538;
  assign N537 = snoop_decode_fetch_op_ & N530;
  assign N538 = ~cache_req_o[115];
  assign N541 = ~snoop_spec;
  assign inval_req = snoop_decode_inval_op_ & N530;
  assign cache_req_v_o = N545 & N546;
  assign N545 = N542 & N544;
  assign N542 = N420 & v_tv_r;
  assign N544 = N543 | inval_req;
  assign N543 = uncached_req | cached_req;
  assign N546 = ~tv_flush_i;
  assign N123 = ~cached_req;
  assign cache_req_o[50] = cached_req;
  assign cache_req_o[48] = N123;
  assign N124 = uncached_req | cached_req;
  assign N125 = ~N124;
  assign N126 = ~cached_req;
  assign N127 = uncached_req & N126;
  assign N128 = ~metadata_hit_r;
  assign N129 = ~cache_req_yumi_i;
  assign N130 = ~complete_recv;
  assign do_recover = N418 & N547;
  assign N547 = ~yumi_o;
  assign tag_mem_bypass = N548 & N135;
  assign N548 = v_tl_r & decode_tl_r_fetch_op_;
  assign tag_mem_fast_read = do_recover | N551;
  assign N551 = N549 & N550;
  assign N549 = yumi_o & decode_lo_fetch_op_;
  assign N550 = ~tag_mem_bypass;
  assign tag_mem_slow_read = tag_mem_pkt_yumi_o & N372;
  assign tag_mem_slow_write = tag_mem_pkt_yumi_o & N374;
  assign tag_mem_v_li = N553 | tag_mem_slow_write;
  assign N553 = N552 | tag_mem_slow_read;
  assign N552 = tag_mem_fast_read | 1'b0;
  assign tag_mem_w_li = 1'b0 | tag_mem_slow_write;
  assign N136 = ~tag_mem_fast_read;
  assign N137 = ~do_recover;
  assign tag_mem_pkt_yumi_o = tag_mem_pkt_v_i & N136;
  assign N144 = ~tag_mem_pkt_i[0];
  assign N147 = ~N146;
  assign N148 = ~tag_mem_pkt_i[1];
  assign N151 = ~N150;
  assign N154 = ~N153;
  assign N156 = tag_mem_pkt_i[2] | N155;
  assign N159 = ~N158;
  assign N162 = ~N161;
  assign N165 = ~N164;
  assign N167 = tag_mem_pkt_i[2] | N166;
  assign N170 = ~N169;
  assign N173 = ~N172;
  assign N176 = ~N175;
  assign N178 = tag_mem_pkt_i[2] | N177;
  assign N181 = ~N180;
  assign N184 = ~N183;
  assign N187 = ~N186;
  assign N189 = tag_mem_pkt_i[2] | N188;
  assign N192 = ~N191;
  assign N195 = ~N194;
  assign N198 = ~N197;
  assign N200 = tag_mem_pkt_i[2] | N199;
  assign N203 = ~N202;
  assign N206 = ~N205;
  assign N209 = ~N208;
  assign N211 = tag_mem_pkt_i[2] | N210;
  assign N214 = ~N213;
  assign N217 = ~N216;
  assign N220 = ~N219;
  assign N222 = tag_mem_pkt_i[2] | N221;
  assign N225 = ~N224;
  assign N228 = ~N227;
  assign N231 = ~N230;
  assign N233 = tag_mem_pkt_i[2] | N232;
  assign N234 = ~tag_mem_pkt_way_r[0];
  assign N235 = ~tag_mem_pkt_way_r[1];
  assign N236 = N234 & N235;
  assign N237 = N234 & tag_mem_pkt_way_r[1];
  assign N238 = tag_mem_pkt_way_r[0] & N235;
  assign N239 = tag_mem_pkt_way_r[0] & tag_mem_pkt_way_r[1];
  assign N240 = ~tag_mem_pkt_way_r[2];
  assign N241 = N236 & N240;
  assign N242 = N236 & tag_mem_pkt_way_r[2];
  assign N243 = N238 & N240;
  assign N244 = N238 & tag_mem_pkt_way_r[2];
  assign N245 = N237 & N240;
  assign N246 = N237 & tag_mem_pkt_way_r[2];
  assign N247 = N239 & N240;
  assign N248 = N239 & tag_mem_pkt_way_r[2];
  assign data_mem_bypass = N555 & N250;
  assign N555 = N554 & N249;
  assign N554 = v_tl_r & decode_tl_r_fetch_op_;
  assign data_mem_slow_read[0] = data_mem_pkt_yumi_o & N377;
  assign data_mem_slow_write[0] = N556 & data_mem_write_bank_mask[0];
  assign N556 = data_mem_pkt_yumi_o & N379;
  assign data_mem_fast_read[0] = do_recover | N560;
  assign N560 = N557 & N559;
  assign N557 = yumi_o & decode_lo_fetch_op_;
  assign N559 = N558 | data_mem_bypass_select[0];
  assign N558 = ~data_mem_bypass;
  assign data_mem_v_li[0] = N561 | data_mem_slow_write[0];
  assign N561 = data_mem_fast_read[0] | data_mem_slow_read[0];
  assign N251 = ~data_mem_fast_read[0];
  assign data_mem_slow_read[1] = data_mem_pkt_yumi_o & N381;
  assign data_mem_slow_write[1] = N562 & data_mem_write_bank_mask[1];
  assign N562 = data_mem_pkt_yumi_o & N383;
  assign data_mem_fast_read[1] = do_recover | N565;
  assign N565 = N563 & N564;
  assign N563 = yumi_o & decode_lo_fetch_op_;
  assign N564 = N558 | data_mem_bypass_select[1];
  assign data_mem_v_li[1] = N566 | data_mem_slow_write[1];
  assign N566 = data_mem_fast_read[1] | data_mem_slow_read[1];
  assign N261 = ~data_mem_fast_read[1];
  assign data_mem_slow_read[2] = data_mem_pkt_yumi_o & N385;
  assign data_mem_slow_write[2] = N567 & data_mem_write_bank_mask[2];
  assign N567 = data_mem_pkt_yumi_o & N387;
  assign data_mem_fast_read[2] = do_recover | N570;
  assign N570 = N568 & N569;
  assign N568 = yumi_o & decode_lo_fetch_op_;
  assign N569 = N558 | data_mem_bypass_select[2];
  assign data_mem_v_li[2] = N571 | data_mem_slow_write[2];
  assign N571 = data_mem_fast_read[2] | data_mem_slow_read[2];
  assign N271 = ~data_mem_fast_read[2];
  assign data_mem_slow_read[3] = data_mem_pkt_yumi_o & N389;
  assign data_mem_slow_write[3] = N572 & data_mem_write_bank_mask[3];
  assign N572 = data_mem_pkt_yumi_o & N391;
  assign data_mem_fast_read[3] = do_recover | N575;
  assign N575 = N573 & N574;
  assign N573 = yumi_o & decode_lo_fetch_op_;
  assign N574 = N558 | data_mem_bypass_select[3];
  assign data_mem_v_li[3] = N576 | data_mem_slow_write[3];
  assign N576 = data_mem_fast_read[3] | data_mem_slow_read[3];
  assign N281 = ~data_mem_fast_read[3];
  assign data_mem_slow_read[4] = data_mem_pkt_yumi_o & N393;
  assign data_mem_slow_write[4] = N577 & data_mem_write_bank_mask[4];
  assign N577 = data_mem_pkt_yumi_o & N395;
  assign data_mem_fast_read[4] = do_recover | N580;
  assign N580 = N578 & N579;
  assign N578 = yumi_o & decode_lo_fetch_op_;
  assign N579 = N558 | data_mem_bypass_select[4];
  assign data_mem_v_li[4] = N581 | data_mem_slow_write[4];
  assign N581 = data_mem_fast_read[4] | data_mem_slow_read[4];
  assign N291 = ~data_mem_fast_read[4];
  assign data_mem_slow_read[5] = data_mem_pkt_yumi_o & N397;
  assign data_mem_slow_write[5] = N582 & data_mem_write_bank_mask[5];
  assign N582 = data_mem_pkt_yumi_o & N399;
  assign data_mem_fast_read[5] = do_recover | N585;
  assign N585 = N583 & N584;
  assign N583 = yumi_o & decode_lo_fetch_op_;
  assign N584 = N558 | data_mem_bypass_select[5];
  assign data_mem_v_li[5] = N586 | data_mem_slow_write[5];
  assign N586 = data_mem_fast_read[5] | data_mem_slow_read[5];
  assign N301 = ~data_mem_fast_read[5];
  assign data_mem_slow_read[6] = data_mem_pkt_yumi_o & N401;
  assign data_mem_slow_write[6] = N587 & data_mem_write_bank_mask[6];
  assign N587 = data_mem_pkt_yumi_o & N403;
  assign data_mem_fast_read[6] = do_recover | N590;
  assign N590 = N588 & N589;
  assign N588 = yumi_o & decode_lo_fetch_op_;
  assign N589 = N558 | data_mem_bypass_select[6];
  assign data_mem_v_li[6] = N591 | data_mem_slow_write[6];
  assign N591 = data_mem_fast_read[6] | data_mem_slow_read[6];
  assign N311 = ~data_mem_fast_read[6];
  assign data_mem_slow_read[7] = data_mem_pkt_yumi_o & N405;
  assign data_mem_slow_write[7] = N592 & data_mem_write_bank_mask[7];
  assign N592 = data_mem_pkt_yumi_o & N407;
  assign data_mem_fast_read[7] = do_recover | N595;
  assign N595 = N593 & N594;
  assign N593 = yumi_o & decode_lo_fetch_op_;
  assign N594 = N558 | data_mem_bypass_select[7];
  assign data_mem_v_li[7] = N596 | data_mem_slow_write[7];
  assign N596 = data_mem_fast_read[7] | data_mem_slow_read[7];
  assign N321 = ~data_mem_fast_read[7];
  assign N331 = data_mem_pkt_v_i & N604;
  assign N604 = ~N603;
  assign N603 = N602 | data_mem_fast_read[0];
  assign N602 = N601 | data_mem_fast_read[1];
  assign N601 = N600 | data_mem_fast_read[2];
  assign N600 = N599 | data_mem_fast_read[3];
  assign N599 = N598 | data_mem_fast_read[4];
  assign N598 = N597 | data_mem_fast_read[5];
  assign N597 = data_mem_fast_read[7] | data_mem_fast_read[6];
  assign stat_mem_fast_read = N605 & cache_req_yumi_i;
  assign N605 = ~snoop_uncached;
  assign stat_mem_fast_write = N606 & yumi_i;
  assign N606 = ~snoop_uncached;
  assign stat_mem_slow_write = stat_mem_pkt_v_i & N409;
  assign stat_mem_pkt_yumi_o = N608 & N609;
  assign N608 = stat_mem_pkt_v_i & N607;
  assign N607 = ~stat_mem_fast_write;
  assign N609 = ~stat_mem_fast_read;
  assign stat_mem_v_li = N610 | stat_mem_pkt_yumi_o;
  assign N610 = stat_mem_fast_read | stat_mem_fast_write;
  assign stat_mem_w_li = stat_mem_fast_write | N611;
  assign N611 = stat_mem_pkt_yumi_o & stat_mem_slow_write;
  assign N332 = stat_mem_fast_write | stat_mem_fast_read;
  assign N333 = ~N332;
  assign pseudo_hit[7] = N341 | N349;
  assign pseudo_hit[6] = N340 | N348;
  assign pseudo_hit[5] = N339 | N347;
  assign pseudo_hit[4] = N338 | N346;
  assign pseudo_hit[3] = N337 | N345;
  assign pseudo_hit[2] = N336 | N344;
  assign pseudo_hit[1] = N335 | N343;
  assign pseudo_hit[0] = N334 | N342;
  assign N350 = N410 & N416;
  assign N351 = N129 & N350;
  assign N352 = ~N351;

  always @(posedge clk_i) begin
    if(reset_i) begin
      state_r_1_sv2v_reg <= 1'b0;
      state_r_0_sv2v_reg <= 1'b0;
    end else if(N352) begin
      state_r_1_sv2v_reg <= state_n[1];
      state_r_0_sv2v_reg <= state_n[0];
    end 
  end


endmodule



module bsg_dff_reset_en_00000038
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [55:0] data_i;
  output [55:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [55:0] data_o;
  wire N0,N1,N2;
  reg data_o_55_sv2v_reg,data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,
  data_o_51_sv2v_reg,data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,
  data_o_47_sv2v_reg,data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,
  data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,
  data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,
  data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,
  data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,
  data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,
  data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,
  data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,
  data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_55_sv2v_reg <= 1'b0;
      data_o_54_sv2v_reg <= 1'b0;
      data_o_53_sv2v_reg <= 1'b0;
      data_o_52_sv2v_reg <= 1'b0;
      data_o_51_sv2v_reg <= 1'b0;
      data_o_50_sv2v_reg <= 1'b0;
      data_o_49_sv2v_reg <= 1'b0;
      data_o_48_sv2v_reg <= 1'b0;
      data_o_47_sv2v_reg <= 1'b0;
      data_o_46_sv2v_reg <= 1'b0;
      data_o_45_sv2v_reg <= 1'b0;
      data_o_44_sv2v_reg <= 1'b0;
      data_o_43_sv2v_reg <= 1'b0;
      data_o_42_sv2v_reg <= 1'b0;
      data_o_41_sv2v_reg <= 1'b0;
      data_o_40_sv2v_reg <= 1'b0;
      data_o_39_sv2v_reg <= 1'b0;
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bp_fe_realigner_00
(
  clk_i,
  reset_i,
  if2_hit_v_i,
  if2_miss_v_i,
  if2_pc_i,
  if2_data_i,
  if2_br_metadata_fwd_i,
  if2_yumi_o,
  redirect_v_i,
  redirect_pc_i,
  redirect_instr_i,
  redirect_br_metadata_fwd_i,
  redirect_resume_i,
  assembled_v_o,
  assembled_pc_o,
  assembled_instr_o,
  assembled_br_metadata_fwd_o,
  assembled_count_o,
  assembled_partial_o,
  assembled_count_i,
  assembled_yumi_i
);

  input [38:0] if2_pc_i;
  input [63:0] if2_data_i;
  input [48:0] if2_br_metadata_fwd_i;
  input [38:0] redirect_pc_i;
  input [15:0] redirect_instr_i;
  input [48:0] redirect_br_metadata_fwd_i;
  output [38:0] assembled_pc_o;
  output [79:0] assembled_instr_o;
  output [48:0] assembled_br_metadata_fwd_o;
  output [2:0] assembled_count_o;
  input [2:0] assembled_count_i;
  input clk_i;
  input reset_i;
  input if2_hit_v_i;
  input if2_miss_v_i;
  input redirect_v_i;
  input redirect_resume_i;
  input assembled_yumi_i;
  output if2_yumi_o;
  output assembled_v_o;
  output assembled_partial_o;
  wire [38:0] assembled_pc_o,partial_pc_n,realigned_pc;
  wire [79:0] assembled_instr_o;
  wire [48:0] assembled_br_metadata_fwd_o;
  wire [2:0] assembled_count_o,if2_count;
  wire if2_yumi_o,assembled_v_o,assembled_partial_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,
  partial_w_v,partial_v_n,realigned_instr_0__15_,realigned_instr_0__14_,
  realigned_instr_0__13_,realigned_instr_0__12_,realigned_instr_0__11_,realigned_instr_0__10_,
  realigned_instr_0__9_,realigned_instr_0__8_,realigned_instr_0__7_,
  realigned_instr_0__6_,realigned_instr_0__5_,realigned_instr_0__4_,realigned_instr_0__3_,
  realigned_instr_0__2_,realigned_instr_0__1_,realigned_instr_0__0_,N9,N10,N11,partial_store,
  N12,N13,N14,partial_drain,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,
  N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,
  N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,
  N68;
  wire [63:0] if2_instr;
  wire [15:0] partial_instr_n;
  wire [2:2] realigned_count;
  assign assembled_br_metadata_fwd_o[48] = if2_br_metadata_fwd_i[48];
  assign assembled_br_metadata_fwd_o[47] = if2_br_metadata_fwd_i[47];
  assign assembled_br_metadata_fwd_o[46] = if2_br_metadata_fwd_i[46];
  assign assembled_br_metadata_fwd_o[45] = if2_br_metadata_fwd_i[45];
  assign assembled_br_metadata_fwd_o[44] = if2_br_metadata_fwd_i[44];
  assign assembled_br_metadata_fwd_o[43] = if2_br_metadata_fwd_i[43];
  assign assembled_br_metadata_fwd_o[42] = if2_br_metadata_fwd_i[42];
  assign assembled_br_metadata_fwd_o[41] = if2_br_metadata_fwd_i[41];
  assign assembled_br_metadata_fwd_o[40] = if2_br_metadata_fwd_i[40];
  assign assembled_br_metadata_fwd_o[39] = if2_br_metadata_fwd_i[39];
  assign assembled_br_metadata_fwd_o[38] = if2_br_metadata_fwd_i[38];
  assign assembled_br_metadata_fwd_o[37] = if2_br_metadata_fwd_i[37];
  assign assembled_br_metadata_fwd_o[36] = if2_br_metadata_fwd_i[36];
  assign assembled_br_metadata_fwd_o[35] = if2_br_metadata_fwd_i[35];
  assign assembled_br_metadata_fwd_o[34] = if2_br_metadata_fwd_i[34];
  assign assembled_br_metadata_fwd_o[33] = if2_br_metadata_fwd_i[33];
  assign assembled_br_metadata_fwd_o[32] = if2_br_metadata_fwd_i[32];
  assign assembled_br_metadata_fwd_o[31] = if2_br_metadata_fwd_i[31];
  assign assembled_br_metadata_fwd_o[30] = if2_br_metadata_fwd_i[30];
  assign assembled_br_metadata_fwd_o[29] = if2_br_metadata_fwd_i[29];
  assign assembled_br_metadata_fwd_o[28] = if2_br_metadata_fwd_i[28];
  assign assembled_br_metadata_fwd_o[27] = if2_br_metadata_fwd_i[27];
  assign assembled_br_metadata_fwd_o[26] = if2_br_metadata_fwd_i[26];
  assign assembled_br_metadata_fwd_o[25] = if2_br_metadata_fwd_i[25];
  assign assembled_br_metadata_fwd_o[24] = if2_br_metadata_fwd_i[24];
  assign assembled_br_metadata_fwd_o[23] = if2_br_metadata_fwd_i[23];
  assign assembled_br_metadata_fwd_o[22] = if2_br_metadata_fwd_i[22];
  assign assembled_br_metadata_fwd_o[21] = if2_br_metadata_fwd_i[21];
  assign assembled_br_metadata_fwd_o[20] = if2_br_metadata_fwd_i[20];
  assign assembled_br_metadata_fwd_o[19] = if2_br_metadata_fwd_i[19];
  assign assembled_br_metadata_fwd_o[18] = if2_br_metadata_fwd_i[18];
  assign assembled_br_metadata_fwd_o[17] = if2_br_metadata_fwd_i[17];
  assign assembled_br_metadata_fwd_o[16] = if2_br_metadata_fwd_i[16];
  assign assembled_br_metadata_fwd_o[15] = if2_br_metadata_fwd_i[15];
  assign assembled_br_metadata_fwd_o[14] = if2_br_metadata_fwd_i[14];
  assign assembled_br_metadata_fwd_o[13] = if2_br_metadata_fwd_i[13];
  assign assembled_br_metadata_fwd_o[12] = if2_br_metadata_fwd_i[12];
  assign assembled_br_metadata_fwd_o[11] = if2_br_metadata_fwd_i[11];
  assign assembled_br_metadata_fwd_o[10] = if2_br_metadata_fwd_i[10];
  assign assembled_br_metadata_fwd_o[9] = if2_br_metadata_fwd_i[9];
  assign assembled_br_metadata_fwd_o[8] = if2_br_metadata_fwd_i[8];
  assign assembled_br_metadata_fwd_o[7] = if2_br_metadata_fwd_i[7];
  assign assembled_br_metadata_fwd_o[6] = if2_br_metadata_fwd_i[6];
  assign assembled_br_metadata_fwd_o[5] = if2_br_metadata_fwd_i[5];
  assign assembled_br_metadata_fwd_o[4] = if2_br_metadata_fwd_i[4];
  assign assembled_br_metadata_fwd_o[3] = if2_br_metadata_fwd_i[3];
  assign assembled_br_metadata_fwd_o[2] = if2_br_metadata_fwd_i[2];
  assign assembled_br_metadata_fwd_o[1] = if2_br_metadata_fwd_i[1];
  assign assembled_br_metadata_fwd_o[0] = if2_br_metadata_fwd_i[0];

  bsg_dff_reset_en_00000038
  partial_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(partial_w_v),
    .data_i({ partial_instr_n, partial_pc_n, partial_v_n }),
    .data_o({ realigned_instr_0__15_, realigned_instr_0__14_, realigned_instr_0__13_, realigned_instr_0__12_, realigned_instr_0__11_, realigned_instr_0__10_, realigned_instr_0__9_, realigned_instr_0__8_, realigned_instr_0__7_, realigned_instr_0__6_, realigned_instr_0__5_, realigned_instr_0__4_, realigned_instr_0__3_, realigned_instr_0__2_, realigned_instr_0__1_, realigned_instr_0__0_, realigned_pc, assembled_partial_o })
  );

  assign partial_store = { N11, N10, N9 } == 1'b1;
  assign partial_drain = { N14, N13, N12 } > 1'b1;
  assign if2_instr = if2_data_i >> { if2_pc_i[2:1], 1'b0, 1'b0, 1'b0, 1'b0 };
  assign { N8, N7, N6 } = { 1'b1, 1'b0, 1'b0 } - if2_pc_i[2:1];
  assign { N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22 } = assembled_pc_o + { assembled_count_i, 1'b0 };
  assign { N11, N10, N9 } = assembled_count_o - assembled_count_i;
  assign { N14, N13, N12 } = assembled_count_o - assembled_count_i;
  assign if2_count = (N0)? { N8, N7, N6 } : 
                     (N1)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = if2_hit_v_i;
  assign N1 = N5;
  assign partial_v_n = (N2)? redirect_resume_i : 
                       (N18)? partial_store : 
                       (N16)? assembled_partial_o : 1'b0;
  assign N2 = redirect_v_i;
  assign partial_pc_n = (N2)? redirect_pc_i : 
                        (N61)? { N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22 } : 
                        (N20)? if2_pc_i : 1'b0;
  assign partial_instr_n = (N2)? redirect_instr_i : 
                           (N64)? if2_data_i[63:48] : 
                           (N63)? if2_data_i[63:48] : 1'b0;
  assign assembled_pc_o = (N3)? realigned_pc : 
                          (N4)? if2_pc_i : 1'b0;
  assign N3 = assembled_partial_o;
  assign N4 = N65;
  assign assembled_instr_o = (N3)? { if2_data_i, realigned_instr_0__15_, realigned_instr_0__14_, realigned_instr_0__13_, realigned_instr_0__12_, realigned_instr_0__11_, realigned_instr_0__10_, realigned_instr_0__9_, realigned_instr_0__8_, realigned_instr_0__7_, realigned_instr_0__6_, realigned_instr_0__5_, realigned_instr_0__4_, realigned_instr_0__3_, realigned_instr_0__2_, realigned_instr_0__1_, realigned_instr_0__0_ } : 
                             (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, if2_instr } : 1'b0;
  assign assembled_count_o = (N3)? { realigned_count[2:2], 1'b0, 1'b1 } : 
                             (N4)? if2_count : 1'b0;
  assign N5 = ~if2_hit_v_i;
  assign realigned_count[2] = if2_hit_v_i;
  assign partial_w_v = N66 | if2_yumi_o;
  assign N66 = redirect_v_i | assembled_yumi_i;
  assign N15 = assembled_yumi_i | redirect_v_i;
  assign N16 = ~N15;
  assign N17 = ~redirect_v_i;
  assign N18 = assembled_yumi_i & N17;
  assign N19 = assembled_yumi_i | redirect_v_i;
  assign N20 = ~N19;
  assign N21 = N61;
  assign N61 = assembled_yumi_i & N17;
  assign N62 = assembled_yumi_i | redirect_v_i;
  assign N63 = ~N62;
  assign N64 = assembled_yumi_i & N17;
  assign N65 = ~assembled_partial_o;
  assign assembled_v_o = if2_hit_v_i | if2_miss_v_i;
  assign if2_yumi_o = N68 & assembled_yumi_i;
  assign N68 = if2_hit_v_i & N67;
  assign N67 = ~partial_drain;

endmodule



module bsg_scan_00000005_1_0
(
  i,
  o
);

  input [4:0] i;
  output [4:0] o;
  wire [4:0] o;
  wire t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__4_ = i[4] | 1'b0;
  assign t_1__3_ = i[3] | i[4];
  assign t_1__2_ = i[2] | i[3];
  assign t_1__1_ = i[1] | i[2];
  assign t_1__0_ = i[0] | i[1];
  assign t_2__4_ = t_1__4_ | 1'b0;
  assign t_2__3_ = t_1__3_ | 1'b0;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign o[4] = t_2__4_ | 1'b0;
  assign o[3] = t_2__3_ | 1'b0;
  assign o[2] = t_2__2_ | 1'b0;
  assign o[1] = t_2__1_ | 1'b0;
  assign o[0] = t_2__0_ | t_2__4_;

endmodule



module bsg_priority_encode_one_hot_out_00000005_0
(
  i,
  o,
  v_o
);

  input [4:0] i;
  output [4:0] o;
  output v_o;
  wire [4:0] o;
  wire v_o,N0,N1,N2,N3;
  wire [3:1] scan_lo;

  bsg_scan_00000005_1_0
  \nw1.scan 
  (
    .i(i),
    .o({ o[4:4], scan_lo, v_o })
  );

  assign o[3] = scan_lo[3] & N0;
  assign N0 = ~o[4];
  assign o[2] = scan_lo[2] & N1;
  assign N1 = ~scan_lo[3];
  assign o[1] = scan_lo[1] & N2;
  assign N2 = ~scan_lo[2];
  assign o[0] = v_o & N3;
  assign N3 = ~scan_lo[1];

endmodule



module bsg_encode_one_hot_00000005_0
(
  i,
  addr_o,
  v_o
);

  input [4:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o,v_2__4_,v_1__6_,v_1__4_,v_1__2_,v_1__0_,addr_2__4_,addr_2__0_;
  assign v_1__0_ = 1'b0 | 1'b0;
  assign v_1__2_ = i[0] | 1'b0;
  assign v_1__4_ = i[2] | i[1];
  assign v_1__6_ = i[4] | i[3];
  assign addr_o[2] = v_1__2_ | v_1__0_;
  assign addr_2__0_ = 1'b0 | 1'b0;
  assign v_2__4_ = v_1__6_ | v_1__4_;
  assign addr_2__4_ = i[1] | i[3];
  assign v_o = v_2__4_ | addr_o[2];
  assign addr_o[1] = v_1__0_ | v_1__4_;
  assign addr_o[0] = addr_2__0_ | addr_2__4_;

endmodule



module bsg_priority_encode_00000005_0
(
  i,
  addr_o,
  v_o
);

  input [4:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [4:0] enc_lo;

  bsg_priority_encode_one_hot_out_00000005_0
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_00000005_0
  b
  (
    .i(enc_lo),
    .addr_o(addr_o)
  );


endmodule



module bsg_scan_00000005_1_1
(
  i,
  o
);

  input [4:0] i;
  output [4:0] o;
  wire [4:0] o;
  wire t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__4_ = i[0] | 1'b0;
  assign t_1__3_ = i[1] | i[0];
  assign t_1__2_ = i[2] | i[1];
  assign t_1__1_ = i[3] | i[2];
  assign t_1__0_ = i[4] | i[3];
  assign t_2__4_ = t_1__4_ | 1'b0;
  assign t_2__3_ = t_1__3_ | 1'b0;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign o[0] = t_2__4_ | 1'b0;
  assign o[1] = t_2__3_ | 1'b0;
  assign o[2] = t_2__2_ | 1'b0;
  assign o[3] = t_2__1_ | 1'b0;
  assign o[4] = t_2__0_ | t_2__4_;

endmodule



module bsg_priority_encode_one_hot_out_00000005_1
(
  i,
  o,
  v_o
);

  input [4:0] i;
  output [4:0] o;
  output v_o;
  wire [4:0] o;
  wire v_o,N0,N1,N2,N3;
  wire [3:1] scan_lo;

  bsg_scan_00000005_1_1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, scan_lo, o[0:0] })
  );

  assign o[4] = v_o & N0;
  assign N0 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N1;
  assign N1 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N2;
  assign N2 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N3;
  assign N3 = ~o[0];

endmodule



module bsg_encode_one_hot_00000005_1
(
  i,
  addr_o,
  v_o
);

  input [4:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o,v_2__0_,v_1__6_,v_1__4_,v_1__2_,v_1__0_,addr_2__4_,addr_2__0_;
  assign v_1__0_ = i[1] | i[0];
  assign v_1__2_ = i[3] | i[2];
  assign v_1__4_ = 1'b0 | i[4];
  assign v_1__6_ = 1'b0 | 1'b0;
  assign v_2__0_ = v_1__2_ | v_1__0_;
  assign addr_2__0_ = i[1] | i[3];
  assign addr_o[2] = v_1__6_ | v_1__4_;
  assign addr_2__4_ = 1'b0 | 1'b0;
  assign v_o = addr_o[2] | v_2__0_;
  assign addr_o[1] = v_1__2_ | v_1__6_;
  assign addr_o[0] = addr_2__0_ | addr_2__4_;

endmodule



module bsg_priority_encode_00000005_1
(
  i,
  addr_o,
  v_o
);

  input [4:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [4:0] enc_lo;

  bsg_priority_encode_one_hot_out_00000005_1
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_00000005_1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o)
  );


endmodule



module bsg_scan_00000006_1_0
(
  i,
  o
);

  input [5:0] i;
  output [5:0] o;
  wire [5:0] o;
  wire t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,
  t_1__1_,t_1__0_;
  assign t_1__5_ = i[5] | 1'b0;
  assign t_1__4_ = i[4] | i[5];
  assign t_1__3_ = i[3] | i[4];
  assign t_1__2_ = i[2] | i[3];
  assign t_1__1_ = i[1] | i[2];
  assign t_1__0_ = i[0] | i[1];
  assign t_2__5_ = t_1__5_ | 1'b0;
  assign t_2__4_ = t_1__4_ | 1'b0;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign o[5] = t_2__5_ | 1'b0;
  assign o[4] = t_2__4_ | 1'b0;
  assign o[3] = t_2__3_ | 1'b0;
  assign o[2] = t_2__2_ | 1'b0;
  assign o[1] = t_2__1_ | t_2__5_;
  assign o[0] = t_2__0_ | t_2__4_;

endmodule



module bsg_priority_encode_one_hot_out_00000006_0
(
  i,
  o,
  v_o
);

  input [5:0] i;
  output [5:0] o;
  output v_o;
  wire [5:0] o;
  wire v_o,N0,N1,N2,N3,N4;
  wire [4:1] scan_lo;

  bsg_scan_00000006_1_0
  \nw1.scan 
  (
    .i(i),
    .o({ o[5:5], scan_lo, v_o })
  );

  assign o[4] = scan_lo[4] & N0;
  assign N0 = ~o[5];
  assign o[3] = scan_lo[3] & N1;
  assign N1 = ~scan_lo[4];
  assign o[2] = scan_lo[2] & N2;
  assign N2 = ~scan_lo[3];
  assign o[1] = scan_lo[1] & N3;
  assign N3 = ~scan_lo[2];
  assign o[0] = v_o & N4;
  assign N4 = ~scan_lo[1];

endmodule



module bsg_encode_one_hot_00000006_0
(
  i,
  addr_o,
  v_o
);

  input [5:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o,v_2__4_,v_1__6_,v_1__4_,v_1__2_,v_1__0_,addr_2__4_,addr_2__0_;
  assign v_1__0_ = 1'b0 | 1'b0;
  assign v_1__2_ = i[1] | i[0];
  assign v_1__4_ = i[3] | i[2];
  assign v_1__6_ = i[5] | i[4];
  assign addr_o[2] = v_1__2_ | v_1__0_;
  assign addr_2__0_ = 1'b0 | i[0];
  assign v_2__4_ = v_1__6_ | v_1__4_;
  assign addr_2__4_ = i[2] | i[4];
  assign v_o = v_2__4_ | addr_o[2];
  assign addr_o[1] = v_1__0_ | v_1__4_;
  assign addr_o[0] = addr_2__0_ | addr_2__4_;

endmodule



module bsg_priority_encode_00000006_0
(
  i,
  addr_o,
  v_o
);

  input [5:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [5:0] enc_lo;

  bsg_priority_encode_one_hot_out_00000006_0
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_00000006_0
  b
  (
    .i(enc_lo),
    .addr_o(addr_o)
  );


endmodule



module bsg_mux_47_00000006
(
  data_i,
  sel_i,
  data_o
);

  input [281:0] data_i;
  input [2:0] sel_i;
  output [46:0] data_o;
  wire [46:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;
  assign N13 = N0 & N1 & N2;
  assign N0 = ~sel_i[2];
  assign N1 = ~sel_i[0];
  assign N2 = ~sel_i[1];
  assign N14 = sel_i[2] & N3;
  assign N3 = ~sel_i[0];
  assign N15 = N4 & sel_i[0] & N5;
  assign N4 = ~sel_i[2];
  assign N5 = ~sel_i[1];
  assign N17 = N6 & sel_i[1];
  assign N6 = ~sel_i[0];
  assign N18 = sel_i[0] & sel_i[1];
  assign N16 = sel_i[2] & sel_i[0];
  assign data_o[46] = (N7)? data_i[46] : 
                      (N8)? data_i[93] : 
                      (N9)? data_i[140] : 
                      (N10)? data_i[187] : 
                      (N11)? data_i[234] : 
                      (N12)? data_i[281] : 1'b0;
  assign N7 = N13;
  assign N8 = N15;
  assign N9 = N17;
  assign N10 = N18;
  assign N11 = N14;
  assign N12 = N16;
  assign data_o[45] = (N7)? data_i[45] : 
                      (N8)? data_i[92] : 
                      (N9)? data_i[139] : 
                      (N10)? data_i[186] : 
                      (N11)? data_i[233] : 
                      (N12)? data_i[280] : 1'b0;
  assign data_o[44] = (N7)? data_i[44] : 
                      (N8)? data_i[91] : 
                      (N9)? data_i[138] : 
                      (N10)? data_i[185] : 
                      (N11)? data_i[232] : 
                      (N12)? data_i[279] : 1'b0;
  assign data_o[43] = (N7)? data_i[43] : 
                      (N8)? data_i[90] : 
                      (N9)? data_i[137] : 
                      (N10)? data_i[184] : 
                      (N11)? data_i[231] : 
                      (N12)? data_i[278] : 1'b0;
  assign data_o[42] = (N7)? data_i[42] : 
                      (N8)? data_i[89] : 
                      (N9)? data_i[136] : 
                      (N10)? data_i[183] : 
                      (N11)? data_i[230] : 
                      (N12)? data_i[277] : 1'b0;
  assign data_o[41] = (N7)? data_i[41] : 
                      (N8)? data_i[88] : 
                      (N9)? data_i[135] : 
                      (N10)? data_i[182] : 
                      (N11)? data_i[229] : 
                      (N12)? data_i[276] : 1'b0;
  assign data_o[40] = (N7)? data_i[40] : 
                      (N8)? data_i[87] : 
                      (N9)? data_i[134] : 
                      (N10)? data_i[181] : 
                      (N11)? data_i[228] : 
                      (N12)? data_i[275] : 1'b0;
  assign data_o[39] = (N7)? data_i[39] : 
                      (N8)? data_i[86] : 
                      (N9)? data_i[133] : 
                      (N10)? data_i[180] : 
                      (N11)? data_i[227] : 
                      (N12)? data_i[274] : 1'b0;
  assign data_o[38] = (N7)? data_i[38] : 
                      (N8)? data_i[85] : 
                      (N9)? data_i[132] : 
                      (N10)? data_i[179] : 
                      (N11)? data_i[226] : 
                      (N12)? data_i[273] : 1'b0;
  assign data_o[37] = (N7)? data_i[37] : 
                      (N8)? data_i[84] : 
                      (N9)? data_i[131] : 
                      (N10)? data_i[178] : 
                      (N11)? data_i[225] : 
                      (N12)? data_i[272] : 1'b0;
  assign data_o[36] = (N7)? data_i[36] : 
                      (N8)? data_i[83] : 
                      (N9)? data_i[130] : 
                      (N10)? data_i[177] : 
                      (N11)? data_i[224] : 
                      (N12)? data_i[271] : 1'b0;
  assign data_o[35] = (N7)? data_i[35] : 
                      (N8)? data_i[82] : 
                      (N9)? data_i[129] : 
                      (N10)? data_i[176] : 
                      (N11)? data_i[223] : 
                      (N12)? data_i[270] : 1'b0;
  assign data_o[34] = (N7)? data_i[34] : 
                      (N8)? data_i[81] : 
                      (N9)? data_i[128] : 
                      (N10)? data_i[175] : 
                      (N11)? data_i[222] : 
                      (N12)? data_i[269] : 1'b0;
  assign data_o[33] = (N7)? data_i[33] : 
                      (N8)? data_i[80] : 
                      (N9)? data_i[127] : 
                      (N10)? data_i[174] : 
                      (N11)? data_i[221] : 
                      (N12)? data_i[268] : 1'b0;
  assign data_o[32] = (N7)? data_i[32] : 
                      (N8)? data_i[79] : 
                      (N9)? data_i[126] : 
                      (N10)? data_i[173] : 
                      (N11)? data_i[220] : 
                      (N12)? data_i[267] : 1'b0;
  assign data_o[31] = (N7)? data_i[31] : 
                      (N8)? data_i[78] : 
                      (N9)? data_i[125] : 
                      (N10)? data_i[172] : 
                      (N11)? data_i[219] : 
                      (N12)? data_i[266] : 1'b0;
  assign data_o[30] = (N7)? data_i[30] : 
                      (N8)? data_i[77] : 
                      (N9)? data_i[124] : 
                      (N10)? data_i[171] : 
                      (N11)? data_i[218] : 
                      (N12)? data_i[265] : 1'b0;
  assign data_o[29] = (N7)? data_i[29] : 
                      (N8)? data_i[76] : 
                      (N9)? data_i[123] : 
                      (N10)? data_i[170] : 
                      (N11)? data_i[217] : 
                      (N12)? data_i[264] : 1'b0;
  assign data_o[28] = (N7)? data_i[28] : 
                      (N8)? data_i[75] : 
                      (N9)? data_i[122] : 
                      (N10)? data_i[169] : 
                      (N11)? data_i[216] : 
                      (N12)? data_i[263] : 1'b0;
  assign data_o[27] = (N7)? data_i[27] : 
                      (N8)? data_i[74] : 
                      (N9)? data_i[121] : 
                      (N10)? data_i[168] : 
                      (N11)? data_i[215] : 
                      (N12)? data_i[262] : 1'b0;
  assign data_o[26] = (N7)? data_i[26] : 
                      (N8)? data_i[73] : 
                      (N9)? data_i[120] : 
                      (N10)? data_i[167] : 
                      (N11)? data_i[214] : 
                      (N12)? data_i[261] : 1'b0;
  assign data_o[25] = (N7)? data_i[25] : 
                      (N8)? data_i[72] : 
                      (N9)? data_i[119] : 
                      (N10)? data_i[166] : 
                      (N11)? data_i[213] : 
                      (N12)? data_i[260] : 1'b0;
  assign data_o[24] = (N7)? data_i[24] : 
                      (N8)? data_i[71] : 
                      (N9)? data_i[118] : 
                      (N10)? data_i[165] : 
                      (N11)? data_i[212] : 
                      (N12)? data_i[259] : 1'b0;
  assign data_o[23] = (N7)? data_i[23] : 
                      (N8)? data_i[70] : 
                      (N9)? data_i[117] : 
                      (N10)? data_i[164] : 
                      (N11)? data_i[211] : 
                      (N12)? data_i[258] : 1'b0;
  assign data_o[22] = (N7)? data_i[22] : 
                      (N8)? data_i[69] : 
                      (N9)? data_i[116] : 
                      (N10)? data_i[163] : 
                      (N11)? data_i[210] : 
                      (N12)? data_i[257] : 1'b0;
  assign data_o[21] = (N7)? data_i[21] : 
                      (N8)? data_i[68] : 
                      (N9)? data_i[115] : 
                      (N10)? data_i[162] : 
                      (N11)? data_i[209] : 
                      (N12)? data_i[256] : 1'b0;
  assign data_o[20] = (N7)? data_i[20] : 
                      (N8)? data_i[67] : 
                      (N9)? data_i[114] : 
                      (N10)? data_i[161] : 
                      (N11)? data_i[208] : 
                      (N12)? data_i[255] : 1'b0;
  assign data_o[19] = (N7)? data_i[19] : 
                      (N8)? data_i[66] : 
                      (N9)? data_i[113] : 
                      (N10)? data_i[160] : 
                      (N11)? data_i[207] : 
                      (N12)? data_i[254] : 1'b0;
  assign data_o[18] = (N7)? data_i[18] : 
                      (N8)? data_i[65] : 
                      (N9)? data_i[112] : 
                      (N10)? data_i[159] : 
                      (N11)? data_i[206] : 
                      (N12)? data_i[253] : 1'b0;
  assign data_o[17] = (N7)? data_i[17] : 
                      (N8)? data_i[64] : 
                      (N9)? data_i[111] : 
                      (N10)? data_i[158] : 
                      (N11)? data_i[205] : 
                      (N12)? data_i[252] : 1'b0;
  assign data_o[16] = (N7)? data_i[16] : 
                      (N8)? data_i[63] : 
                      (N9)? data_i[110] : 
                      (N10)? data_i[157] : 
                      (N11)? data_i[204] : 
                      (N12)? data_i[251] : 1'b0;
  assign data_o[15] = (N7)? data_i[15] : 
                      (N8)? data_i[62] : 
                      (N9)? data_i[109] : 
                      (N10)? data_i[156] : 
                      (N11)? data_i[203] : 
                      (N12)? data_i[250] : 1'b0;
  assign data_o[14] = (N7)? data_i[14] : 
                      (N8)? data_i[61] : 
                      (N9)? data_i[108] : 
                      (N10)? data_i[155] : 
                      (N11)? data_i[202] : 
                      (N12)? data_i[249] : 1'b0;
  assign data_o[13] = (N7)? data_i[13] : 
                      (N8)? data_i[60] : 
                      (N9)? data_i[107] : 
                      (N10)? data_i[154] : 
                      (N11)? data_i[201] : 
                      (N12)? data_i[248] : 1'b0;
  assign data_o[12] = (N7)? data_i[12] : 
                      (N8)? data_i[59] : 
                      (N9)? data_i[106] : 
                      (N10)? data_i[153] : 
                      (N11)? data_i[200] : 
                      (N12)? data_i[247] : 1'b0;
  assign data_o[11] = (N7)? data_i[11] : 
                      (N8)? data_i[58] : 
                      (N9)? data_i[105] : 
                      (N10)? data_i[152] : 
                      (N11)? data_i[199] : 
                      (N12)? data_i[246] : 1'b0;
  assign data_o[10] = (N7)? data_i[10] : 
                      (N8)? data_i[57] : 
                      (N9)? data_i[104] : 
                      (N10)? data_i[151] : 
                      (N11)? data_i[198] : 
                      (N12)? data_i[245] : 1'b0;
  assign data_o[9] = (N7)? data_i[9] : 
                     (N8)? data_i[56] : 
                     (N9)? data_i[103] : 
                     (N10)? data_i[150] : 
                     (N11)? data_i[197] : 
                     (N12)? data_i[244] : 1'b0;
  assign data_o[8] = (N7)? data_i[8] : 
                     (N8)? data_i[55] : 
                     (N9)? data_i[102] : 
                     (N10)? data_i[149] : 
                     (N11)? data_i[196] : 
                     (N12)? data_i[243] : 1'b0;
  assign data_o[7] = (N7)? data_i[7] : 
                     (N8)? data_i[54] : 
                     (N9)? data_i[101] : 
                     (N10)? data_i[148] : 
                     (N11)? data_i[195] : 
                     (N12)? data_i[242] : 1'b0;
  assign data_o[6] = (N7)? data_i[6] : 
                     (N8)? data_i[53] : 
                     (N9)? data_i[100] : 
                     (N10)? data_i[147] : 
                     (N11)? data_i[194] : 
                     (N12)? data_i[241] : 1'b0;
  assign data_o[5] = (N7)? data_i[5] : 
                     (N8)? data_i[52] : 
                     (N9)? data_i[99] : 
                     (N10)? data_i[146] : 
                     (N11)? data_i[193] : 
                     (N12)? data_i[240] : 1'b0;
  assign data_o[4] = (N7)? data_i[4] : 
                     (N8)? data_i[51] : 
                     (N9)? data_i[98] : 
                     (N10)? data_i[145] : 
                     (N11)? data_i[192] : 
                     (N12)? data_i[239] : 1'b0;
  assign data_o[3] = (N7)? data_i[3] : 
                     (N8)? data_i[50] : 
                     (N9)? data_i[97] : 
                     (N10)? data_i[144] : 
                     (N11)? data_i[191] : 
                     (N12)? data_i[238] : 1'b0;
  assign data_o[2] = (N7)? data_i[2] : 
                     (N8)? data_i[49] : 
                     (N9)? data_i[96] : 
                     (N10)? data_i[143] : 
                     (N11)? data_i[190] : 
                     (N12)? data_i[237] : 1'b0;
  assign data_o[1] = (N7)? data_i[1] : 
                     (N8)? data_i[48] : 
                     (N9)? data_i[95] : 
                     (N10)? data_i[142] : 
                     (N11)? data_i[189] : 
                     (N12)? data_i[236] : 1'b0;
  assign data_o[0] = (N7)? data_i[0] : 
                     (N8)? data_i[47] : 
                     (N9)? data_i[94] : 
                     (N10)? data_i[141] : 
                     (N11)? data_i[188] : 
                     (N12)? data_i[235] : 1'b0;

endmodule



module bp_fe_scan_00
(
  assembled_v_i,
  assembled_pc_i,
  assembled_instr_i,
  assembled_br_metadata_fwd_i,
  assembled_count_i,
  assembled_partial_i,
  assembled_count_o,
  assembled_yumi_o,
  fetch_v_o,
  fetch_pc_o,
  fetch_instr_o,
  fetch_br_metadata_fwd_o,
  fetch_count_o,
  fetch_partial_o,
  fetch_scan_o,
  fetch_startup_o,
  fetch_catchup_o,
  fetch_rebase_o,
  fetch_linear_o,
  fetch_taken_i,
  fetch_yumi_i
);

  input [38:0] assembled_pc_i;
  input [79:0] assembled_instr_i;
  input [48:0] assembled_br_metadata_fwd_i;
  input [2:0] assembled_count_i;
  output [2:0] assembled_count_o;
  output [38:0] fetch_pc_o;
  output [79:0] fetch_instr_o;
  output [48:0] fetch_br_metadata_fwd_o;
  output [2:0] fetch_count_o;
  output [124:0] fetch_scan_o;
  input assembled_v_i;
  input assembled_partial_i;
  input fetch_taken_i;
  input fetch_yumi_i;
  output assembled_yumi_o;
  output fetch_v_o;
  output fetch_partial_o;
  output fetch_startup_o;
  output fetch_catchup_o;
  output fetch_rebase_o;
  output fetch_linear_o;
  wire [2:0] assembled_count_o,fetch_count_o,complete_addr,linear_sel,linear_count,
  branch_sel,branch_count,last_branch_addr,last_branch_sel,next_sel;
  wire [38:0] fetch_pc_o,\scan_0_.imm ,\scan_1_.imm ,\scan_2_.imm ,\scan_3_.imm ,
  \scan_4_.imm ,\scan_5_.imm ;
  wire [79:0] fetch_instr_o;
  wire [48:0] fetch_br_metadata_fwd_o;
  wire [124:0] fetch_scan_o;
  wire assembled_yumi_o,fetch_v_o,fetch_partial_o,fetch_startup_o,fetch_catchup_o,
  fetch_rebase_o,fetch_linear_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,
  N16,N17,N18,N19,N20,N21,N22,N23,N24,full1_5_,full1_4_,full1_3_,full1_2_,full1_1_,
  full1_0_,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  \scan_0_.is_br ,N39,N40,N41,N42,N43,N44,N45,N46,N47,\scan_0_.is_jal ,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,\scan_0_.is_jalr ,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,
  \scan_0_.is_link_dest ,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  \scan_0_.is_link_src ,N82,\scan_0_.is_link_match ,\scan_0_.is_call ,\scan_0_.is_return ,
  N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,\scan_0_.is_cbr ,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,
  N147,N148,\scan_0_.is_cj ,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,
  N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,
  \scan_0_.is_cjr ,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,
  N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,
  \scan_0_.is_cjalr ,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  \scan_0_.is_clink_src ,\scan_0_.is_clink_match ,\scan_0_.is_ccall ,\scan_0_.is_creturn ,N214,
  N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,
  N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,
  N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,
  N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,
  N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,
  N295,N296,N297,N298,N299,N300,decode_lo_5__br_,decode_lo_5__jal_,
  decode_lo_5__jalr_,decode_lo_5__call_,decode_lo_5___return_,decode_lo_5__full1_,
  decode_lo_5__full2_,decode_lo_5__comp_,decode_lo_4__br_,decode_lo_4__jal_,decode_lo_4__jalr_,
  decode_lo_4__call_,decode_lo_4___return_,decode_lo_4__full1_,decode_lo_4__full2_,
  decode_lo_4__comp_,decode_lo_3__br_,decode_lo_3__jal_,decode_lo_3__jalr_,
  decode_lo_3__call_,decode_lo_3___return_,decode_lo_3__full1_,decode_lo_3__full2_,
  decode_lo_3__comp_,decode_lo_2__br_,decode_lo_2__jal_,decode_lo_2__jalr_,
  decode_lo_2__call_,decode_lo_2___return_,decode_lo_2__full1_,decode_lo_2__full2_,
  decode_lo_2__comp_,decode_lo_1__br_,decode_lo_1__jal_,decode_lo_1__jalr_,decode_lo_1__call_,
  decode_lo_1___return_,decode_lo_1__full1_,decode_lo_1__full2_,decode_lo_1__comp_,
  decode_lo_0__br_,decode_lo_0__jal_,decode_lo_0__jalr_,decode_lo_0__call_,
  decode_lo_0___return_,decode_lo_0__full1_,decode_lo_0__full2_,decode_lo_0__comp_,N301,
  N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,\scan_1_.is_br ,
  N315,N316,N317,N318,N319,N320,N321,N322,N323,\scan_1_.is_jal ,N324,N325,N326,
  N327,N328,N329,N330,N331,N332,N333,\scan_1_.is_jalr ,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,\scan_1_.is_link_dest ,N346,N347,N348,N349,N350,
  N351,N352,N353,N354,N355,N356,N357,\scan_1_.is_link_src ,N358,
  \scan_1_.is_link_match ,\scan_1_.is_call ,\scan_1_.is_return ,N359,N360,N361,N362,N363,N364,N365,
  N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,
  N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,
  N398,N399,N400,N401,N402,N403,\scan_1_.is_cbr ,N404,N405,N406,N407,N408,N409,N410,
  N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,
  \scan_1_.is_cj ,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,
  N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,\scan_1_.is_cjr ,
  N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,
  N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,\scan_1_.is_cjalr ,N480,
  N481,N482,N483,N484,N485,N486,N487,N488,N489,\scan_1_.is_clink_src ,
  \scan_1_.is_clink_match ,\scan_1_.is_ccall ,\scan_1_.is_creturn ,N490,N491,N492,N493,N494,
  N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,
  N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,
  N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,
  N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,
  N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,
  N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,
  \scan_2_.is_br ,N591,N592,N593,N594,N595,N596,N597,N598,N599,\scan_2_.is_jal ,
  N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,\scan_2_.is_jalr ,N610,N611,N612,
  N613,N614,N615,N616,N617,N618,N619,N620,N621,\scan_2_.is_link_dest ,N622,N623,
  N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,\scan_2_.is_link_src ,N634,
  \scan_2_.is_link_match ,\scan_2_.is_call ,\scan_2_.is_return ,N635,N636,N637,N638,
  N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,
  N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,
  N671,N672,N673,N674,N675,N676,N677,N678,N679,\scan_2_.is_cbr ,N680,N681,N682,N683,
  N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,
  N700,\scan_2_.is_cj ,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,
  N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,
  \scan_2_.is_cjr ,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,
  N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,
  \scan_2_.is_cjalr ,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,
  \scan_2_.is_clink_src ,\scan_2_.is_clink_match ,\scan_2_.is_ccall ,\scan_2_.is_creturn ,N766,N767,
  N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,
  N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,
  N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,
  N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,
  N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,
  N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,
  N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,
  N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,
  N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,
  N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,
  N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,
  N944,N945,\scan_3_.is_br ,N946,N947,N948,N949,N950,N951,N952,N953,N954,
  \scan_3_.is_jal ,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,\scan_3_.is_jalr ,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,\scan_3_.is_link_dest ,
  N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,\scan_3_.is_link_src ,
  N989,\scan_3_.is_link_match ,\scan_3_.is_call ,\scan_3_.is_return ,N990,N991,
  N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,
  N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,
  N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,
  N1034,\scan_3_.is_cbr ,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,
  N1044,N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,
  \scan_3_.is_cj ,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,
  N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,
  N1081,N1082,\scan_3_.is_cjr ,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091,
  N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,\scan_3_.is_cjalr ,N1111,N1112,N1113,N1114,
  N1115,N1116,N1117,N1118,N1119,N1120,\scan_3_.is_clink_src ,\scan_3_.is_clink_match ,
  \scan_3_.is_ccall ,\scan_3_.is_creturn ,N1121,N1122,N1123,N1124,N1125,N1126,
  N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,
  N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,
  N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,
  N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,
  N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,
  N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,
  N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,
  N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,
  N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,
  N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,
  N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,
  N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,
  N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,
  \scan_4_.is_br ,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,
  \scan_4_.is_jal ,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,N1318,N1319,
  \scan_4_.is_jalr ,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,N1331,
  \scan_4_.is_link_dest ,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,
  N1342,N1343,\scan_4_.is_link_src ,N1344,\scan_4_.is_link_match ,
  \scan_4_.is_call ,\scan_4_.is_return ,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,
  N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,
  N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,
  N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,\scan_4_.is_cbr ,N1390,N1391,
  N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,
  N1405,N1406,N1407,N1408,N1409,N1410,\scan_4_.is_cj ,N1411,N1412,N1413,N1414,N1415,
  N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,
  N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,\scan_4_.is_cjr ,N1438,
  N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,N1451,N1452,
  N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,N1465,
  \scan_4_.is_cjalr ,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,
  \scan_4_.is_clink_src ,\scan_4_.is_clink_match ,\scan_4_.is_ccall ,
  \scan_4_.is_creturn ,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,
  N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,
  N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,
  N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,
  N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,
  N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,
  N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,
  N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,
  N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,
  N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,
  N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,
  N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,
  N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,
  \scan_5_.curr_instr_rs1_addr__0_ ,\scan_5_.curr_instr_funct3__2_ ,\scan_5_.curr_instr_funct3__1_ ,
  \scan_5_.curr_instr_funct3__0_ ,\scan_5_.curr_instr_rd_addr__4_ ,
  \scan_5_.curr_instr_rd_addr__3_ ,\scan_5_.curr_instr_rd_addr__2_ ,\scan_5_.curr_instr_rd_addr__1_ ,
  \scan_5_.curr_instr_rd_addr__0_ ,\scan_5_.curr_instr_opcode__6_ ,
  \scan_5_.curr_instr_opcode__5_ ,\scan_5_.curr_instr_opcode__4_ ,
  \scan_5_.curr_instr_opcode__3_ ,\scan_5_.curr_instr_opcode__2_ ,\scan_5_.curr_instr_opcode__1_ ,
  \scan_5_.curr_instr_opcode__0_ ,N1645,N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,
  N1655,\scan_5_.is_br ,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,
  \scan_5_.is_jal ,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,
  \scan_5_.is_jalr ,N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,
  \scan_5_.is_link_dest ,N1687,N1688,\scan_5_.is_link_match ,\scan_5_.is_call ,
  \scan_5_.is_return ,N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,
  N1699,N1700,N1701,\scan_5_.is_cbr ,N1702,N1703,N1704,N1705,N1706,\scan_5_.is_cj ,
  N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,
  \scan_5_.is_cjr ,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,
  \scan_5_.is_cjalr ,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,
  \scan_5_.is_clink_src ,\scan_5_.is_clink_match ,\scan_5_.is_ccall ,\scan_5_.is_creturn ,
  N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,
  N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,
  N1766,N1767,N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,
  N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,
  N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,
  N1806,N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,
  N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,
  N1833,N1834,N1835,N1836,N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,
  N1846,N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,
  any_complete,N1858,N1859,N1860,N1861,any_branch,N1862,N1863,N1864,N1865,any_last_branch,
  N1866,double_branch,branch_decode_lo_br_,branch_decode_lo_jal_,
  branch_decode_lo_jalr_,branch_decode_lo_call_,branch_decode_lo__return_,branch_decode_lo_full1_,
  branch_decode_lo_full2_,branch_decode_lo_comp_,N1867,N1868,N1869,N1870,N1871,N1872,
  assembled_startup,N1873,assembled_catchup,N1874,assembled_rebase,N1875,
  assembled_linear,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,
  N1888,N1889,N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,
  N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,
  N1915,N1916,N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,
  N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,
  N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,
  N1955,N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,
  N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,
  N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,
  N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,
  N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,
  N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,
  N2035,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,
  N2048,N2049,N2050,N2051,N2052,N2053,N2054;
  wire [31:0] \scan_0_.curr_instr ,\scan_1_.curr_instr ,\scan_2_.curr_instr ,
  \scan_3_.curr_instr ,\scan_4_.curr_instr ;
  wire [5:0] branch;
  wire [4:0] complete;
  wire [46:0] next_decode_lo;
  assign fetch_scan_o[39] = 1'b0;
  assign fetch_scan_o[43] = 1'b0;
  assign fetch_scan_o[44] = 1'b0;
  assign fetch_scan_o[45] = 1'b0;
  assign fetch_scan_o[46] = 1'b0;
  assign fetch_scan_o[47] = 1'b0;
  assign fetch_scan_o[48] = 1'b0;
  assign fetch_scan_o[49] = 1'b0;
  assign fetch_scan_o[50] = 1'b0;
  assign fetch_scan_o[51] = 1'b0;
  assign fetch_scan_o[52] = 1'b0;
  assign fetch_scan_o[53] = 1'b0;
  assign fetch_scan_o[54] = 1'b0;
  assign fetch_scan_o[55] = 1'b0;
  assign fetch_scan_o[56] = 1'b0;
  assign fetch_scan_o[57] = 1'b0;
  assign fetch_scan_o[58] = 1'b0;
  assign fetch_scan_o[59] = 1'b0;
  assign fetch_scan_o[60] = 1'b0;
  assign fetch_scan_o[61] = 1'b0;
  assign fetch_scan_o[62] = 1'b0;
  assign fetch_scan_o[63] = 1'b0;
  assign fetch_scan_o[64] = 1'b0;
  assign fetch_scan_o[65] = 1'b0;
  assign fetch_scan_o[66] = 1'b0;
  assign fetch_scan_o[67] = 1'b0;
  assign fetch_scan_o[68] = 1'b0;
  assign fetch_scan_o[69] = 1'b0;
  assign fetch_scan_o[70] = 1'b0;
  assign fetch_scan_o[71] = 1'b0;
  assign fetch_scan_o[72] = 1'b0;
  assign fetch_scan_o[73] = 1'b0;
  assign fetch_scan_o[74] = 1'b0;
  assign fetch_scan_o[75] = 1'b0;
  assign fetch_scan_o[76] = 1'b0;
  assign fetch_scan_o[77] = 1'b0;
  assign fetch_scan_o[78] = 1'b0;
  assign fetch_scan_o[83] = 1'b0;
  assign fetch_scan_o[84] = 1'b0;
  assign fetch_scan_o[85] = 1'b0;
  assign fetch_scan_o[86] = 1'b0;
  assign fetch_scan_o[87] = 1'b0;
  assign fetch_scan_o[88] = 1'b0;
  assign fetch_scan_o[89] = 1'b0;
  assign fetch_scan_o[90] = 1'b0;
  assign fetch_scan_o[91] = 1'b0;
  assign fetch_scan_o[92] = 1'b0;
  assign fetch_scan_o[93] = 1'b0;
  assign fetch_scan_o[94] = 1'b0;
  assign fetch_scan_o[95] = 1'b0;
  assign fetch_scan_o[96] = 1'b0;
  assign fetch_scan_o[97] = 1'b0;
  assign fetch_scan_o[98] = 1'b0;
  assign fetch_scan_o[99] = 1'b0;
  assign fetch_scan_o[100] = 1'b0;
  assign fetch_scan_o[101] = 1'b0;
  assign fetch_scan_o[102] = 1'b0;
  assign fetch_scan_o[103] = 1'b0;
  assign fetch_scan_o[104] = 1'b0;
  assign fetch_scan_o[105] = 1'b0;
  assign fetch_scan_o[106] = 1'b0;
  assign fetch_scan_o[107] = 1'b0;
  assign fetch_scan_o[108] = 1'b0;
  assign fetch_scan_o[109] = 1'b0;
  assign fetch_scan_o[110] = 1'b0;
  assign fetch_scan_o[111] = 1'b0;
  assign fetch_scan_o[112] = 1'b0;
  assign fetch_scan_o[113] = 1'b0;
  assign fetch_scan_o[114] = 1'b0;
  assign fetch_scan_o[115] = 1'b0;
  assign fetch_scan_o[116] = 1'b0;
  assign fetch_scan_o[122] = 1'b0;
  assign fetch_scan_o[123] = 1'b0;
  assign fetch_scan_o[124] = 1'b0;
  assign assembled_yumi_o = fetch_yumi_i;
  assign fetch_v_o = assembled_v_i;
  assign fetch_pc_o[38] = assembled_pc_i[38];
  assign fetch_pc_o[37] = assembled_pc_i[37];
  assign fetch_pc_o[36] = assembled_pc_i[36];
  assign fetch_pc_o[35] = assembled_pc_i[35];
  assign fetch_pc_o[34] = assembled_pc_i[34];
  assign fetch_pc_o[33] = assembled_pc_i[33];
  assign fetch_pc_o[32] = assembled_pc_i[32];
  assign fetch_pc_o[31] = assembled_pc_i[31];
  assign fetch_pc_o[30] = assembled_pc_i[30];
  assign fetch_pc_o[29] = assembled_pc_i[29];
  assign fetch_pc_o[28] = assembled_pc_i[28];
  assign fetch_pc_o[27] = assembled_pc_i[27];
  assign fetch_pc_o[26] = assembled_pc_i[26];
  assign fetch_pc_o[25] = assembled_pc_i[25];
  assign fetch_pc_o[24] = assembled_pc_i[24];
  assign fetch_pc_o[23] = assembled_pc_i[23];
  assign fetch_pc_o[22] = assembled_pc_i[22];
  assign fetch_pc_o[21] = assembled_pc_i[21];
  assign fetch_pc_o[20] = assembled_pc_i[20];
  assign fetch_pc_o[19] = assembled_pc_i[19];
  assign fetch_pc_o[18] = assembled_pc_i[18];
  assign fetch_pc_o[17] = assembled_pc_i[17];
  assign fetch_pc_o[16] = assembled_pc_i[16];
  assign fetch_pc_o[15] = assembled_pc_i[15];
  assign fetch_pc_o[14] = assembled_pc_i[14];
  assign fetch_pc_o[13] = assembled_pc_i[13];
  assign fetch_pc_o[12] = assembled_pc_i[12];
  assign fetch_pc_o[11] = assembled_pc_i[11];
  assign fetch_pc_o[10] = assembled_pc_i[10];
  assign fetch_pc_o[9] = assembled_pc_i[9];
  assign fetch_pc_o[8] = assembled_pc_i[8];
  assign fetch_pc_o[7] = assembled_pc_i[7];
  assign fetch_pc_o[6] = assembled_pc_i[6];
  assign fetch_pc_o[5] = assembled_pc_i[5];
  assign fetch_pc_o[4] = assembled_pc_i[4];
  assign fetch_pc_o[3] = assembled_pc_i[3];
  assign fetch_pc_o[2] = assembled_pc_i[2];
  assign fetch_pc_o[1] = assembled_pc_i[1];
  assign fetch_pc_o[0] = assembled_pc_i[0];
  assign fetch_instr_o[79] = assembled_instr_i[79];
  assign fetch_instr_o[78] = assembled_instr_i[78];
  assign fetch_instr_o[77] = assembled_instr_i[77];
  assign fetch_instr_o[76] = assembled_instr_i[76];
  assign fetch_instr_o[75] = assembled_instr_i[75];
  assign fetch_instr_o[74] = assembled_instr_i[74];
  assign fetch_instr_o[73] = assembled_instr_i[73];
  assign fetch_instr_o[72] = assembled_instr_i[72];
  assign fetch_instr_o[71] = assembled_instr_i[71];
  assign fetch_instr_o[70] = assembled_instr_i[70];
  assign fetch_instr_o[69] = assembled_instr_i[69];
  assign fetch_instr_o[68] = assembled_instr_i[68];
  assign fetch_instr_o[67] = assembled_instr_i[67];
  assign fetch_instr_o[66] = assembled_instr_i[66];
  assign fetch_instr_o[65] = assembled_instr_i[65];
  assign fetch_instr_o[64] = assembled_instr_i[64];
  assign fetch_instr_o[63] = assembled_instr_i[63];
  assign fetch_instr_o[62] = assembled_instr_i[62];
  assign fetch_instr_o[61] = assembled_instr_i[61];
  assign fetch_instr_o[60] = assembled_instr_i[60];
  assign fetch_instr_o[59] = assembled_instr_i[59];
  assign fetch_instr_o[58] = assembled_instr_i[58];
  assign fetch_instr_o[57] = assembled_instr_i[57];
  assign fetch_instr_o[56] = assembled_instr_i[56];
  assign fetch_instr_o[55] = assembled_instr_i[55];
  assign fetch_instr_o[54] = assembled_instr_i[54];
  assign fetch_instr_o[53] = assembled_instr_i[53];
  assign fetch_instr_o[52] = assembled_instr_i[52];
  assign fetch_instr_o[51] = assembled_instr_i[51];
  assign fetch_instr_o[50] = assembled_instr_i[50];
  assign fetch_instr_o[49] = assembled_instr_i[49];
  assign fetch_instr_o[48] = assembled_instr_i[48];
  assign fetch_instr_o[47] = assembled_instr_i[47];
  assign fetch_instr_o[46] = assembled_instr_i[46];
  assign fetch_instr_o[45] = assembled_instr_i[45];
  assign fetch_instr_o[44] = assembled_instr_i[44];
  assign fetch_instr_o[43] = assembled_instr_i[43];
  assign fetch_instr_o[42] = assembled_instr_i[42];
  assign fetch_instr_o[41] = assembled_instr_i[41];
  assign fetch_instr_o[40] = assembled_instr_i[40];
  assign fetch_instr_o[39] = assembled_instr_i[39];
  assign fetch_instr_o[38] = assembled_instr_i[38];
  assign fetch_instr_o[37] = assembled_instr_i[37];
  assign fetch_instr_o[36] = assembled_instr_i[36];
  assign fetch_instr_o[35] = assembled_instr_i[35];
  assign fetch_instr_o[34] = assembled_instr_i[34];
  assign fetch_instr_o[33] = assembled_instr_i[33];
  assign fetch_instr_o[32] = assembled_instr_i[32];
  assign fetch_instr_o[31] = assembled_instr_i[31];
  assign fetch_instr_o[30] = assembled_instr_i[30];
  assign fetch_instr_o[29] = assembled_instr_i[29];
  assign fetch_instr_o[28] = assembled_instr_i[28];
  assign fetch_instr_o[27] = assembled_instr_i[27];
  assign fetch_instr_o[26] = assembled_instr_i[26];
  assign fetch_instr_o[25] = assembled_instr_i[25];
  assign fetch_instr_o[24] = assembled_instr_i[24];
  assign fetch_instr_o[23] = assembled_instr_i[23];
  assign fetch_instr_o[22] = assembled_instr_i[22];
  assign fetch_instr_o[21] = assembled_instr_i[21];
  assign fetch_instr_o[20] = assembled_instr_i[20];
  assign fetch_instr_o[19] = assembled_instr_i[19];
  assign fetch_instr_o[18] = assembled_instr_i[18];
  assign fetch_instr_o[17] = assembled_instr_i[17];
  assign fetch_instr_o[16] = assembled_instr_i[16];
  assign fetch_instr_o[15] = assembled_instr_i[15];
  assign fetch_instr_o[14] = assembled_instr_i[14];
  assign fetch_instr_o[13] = assembled_instr_i[13];
  assign fetch_instr_o[12] = assembled_instr_i[12];
  assign fetch_instr_o[11] = assembled_instr_i[11];
  assign fetch_instr_o[10] = assembled_instr_i[10];
  assign fetch_instr_o[9] = assembled_instr_i[9];
  assign fetch_instr_o[8] = assembled_instr_i[8];
  assign fetch_instr_o[7] = assembled_instr_i[7];
  assign fetch_instr_o[6] = assembled_instr_i[6];
  assign fetch_instr_o[5] = assembled_instr_i[5];
  assign fetch_instr_o[4] = assembled_instr_i[4];
  assign fetch_instr_o[3] = assembled_instr_i[3];
  assign fetch_instr_o[2] = assembled_instr_i[2];
  assign fetch_instr_o[1] = assembled_instr_i[1];
  assign fetch_instr_o[0] = assembled_instr_i[0];
  assign fetch_br_metadata_fwd_o[48] = assembled_br_metadata_fwd_i[48];
  assign fetch_br_metadata_fwd_o[47] = assembled_br_metadata_fwd_i[47];
  assign fetch_br_metadata_fwd_o[46] = assembled_br_metadata_fwd_i[46];
  assign fetch_br_metadata_fwd_o[45] = assembled_br_metadata_fwd_i[45];
  assign fetch_br_metadata_fwd_o[44] = assembled_br_metadata_fwd_i[44];
  assign fetch_br_metadata_fwd_o[43] = assembled_br_metadata_fwd_i[43];
  assign fetch_br_metadata_fwd_o[42] = assembled_br_metadata_fwd_i[42];
  assign fetch_br_metadata_fwd_o[41] = assembled_br_metadata_fwd_i[41];
  assign fetch_br_metadata_fwd_o[40] = assembled_br_metadata_fwd_i[40];
  assign fetch_br_metadata_fwd_o[39] = assembled_br_metadata_fwd_i[39];
  assign fetch_br_metadata_fwd_o[38] = assembled_br_metadata_fwd_i[38];
  assign fetch_br_metadata_fwd_o[37] = assembled_br_metadata_fwd_i[37];
  assign fetch_br_metadata_fwd_o[36] = assembled_br_metadata_fwd_i[36];
  assign fetch_br_metadata_fwd_o[35] = assembled_br_metadata_fwd_i[35];
  assign fetch_br_metadata_fwd_o[34] = assembled_br_metadata_fwd_i[34];
  assign fetch_br_metadata_fwd_o[33] = assembled_br_metadata_fwd_i[33];
  assign fetch_br_metadata_fwd_o[32] = assembled_br_metadata_fwd_i[32];
  assign fetch_br_metadata_fwd_o[31] = assembled_br_metadata_fwd_i[31];
  assign fetch_br_metadata_fwd_o[30] = assembled_br_metadata_fwd_i[30];
  assign fetch_br_metadata_fwd_o[29] = assembled_br_metadata_fwd_i[29];
  assign fetch_br_metadata_fwd_o[28] = assembled_br_metadata_fwd_i[28];
  assign fetch_br_metadata_fwd_o[27] = assembled_br_metadata_fwd_i[27];
  assign fetch_br_metadata_fwd_o[26] = assembled_br_metadata_fwd_i[26];
  assign fetch_br_metadata_fwd_o[25] = assembled_br_metadata_fwd_i[25];
  assign fetch_br_metadata_fwd_o[24] = assembled_br_metadata_fwd_i[24];
  assign fetch_br_metadata_fwd_o[23] = assembled_br_metadata_fwd_i[23];
  assign fetch_br_metadata_fwd_o[22] = assembled_br_metadata_fwd_i[22];
  assign fetch_br_metadata_fwd_o[21] = assembled_br_metadata_fwd_i[21];
  assign fetch_br_metadata_fwd_o[20] = assembled_br_metadata_fwd_i[20];
  assign fetch_br_metadata_fwd_o[19] = assembled_br_metadata_fwd_i[19];
  assign fetch_br_metadata_fwd_o[18] = assembled_br_metadata_fwd_i[18];
  assign fetch_br_metadata_fwd_o[17] = assembled_br_metadata_fwd_i[17];
  assign fetch_br_metadata_fwd_o[16] = assembled_br_metadata_fwd_i[16];
  assign fetch_br_metadata_fwd_o[15] = assembled_br_metadata_fwd_i[15];
  assign fetch_br_metadata_fwd_o[14] = assembled_br_metadata_fwd_i[14];
  assign fetch_br_metadata_fwd_o[13] = assembled_br_metadata_fwd_i[13];
  assign fetch_br_metadata_fwd_o[12] = assembled_br_metadata_fwd_i[12];
  assign fetch_br_metadata_fwd_o[11] = assembled_br_metadata_fwd_i[11];
  assign fetch_br_metadata_fwd_o[10] = assembled_br_metadata_fwd_i[10];
  assign fetch_br_metadata_fwd_o[9] = assembled_br_metadata_fwd_i[9];
  assign fetch_br_metadata_fwd_o[8] = assembled_br_metadata_fwd_i[8];
  assign fetch_br_metadata_fwd_o[7] = assembled_br_metadata_fwd_i[7];
  assign fetch_br_metadata_fwd_o[6] = assembled_br_metadata_fwd_i[6];
  assign fetch_br_metadata_fwd_o[5] = assembled_br_metadata_fwd_i[5];
  assign fetch_br_metadata_fwd_o[4] = assembled_br_metadata_fwd_i[4];
  assign fetch_br_metadata_fwd_o[3] = assembled_br_metadata_fwd_i[3];
  assign fetch_br_metadata_fwd_o[2] = assembled_br_metadata_fwd_i[2];
  assign fetch_br_metadata_fwd_o[1] = assembled_br_metadata_fwd_i[1];
  assign fetch_br_metadata_fwd_o[0] = assembled_br_metadata_fwd_i[0];
  assign fetch_partial_o = assembled_partial_i;
  assign N25 = 1'b0 < assembled_count_i;
  assign N28 = ~\scan_0_.curr_instr [6];
  assign N29 = ~\scan_0_.curr_instr [5];
  assign N30 = ~\scan_0_.curr_instr [1];
  assign N31 = ~\scan_0_.curr_instr [0];
  assign N32 = N29 | N28;
  assign N33 = \scan_0_.curr_instr [4] | N32;
  assign N34 = \scan_0_.curr_instr [3] | N33;
  assign N35 = \scan_0_.curr_instr [2] | N34;
  assign N36 = N30 | N35;
  assign N37 = N31 | N36;
  assign N38 = ~N37;
  assign N39 = ~\scan_0_.curr_instr [3];
  assign N40 = ~\scan_0_.curr_instr [2];
  assign N41 = N29 | N28;
  assign N42 = \scan_0_.curr_instr [4] | N41;
  assign N43 = N39 | N42;
  assign N44 = N40 | N43;
  assign N45 = N30 | N44;
  assign N46 = N31 | N45;
  assign N47 = ~N46;
  assign N48 = \scan_0_.curr_instr [13] | \scan_0_.curr_instr [14];
  assign N49 = \scan_0_.curr_instr [12] | N48;
  assign N50 = N28 | N49;
  assign N51 = N29 | N50;
  assign N52 = \scan_0_.curr_instr [4] | N51;
  assign N53 = \scan_0_.curr_instr [3] | N52;
  assign N54 = N40 | N53;
  assign N55 = N30 | N54;
  assign N56 = N31 | N55;
  assign N57 = ~N56;
  assign N58 = ~\scan_0_.curr_instr [7];
  assign N59 = \scan_0_.curr_instr [10] | \scan_0_.curr_instr [11];
  assign N60 = \scan_0_.curr_instr [9] | N59;
  assign N61 = \scan_0_.curr_instr [8] | N60;
  assign N62 = N58 | N61;
  assign N63 = ~N62;
  assign N64 = ~\scan_0_.curr_instr [9];
  assign N65 = \scan_0_.curr_instr [10] | \scan_0_.curr_instr [11];
  assign N66 = N64 | N65;
  assign N67 = \scan_0_.curr_instr [8] | N66;
  assign N68 = N58 | N67;
  assign N69 = ~N68;
  assign \scan_0_.is_link_dest  = N63 | N69;
  assign N70 = ~\scan_0_.curr_instr [15];
  assign N71 = \scan_0_.curr_instr [18] | \scan_0_.curr_instr [19];
  assign N72 = \scan_0_.curr_instr [17] | N71;
  assign N73 = \scan_0_.curr_instr [16] | N72;
  assign N74 = N70 | N73;
  assign N75 = ~N74;
  assign N76 = ~\scan_0_.curr_instr [17];
  assign N77 = \scan_0_.curr_instr [18] | \scan_0_.curr_instr [19];
  assign N78 = N76 | N77;
  assign N79 = \scan_0_.curr_instr [16] | N78;
  assign N80 = N70 | N79;
  assign N81 = ~N80;
  assign \scan_0_.is_link_src  = N75 | N81;
  assign N82 = \scan_0_.curr_instr [11:7] == \scan_0_.curr_instr [19:15];
  assign N83 = ~\scan_0_.curr_instr [14];
  assign N84 = \scan_0_.curr_instr [30] | \scan_0_.curr_instr [31];
  assign N85 = \scan_0_.curr_instr [29] | N84;
  assign N86 = \scan_0_.curr_instr [28] | N85;
  assign N87 = \scan_0_.curr_instr [27] | N86;
  assign N88 = \scan_0_.curr_instr [26] | N87;
  assign N89 = \scan_0_.curr_instr [25] | N88;
  assign N90 = \scan_0_.curr_instr [24] | N89;
  assign N91 = \scan_0_.curr_instr [23] | N90;
  assign N92 = \scan_0_.curr_instr [22] | N91;
  assign N93 = \scan_0_.curr_instr [21] | N92;
  assign N94 = \scan_0_.curr_instr [20] | N93;
  assign N95 = \scan_0_.curr_instr [19] | N94;
  assign N96 = \scan_0_.curr_instr [18] | N95;
  assign N97 = \scan_0_.curr_instr [17] | N96;
  assign N98 = \scan_0_.curr_instr [16] | N97;
  assign N99 = N70 | N98;
  assign N100 = N83 | N99;
  assign N101 = \scan_0_.curr_instr [13] | N100;
  assign N102 = \scan_0_.curr_instr [1] | N101;
  assign N103 = N31 | N102;
  assign N104 = ~N103;
  assign N105 = ~\scan_0_.curr_instr [13];
  assign N106 = \scan_0_.curr_instr [30] | \scan_0_.curr_instr [31];
  assign N107 = \scan_0_.curr_instr [29] | N106;
  assign N108 = \scan_0_.curr_instr [28] | N107;
  assign N109 = \scan_0_.curr_instr [27] | N108;
  assign N110 = \scan_0_.curr_instr [26] | N109;
  assign N111 = \scan_0_.curr_instr [25] | N110;
  assign N112 = \scan_0_.curr_instr [24] | N111;
  assign N113 = \scan_0_.curr_instr [23] | N112;
  assign N114 = \scan_0_.curr_instr [22] | N113;
  assign N115 = \scan_0_.curr_instr [21] | N114;
  assign N116 = \scan_0_.curr_instr [20] | N115;
  assign N117 = \scan_0_.curr_instr [19] | N116;
  assign N118 = \scan_0_.curr_instr [18] | N117;
  assign N119 = \scan_0_.curr_instr [17] | N118;
  assign N120 = \scan_0_.curr_instr [16] | N119;
  assign N121 = N70 | N120;
  assign N122 = N83 | N121;
  assign N123 = N105 | N122;
  assign N124 = \scan_0_.curr_instr [1] | N123;
  assign N125 = N31 | N124;
  assign N126 = ~N125;
  assign N127 = N104 | N126;
  assign N128 = \scan_0_.curr_instr [30] | \scan_0_.curr_instr [31];
  assign N129 = \scan_0_.curr_instr [29] | N128;
  assign N130 = \scan_0_.curr_instr [28] | N129;
  assign N131 = \scan_0_.curr_instr [27] | N130;
  assign N132 = \scan_0_.curr_instr [26] | N131;
  assign N133 = \scan_0_.curr_instr [25] | N132;
  assign N134 = \scan_0_.curr_instr [24] | N133;
  assign N135 = \scan_0_.curr_instr [23] | N134;
  assign N136 = \scan_0_.curr_instr [22] | N135;
  assign N137 = \scan_0_.curr_instr [21] | N136;
  assign N138 = \scan_0_.curr_instr [20] | N137;
  assign N139 = \scan_0_.curr_instr [19] | N138;
  assign N140 = \scan_0_.curr_instr [18] | N139;
  assign N141 = \scan_0_.curr_instr [17] | N140;
  assign N142 = \scan_0_.curr_instr [16] | N141;
  assign N143 = N70 | N142;
  assign N144 = \scan_0_.curr_instr [14] | N143;
  assign N145 = N105 | N144;
  assign N146 = \scan_0_.curr_instr [1] | N145;
  assign N147 = N31 | N146;
  assign N148 = ~N147;
  assign N149 = \scan_0_.curr_instr [30] | \scan_0_.curr_instr [31];
  assign N150 = \scan_0_.curr_instr [29] | N149;
  assign N151 = \scan_0_.curr_instr [28] | N150;
  assign N152 = \scan_0_.curr_instr [27] | N151;
  assign N153 = \scan_0_.curr_instr [26] | N152;
  assign N154 = \scan_0_.curr_instr [25] | N153;
  assign N155 = \scan_0_.curr_instr [24] | N154;
  assign N156 = \scan_0_.curr_instr [23] | N155;
  assign N157 = \scan_0_.curr_instr [22] | N156;
  assign N158 = \scan_0_.curr_instr [21] | N157;
  assign N159 = \scan_0_.curr_instr [20] | N158;
  assign N160 = \scan_0_.curr_instr [19] | N159;
  assign N161 = \scan_0_.curr_instr [18] | N160;
  assign N162 = \scan_0_.curr_instr [17] | N161;
  assign N163 = \scan_0_.curr_instr [16] | N162;
  assign N164 = N70 | N163;
  assign N165 = \scan_0_.curr_instr [14] | N164;
  assign N166 = \scan_0_.curr_instr [13] | N165;
  assign N167 = \scan_0_.curr_instr [12] | N166;
  assign N168 = \scan_0_.curr_instr [6] | N167;
  assign N169 = \scan_0_.curr_instr [5] | N168;
  assign N170 = \scan_0_.curr_instr [4] | N169;
  assign N171 = \scan_0_.curr_instr [3] | N170;
  assign N172 = \scan_0_.curr_instr [2] | N171;
  assign N173 = N30 | N172;
  assign N174 = \scan_0_.curr_instr [0] | N173;
  assign N175 = ~N174;
  assign N176 = ~\scan_0_.curr_instr [12];
  assign N177 = \scan_0_.curr_instr [30] | \scan_0_.curr_instr [31];
  assign N178 = \scan_0_.curr_instr [29] | N177;
  assign N179 = \scan_0_.curr_instr [28] | N178;
  assign N180 = \scan_0_.curr_instr [27] | N179;
  assign N181 = \scan_0_.curr_instr [26] | N180;
  assign N182 = \scan_0_.curr_instr [25] | N181;
  assign N183 = \scan_0_.curr_instr [24] | N182;
  assign N184 = \scan_0_.curr_instr [23] | N183;
  assign N185 = \scan_0_.curr_instr [22] | N184;
  assign N186 = \scan_0_.curr_instr [21] | N185;
  assign N187 = \scan_0_.curr_instr [20] | N186;
  assign N188 = \scan_0_.curr_instr [19] | N187;
  assign N189 = \scan_0_.curr_instr [18] | N188;
  assign N190 = \scan_0_.curr_instr [17] | N189;
  assign N191 = \scan_0_.curr_instr [16] | N190;
  assign N192 = N70 | N191;
  assign N193 = \scan_0_.curr_instr [14] | N192;
  assign N194 = \scan_0_.curr_instr [13] | N193;
  assign N195 = N176 | N194;
  assign N196 = \scan_0_.curr_instr [6] | N195;
  assign N197 = \scan_0_.curr_instr [5] | N196;
  assign N198 = \scan_0_.curr_instr [4] | N197;
  assign N199 = \scan_0_.curr_instr [3] | N198;
  assign N200 = \scan_0_.curr_instr [2] | N199;
  assign N201 = N30 | N200;
  assign N202 = \scan_0_.curr_instr [0] | N201;
  assign N203 = ~N202;
  assign N204 = \scan_0_.curr_instr [10] | \scan_0_.curr_instr [11];
  assign N205 = \scan_0_.curr_instr [9] | N204;
  assign N206 = \scan_0_.curr_instr [8] | N205;
  assign N207 = N58 | N206;
  assign N208 = ~N207;
  assign N209 = \scan_0_.curr_instr [10] | \scan_0_.curr_instr [11];
  assign N210 = N64 | N209;
  assign N211 = \scan_0_.curr_instr [8] | N210;
  assign N212 = N58 | N211;
  assign N213 = ~N212;
  assign \scan_0_.is_clink_src  = N208 | N213;
  assign N301 = 1'b1 < assembled_count_i;
  assign N304 = ~\scan_1_.curr_instr [6];
  assign N305 = ~\scan_1_.curr_instr [5];
  assign N306 = ~\scan_1_.curr_instr [1];
  assign N307 = ~\scan_1_.curr_instr [0];
  assign N308 = N305 | N304;
  assign N309 = \scan_1_.curr_instr [4] | N308;
  assign N310 = \scan_1_.curr_instr [3] | N309;
  assign N311 = \scan_1_.curr_instr [2] | N310;
  assign N312 = N306 | N311;
  assign N313 = N307 | N312;
  assign N314 = ~N313;
  assign N315 = ~\scan_1_.curr_instr [3];
  assign N316 = ~\scan_1_.curr_instr [2];
  assign N317 = N305 | N304;
  assign N318 = \scan_1_.curr_instr [4] | N317;
  assign N319 = N315 | N318;
  assign N320 = N316 | N319;
  assign N321 = N306 | N320;
  assign N322 = N307 | N321;
  assign N323 = ~N322;
  assign N324 = \scan_1_.curr_instr [13] | \scan_1_.curr_instr [14];
  assign N325 = \scan_1_.curr_instr [12] | N324;
  assign N326 = N304 | N325;
  assign N327 = N305 | N326;
  assign N328 = \scan_1_.curr_instr [4] | N327;
  assign N329 = \scan_1_.curr_instr [3] | N328;
  assign N330 = N316 | N329;
  assign N331 = N306 | N330;
  assign N332 = N307 | N331;
  assign N333 = ~N332;
  assign N334 = ~\scan_1_.curr_instr [7];
  assign N335 = \scan_1_.curr_instr [10] | \scan_1_.curr_instr [11];
  assign N336 = \scan_1_.curr_instr [9] | N335;
  assign N337 = \scan_1_.curr_instr [8] | N336;
  assign N338 = N334 | N337;
  assign N339 = ~N338;
  assign N340 = ~\scan_1_.curr_instr [9];
  assign N341 = \scan_1_.curr_instr [10] | \scan_1_.curr_instr [11];
  assign N342 = N340 | N341;
  assign N343 = \scan_1_.curr_instr [8] | N342;
  assign N344 = N334 | N343;
  assign N345 = ~N344;
  assign \scan_1_.is_link_dest  = N339 | N345;
  assign N346 = ~\scan_1_.curr_instr [15];
  assign N347 = \scan_1_.curr_instr [18] | \scan_1_.curr_instr [19];
  assign N348 = \scan_1_.curr_instr [17] | N347;
  assign N349 = \scan_1_.curr_instr [16] | N348;
  assign N350 = N346 | N349;
  assign N351 = ~N350;
  assign N352 = ~\scan_1_.curr_instr [17];
  assign N353 = \scan_1_.curr_instr [18] | \scan_1_.curr_instr [19];
  assign N354 = N352 | N353;
  assign N355 = \scan_1_.curr_instr [16] | N354;
  assign N356 = N346 | N355;
  assign N357 = ~N356;
  assign \scan_1_.is_link_src  = N351 | N357;
  assign N358 = \scan_1_.curr_instr [11:7] == \scan_1_.curr_instr [19:15];
  assign N359 = ~\scan_1_.curr_instr [14];
  assign N360 = \scan_1_.curr_instr [30] | \scan_1_.curr_instr [31];
  assign N361 = \scan_1_.curr_instr [29] | N360;
  assign N362 = \scan_1_.curr_instr [28] | N361;
  assign N363 = \scan_1_.curr_instr [27] | N362;
  assign N364 = \scan_1_.curr_instr [26] | N363;
  assign N365 = \scan_1_.curr_instr [25] | N364;
  assign N366 = \scan_1_.curr_instr [24] | N365;
  assign N367 = \scan_1_.curr_instr [23] | N366;
  assign N368 = \scan_1_.curr_instr [22] | N367;
  assign N369 = \scan_1_.curr_instr [21] | N368;
  assign N370 = \scan_1_.curr_instr [20] | N369;
  assign N371 = \scan_1_.curr_instr [19] | N370;
  assign N372 = \scan_1_.curr_instr [18] | N371;
  assign N373 = \scan_1_.curr_instr [17] | N372;
  assign N374 = \scan_1_.curr_instr [16] | N373;
  assign N375 = N346 | N374;
  assign N376 = N359 | N375;
  assign N377 = \scan_1_.curr_instr [13] | N376;
  assign N378 = \scan_1_.curr_instr [1] | N377;
  assign N379 = N307 | N378;
  assign N380 = ~N379;
  assign N381 = ~\scan_1_.curr_instr [13];
  assign N382 = \scan_1_.curr_instr [30] | \scan_1_.curr_instr [31];
  assign N383 = \scan_1_.curr_instr [29] | N382;
  assign N384 = \scan_1_.curr_instr [28] | N383;
  assign N385 = \scan_1_.curr_instr [27] | N384;
  assign N386 = \scan_1_.curr_instr [26] | N385;
  assign N387 = \scan_1_.curr_instr [25] | N386;
  assign N388 = \scan_1_.curr_instr [24] | N387;
  assign N389 = \scan_1_.curr_instr [23] | N388;
  assign N390 = \scan_1_.curr_instr [22] | N389;
  assign N391 = \scan_1_.curr_instr [21] | N390;
  assign N392 = \scan_1_.curr_instr [20] | N391;
  assign N393 = \scan_1_.curr_instr [19] | N392;
  assign N394 = \scan_1_.curr_instr [18] | N393;
  assign N395 = \scan_1_.curr_instr [17] | N394;
  assign N396 = \scan_1_.curr_instr [16] | N395;
  assign N397 = N346 | N396;
  assign N398 = N359 | N397;
  assign N399 = N381 | N398;
  assign N400 = \scan_1_.curr_instr [1] | N399;
  assign N401 = N307 | N400;
  assign N402 = ~N401;
  assign N403 = N380 | N402;
  assign N404 = \scan_1_.curr_instr [30] | \scan_1_.curr_instr [31];
  assign N405 = \scan_1_.curr_instr [29] | N404;
  assign N406 = \scan_1_.curr_instr [28] | N405;
  assign N407 = \scan_1_.curr_instr [27] | N406;
  assign N408 = \scan_1_.curr_instr [26] | N407;
  assign N409 = \scan_1_.curr_instr [25] | N408;
  assign N410 = \scan_1_.curr_instr [24] | N409;
  assign N411 = \scan_1_.curr_instr [23] | N410;
  assign N412 = \scan_1_.curr_instr [22] | N411;
  assign N413 = \scan_1_.curr_instr [21] | N412;
  assign N414 = \scan_1_.curr_instr [20] | N413;
  assign N415 = \scan_1_.curr_instr [19] | N414;
  assign N416 = \scan_1_.curr_instr [18] | N415;
  assign N417 = \scan_1_.curr_instr [17] | N416;
  assign N418 = \scan_1_.curr_instr [16] | N417;
  assign N419 = N346 | N418;
  assign N420 = \scan_1_.curr_instr [14] | N419;
  assign N421 = N381 | N420;
  assign N422 = \scan_1_.curr_instr [1] | N421;
  assign N423 = N307 | N422;
  assign N424 = ~N423;
  assign N425 = \scan_1_.curr_instr [30] | \scan_1_.curr_instr [31];
  assign N426 = \scan_1_.curr_instr [29] | N425;
  assign N427 = \scan_1_.curr_instr [28] | N426;
  assign N428 = \scan_1_.curr_instr [27] | N427;
  assign N429 = \scan_1_.curr_instr [26] | N428;
  assign N430 = \scan_1_.curr_instr [25] | N429;
  assign N431 = \scan_1_.curr_instr [24] | N430;
  assign N432 = \scan_1_.curr_instr [23] | N431;
  assign N433 = \scan_1_.curr_instr [22] | N432;
  assign N434 = \scan_1_.curr_instr [21] | N433;
  assign N435 = \scan_1_.curr_instr [20] | N434;
  assign N436 = \scan_1_.curr_instr [19] | N435;
  assign N437 = \scan_1_.curr_instr [18] | N436;
  assign N438 = \scan_1_.curr_instr [17] | N437;
  assign N439 = \scan_1_.curr_instr [16] | N438;
  assign N440 = N346 | N439;
  assign N441 = \scan_1_.curr_instr [14] | N440;
  assign N442 = \scan_1_.curr_instr [13] | N441;
  assign N443 = \scan_1_.curr_instr [12] | N442;
  assign N444 = \scan_1_.curr_instr [6] | N443;
  assign N445 = \scan_1_.curr_instr [5] | N444;
  assign N446 = \scan_1_.curr_instr [4] | N445;
  assign N447 = \scan_1_.curr_instr [3] | N446;
  assign N448 = \scan_1_.curr_instr [2] | N447;
  assign N449 = N306 | N448;
  assign N450 = \scan_1_.curr_instr [0] | N449;
  assign N451 = ~N450;
  assign N452 = ~\scan_1_.curr_instr [12];
  assign N453 = \scan_1_.curr_instr [30] | \scan_1_.curr_instr [31];
  assign N454 = \scan_1_.curr_instr [29] | N453;
  assign N455 = \scan_1_.curr_instr [28] | N454;
  assign N456 = \scan_1_.curr_instr [27] | N455;
  assign N457 = \scan_1_.curr_instr [26] | N456;
  assign N458 = \scan_1_.curr_instr [25] | N457;
  assign N459 = \scan_1_.curr_instr [24] | N458;
  assign N460 = \scan_1_.curr_instr [23] | N459;
  assign N461 = \scan_1_.curr_instr [22] | N460;
  assign N462 = \scan_1_.curr_instr [21] | N461;
  assign N463 = \scan_1_.curr_instr [20] | N462;
  assign N464 = \scan_1_.curr_instr [19] | N463;
  assign N465 = \scan_1_.curr_instr [18] | N464;
  assign N466 = \scan_1_.curr_instr [17] | N465;
  assign N467 = \scan_1_.curr_instr [16] | N466;
  assign N468 = N346 | N467;
  assign N469 = \scan_1_.curr_instr [14] | N468;
  assign N470 = \scan_1_.curr_instr [13] | N469;
  assign N471 = N452 | N470;
  assign N472 = \scan_1_.curr_instr [6] | N471;
  assign N473 = \scan_1_.curr_instr [5] | N472;
  assign N474 = \scan_1_.curr_instr [4] | N473;
  assign N475 = \scan_1_.curr_instr [3] | N474;
  assign N476 = \scan_1_.curr_instr [2] | N475;
  assign N477 = N306 | N476;
  assign N478 = \scan_1_.curr_instr [0] | N477;
  assign N479 = ~N478;
  assign N480 = \scan_1_.curr_instr [10] | \scan_1_.curr_instr [11];
  assign N481 = \scan_1_.curr_instr [9] | N480;
  assign N482 = \scan_1_.curr_instr [8] | N481;
  assign N483 = N334 | N482;
  assign N484 = ~N483;
  assign N485 = \scan_1_.curr_instr [10] | \scan_1_.curr_instr [11];
  assign N486 = N340 | N485;
  assign N487 = \scan_1_.curr_instr [8] | N486;
  assign N488 = N334 | N487;
  assign N489 = ~N488;
  assign \scan_1_.is_clink_src  = N484 | N489;
  assign N577 = { 1'b1, 1'b0 } < assembled_count_i;
  assign N580 = ~\scan_2_.curr_instr [6];
  assign N581 = ~\scan_2_.curr_instr [5];
  assign N582 = ~\scan_2_.curr_instr [1];
  assign N583 = ~\scan_2_.curr_instr [0];
  assign N584 = N581 | N580;
  assign N585 = \scan_2_.curr_instr [4] | N584;
  assign N586 = \scan_2_.curr_instr [3] | N585;
  assign N587 = \scan_2_.curr_instr [2] | N586;
  assign N588 = N582 | N587;
  assign N589 = N583 | N588;
  assign N590 = ~N589;
  assign N591 = ~\scan_2_.curr_instr [3];
  assign N592 = ~\scan_2_.curr_instr [2];
  assign N593 = N581 | N580;
  assign N594 = \scan_2_.curr_instr [4] | N593;
  assign N595 = N591 | N594;
  assign N596 = N592 | N595;
  assign N597 = N582 | N596;
  assign N598 = N583 | N597;
  assign N599 = ~N598;
  assign N600 = \scan_2_.curr_instr [13] | \scan_2_.curr_instr [14];
  assign N601 = \scan_2_.curr_instr [12] | N600;
  assign N602 = N580 | N601;
  assign N603 = N581 | N602;
  assign N604 = \scan_2_.curr_instr [4] | N603;
  assign N605 = \scan_2_.curr_instr [3] | N604;
  assign N606 = N592 | N605;
  assign N607 = N582 | N606;
  assign N608 = N583 | N607;
  assign N609 = ~N608;
  assign N610 = ~\scan_2_.curr_instr [7];
  assign N611 = \scan_2_.curr_instr [10] | \scan_2_.curr_instr [11];
  assign N612 = \scan_2_.curr_instr [9] | N611;
  assign N613 = \scan_2_.curr_instr [8] | N612;
  assign N614 = N610 | N613;
  assign N615 = ~N614;
  assign N616 = ~\scan_2_.curr_instr [9];
  assign N617 = \scan_2_.curr_instr [10] | \scan_2_.curr_instr [11];
  assign N618 = N616 | N617;
  assign N619 = \scan_2_.curr_instr [8] | N618;
  assign N620 = N610 | N619;
  assign N621 = ~N620;
  assign \scan_2_.is_link_dest  = N615 | N621;
  assign N622 = ~\scan_2_.curr_instr [15];
  assign N623 = \scan_2_.curr_instr [18] | \scan_2_.curr_instr [19];
  assign N624 = \scan_2_.curr_instr [17] | N623;
  assign N625 = \scan_2_.curr_instr [16] | N624;
  assign N626 = N622 | N625;
  assign N627 = ~N626;
  assign N628 = ~\scan_2_.curr_instr [17];
  assign N629 = \scan_2_.curr_instr [18] | \scan_2_.curr_instr [19];
  assign N630 = N628 | N629;
  assign N631 = \scan_2_.curr_instr [16] | N630;
  assign N632 = N622 | N631;
  assign N633 = ~N632;
  assign \scan_2_.is_link_src  = N627 | N633;
  assign N634 = \scan_2_.curr_instr [11:7] == \scan_2_.curr_instr [19:15];
  assign N635 = ~\scan_2_.curr_instr [14];
  assign N636 = \scan_2_.curr_instr [30] | \scan_2_.curr_instr [31];
  assign N637 = \scan_2_.curr_instr [29] | N636;
  assign N638 = \scan_2_.curr_instr [28] | N637;
  assign N639 = \scan_2_.curr_instr [27] | N638;
  assign N640 = \scan_2_.curr_instr [26] | N639;
  assign N641 = \scan_2_.curr_instr [25] | N640;
  assign N642 = \scan_2_.curr_instr [24] | N641;
  assign N643 = \scan_2_.curr_instr [23] | N642;
  assign N644 = \scan_2_.curr_instr [22] | N643;
  assign N645 = \scan_2_.curr_instr [21] | N644;
  assign N646 = \scan_2_.curr_instr [20] | N645;
  assign N647 = \scan_2_.curr_instr [19] | N646;
  assign N648 = \scan_2_.curr_instr [18] | N647;
  assign N649 = \scan_2_.curr_instr [17] | N648;
  assign N650 = \scan_2_.curr_instr [16] | N649;
  assign N651 = N622 | N650;
  assign N652 = N635 | N651;
  assign N653 = \scan_2_.curr_instr [13] | N652;
  assign N654 = \scan_2_.curr_instr [1] | N653;
  assign N655 = N583 | N654;
  assign N656 = ~N655;
  assign N657 = ~\scan_2_.curr_instr [13];
  assign N658 = \scan_2_.curr_instr [30] | \scan_2_.curr_instr [31];
  assign N659 = \scan_2_.curr_instr [29] | N658;
  assign N660 = \scan_2_.curr_instr [28] | N659;
  assign N661 = \scan_2_.curr_instr [27] | N660;
  assign N662 = \scan_2_.curr_instr [26] | N661;
  assign N663 = \scan_2_.curr_instr [25] | N662;
  assign N664 = \scan_2_.curr_instr [24] | N663;
  assign N665 = \scan_2_.curr_instr [23] | N664;
  assign N666 = \scan_2_.curr_instr [22] | N665;
  assign N667 = \scan_2_.curr_instr [21] | N666;
  assign N668 = \scan_2_.curr_instr [20] | N667;
  assign N669 = \scan_2_.curr_instr [19] | N668;
  assign N670 = \scan_2_.curr_instr [18] | N669;
  assign N671 = \scan_2_.curr_instr [17] | N670;
  assign N672 = \scan_2_.curr_instr [16] | N671;
  assign N673 = N622 | N672;
  assign N674 = N635 | N673;
  assign N675 = N657 | N674;
  assign N676 = \scan_2_.curr_instr [1] | N675;
  assign N677 = N583 | N676;
  assign N678 = ~N677;
  assign N679 = N656 | N678;
  assign N680 = \scan_2_.curr_instr [30] | \scan_2_.curr_instr [31];
  assign N681 = \scan_2_.curr_instr [29] | N680;
  assign N682 = \scan_2_.curr_instr [28] | N681;
  assign N683 = \scan_2_.curr_instr [27] | N682;
  assign N684 = \scan_2_.curr_instr [26] | N683;
  assign N685 = \scan_2_.curr_instr [25] | N684;
  assign N686 = \scan_2_.curr_instr [24] | N685;
  assign N687 = \scan_2_.curr_instr [23] | N686;
  assign N688 = \scan_2_.curr_instr [22] | N687;
  assign N689 = \scan_2_.curr_instr [21] | N688;
  assign N690 = \scan_2_.curr_instr [20] | N689;
  assign N691 = \scan_2_.curr_instr [19] | N690;
  assign N692 = \scan_2_.curr_instr [18] | N691;
  assign N693 = \scan_2_.curr_instr [17] | N692;
  assign N694 = \scan_2_.curr_instr [16] | N693;
  assign N695 = N622 | N694;
  assign N696 = \scan_2_.curr_instr [14] | N695;
  assign N697 = N657 | N696;
  assign N698 = \scan_2_.curr_instr [1] | N697;
  assign N699 = N583 | N698;
  assign N700 = ~N699;
  assign N701 = \scan_2_.curr_instr [30] | \scan_2_.curr_instr [31];
  assign N702 = \scan_2_.curr_instr [29] | N701;
  assign N703 = \scan_2_.curr_instr [28] | N702;
  assign N704 = \scan_2_.curr_instr [27] | N703;
  assign N705 = \scan_2_.curr_instr [26] | N704;
  assign N706 = \scan_2_.curr_instr [25] | N705;
  assign N707 = \scan_2_.curr_instr [24] | N706;
  assign N708 = \scan_2_.curr_instr [23] | N707;
  assign N709 = \scan_2_.curr_instr [22] | N708;
  assign N710 = \scan_2_.curr_instr [21] | N709;
  assign N711 = \scan_2_.curr_instr [20] | N710;
  assign N712 = \scan_2_.curr_instr [19] | N711;
  assign N713 = \scan_2_.curr_instr [18] | N712;
  assign N714 = \scan_2_.curr_instr [17] | N713;
  assign N715 = \scan_2_.curr_instr [16] | N714;
  assign N716 = N622 | N715;
  assign N717 = \scan_2_.curr_instr [14] | N716;
  assign N718 = \scan_2_.curr_instr [13] | N717;
  assign N719 = \scan_2_.curr_instr [12] | N718;
  assign N720 = \scan_2_.curr_instr [6] | N719;
  assign N721 = \scan_2_.curr_instr [5] | N720;
  assign N722 = \scan_2_.curr_instr [4] | N721;
  assign N723 = \scan_2_.curr_instr [3] | N722;
  assign N724 = \scan_2_.curr_instr [2] | N723;
  assign N725 = N582 | N724;
  assign N726 = \scan_2_.curr_instr [0] | N725;
  assign N727 = ~N726;
  assign N728 = ~\scan_2_.curr_instr [12];
  assign N729 = \scan_2_.curr_instr [30] | \scan_2_.curr_instr [31];
  assign N730 = \scan_2_.curr_instr [29] | N729;
  assign N731 = \scan_2_.curr_instr [28] | N730;
  assign N732 = \scan_2_.curr_instr [27] | N731;
  assign N733 = \scan_2_.curr_instr [26] | N732;
  assign N734 = \scan_2_.curr_instr [25] | N733;
  assign N735 = \scan_2_.curr_instr [24] | N734;
  assign N736 = \scan_2_.curr_instr [23] | N735;
  assign N737 = \scan_2_.curr_instr [22] | N736;
  assign N738 = \scan_2_.curr_instr [21] | N737;
  assign N739 = \scan_2_.curr_instr [20] | N738;
  assign N740 = \scan_2_.curr_instr [19] | N739;
  assign N741 = \scan_2_.curr_instr [18] | N740;
  assign N742 = \scan_2_.curr_instr [17] | N741;
  assign N743 = \scan_2_.curr_instr [16] | N742;
  assign N744 = N622 | N743;
  assign N745 = \scan_2_.curr_instr [14] | N744;
  assign N746 = \scan_2_.curr_instr [13] | N745;
  assign N747 = N728 | N746;
  assign N748 = \scan_2_.curr_instr [6] | N747;
  assign N749 = \scan_2_.curr_instr [5] | N748;
  assign N750 = \scan_2_.curr_instr [4] | N749;
  assign N751 = \scan_2_.curr_instr [3] | N750;
  assign N752 = \scan_2_.curr_instr [2] | N751;
  assign N753 = N582 | N752;
  assign N754 = \scan_2_.curr_instr [0] | N753;
  assign N755 = ~N754;
  assign N756 = \scan_2_.curr_instr [10] | \scan_2_.curr_instr [11];
  assign N757 = \scan_2_.curr_instr [9] | N756;
  assign N758 = \scan_2_.curr_instr [8] | N757;
  assign N759 = N610 | N758;
  assign N760 = ~N759;
  assign N761 = \scan_2_.curr_instr [10] | \scan_2_.curr_instr [11];
  assign N762 = N616 | N761;
  assign N763 = \scan_2_.curr_instr [8] | N762;
  assign N764 = N610 | N763;
  assign N765 = ~N764;
  assign \scan_2_.is_clink_src  = N760 | N765;
  assign N932 = { 1'b1, 1'b1 } < assembled_count_i;
  assign N935 = ~\scan_3_.curr_instr [6];
  assign N936 = ~\scan_3_.curr_instr [5];
  assign N937 = ~\scan_3_.curr_instr [1];
  assign N938 = ~\scan_3_.curr_instr [0];
  assign N939 = N936 | N935;
  assign N940 = \scan_3_.curr_instr [4] | N939;
  assign N941 = \scan_3_.curr_instr [3] | N940;
  assign N942 = \scan_3_.curr_instr [2] | N941;
  assign N943 = N937 | N942;
  assign N944 = N938 | N943;
  assign N945 = ~N944;
  assign N946 = ~\scan_3_.curr_instr [3];
  assign N947 = ~\scan_3_.curr_instr [2];
  assign N948 = N936 | N935;
  assign N949 = \scan_3_.curr_instr [4] | N948;
  assign N950 = N946 | N949;
  assign N951 = N947 | N950;
  assign N952 = N937 | N951;
  assign N953 = N938 | N952;
  assign N954 = ~N953;
  assign N955 = \scan_3_.curr_instr [13] | \scan_3_.curr_instr [14];
  assign N956 = \scan_3_.curr_instr [12] | N955;
  assign N957 = N935 | N956;
  assign N958 = N936 | N957;
  assign N959 = \scan_3_.curr_instr [4] | N958;
  assign N960 = \scan_3_.curr_instr [3] | N959;
  assign N961 = N947 | N960;
  assign N962 = N937 | N961;
  assign N963 = N938 | N962;
  assign N964 = ~N963;
  assign N965 = ~\scan_3_.curr_instr [7];
  assign N966 = \scan_3_.curr_instr [10] | \scan_3_.curr_instr [11];
  assign N967 = \scan_3_.curr_instr [9] | N966;
  assign N968 = \scan_3_.curr_instr [8] | N967;
  assign N969 = N965 | N968;
  assign N970 = ~N969;
  assign N971 = ~\scan_3_.curr_instr [9];
  assign N972 = \scan_3_.curr_instr [10] | \scan_3_.curr_instr [11];
  assign N973 = N971 | N972;
  assign N974 = \scan_3_.curr_instr [8] | N973;
  assign N975 = N965 | N974;
  assign N976 = ~N975;
  assign \scan_3_.is_link_dest  = N970 | N976;
  assign N977 = ~\scan_3_.curr_instr [15];
  assign N978 = \scan_3_.curr_instr [18] | \scan_3_.curr_instr [19];
  assign N979 = \scan_3_.curr_instr [17] | N978;
  assign N980 = \scan_3_.curr_instr [16] | N979;
  assign N981 = N977 | N980;
  assign N982 = ~N981;
  assign N983 = ~\scan_3_.curr_instr [17];
  assign N984 = \scan_3_.curr_instr [18] | \scan_3_.curr_instr [19];
  assign N985 = N983 | N984;
  assign N986 = \scan_3_.curr_instr [16] | N985;
  assign N987 = N977 | N986;
  assign N988 = ~N987;
  assign \scan_3_.is_link_src  = N982 | N988;
  assign N989 = \scan_3_.curr_instr [11:7] == \scan_3_.curr_instr [19:15];
  assign N990 = ~\scan_3_.curr_instr [14];
  assign N991 = \scan_3_.curr_instr [30] | \scan_3_.curr_instr [31];
  assign N992 = \scan_3_.curr_instr [29] | N991;
  assign N993 = \scan_3_.curr_instr [28] | N992;
  assign N994 = \scan_3_.curr_instr [27] | N993;
  assign N995 = \scan_3_.curr_instr [26] | N994;
  assign N996 = \scan_3_.curr_instr [25] | N995;
  assign N997 = \scan_3_.curr_instr [24] | N996;
  assign N998 = \scan_3_.curr_instr [23] | N997;
  assign N999 = \scan_3_.curr_instr [22] | N998;
  assign N1000 = \scan_3_.curr_instr [21] | N999;
  assign N1001 = \scan_3_.curr_instr [20] | N1000;
  assign N1002 = \scan_3_.curr_instr [19] | N1001;
  assign N1003 = \scan_3_.curr_instr [18] | N1002;
  assign N1004 = \scan_3_.curr_instr [17] | N1003;
  assign N1005 = \scan_3_.curr_instr [16] | N1004;
  assign N1006 = N977 | N1005;
  assign N1007 = N990 | N1006;
  assign N1008 = \scan_3_.curr_instr [13] | N1007;
  assign N1009 = \scan_3_.curr_instr [1] | N1008;
  assign N1010 = N938 | N1009;
  assign N1011 = ~N1010;
  assign N1012 = ~\scan_3_.curr_instr [13];
  assign N1013 = \scan_3_.curr_instr [30] | \scan_3_.curr_instr [31];
  assign N1014 = \scan_3_.curr_instr [29] | N1013;
  assign N1015 = \scan_3_.curr_instr [28] | N1014;
  assign N1016 = \scan_3_.curr_instr [27] | N1015;
  assign N1017 = \scan_3_.curr_instr [26] | N1016;
  assign N1018 = \scan_3_.curr_instr [25] | N1017;
  assign N1019 = \scan_3_.curr_instr [24] | N1018;
  assign N1020 = \scan_3_.curr_instr [23] | N1019;
  assign N1021 = \scan_3_.curr_instr [22] | N1020;
  assign N1022 = \scan_3_.curr_instr [21] | N1021;
  assign N1023 = \scan_3_.curr_instr [20] | N1022;
  assign N1024 = \scan_3_.curr_instr [19] | N1023;
  assign N1025 = \scan_3_.curr_instr [18] | N1024;
  assign N1026 = \scan_3_.curr_instr [17] | N1025;
  assign N1027 = \scan_3_.curr_instr [16] | N1026;
  assign N1028 = N977 | N1027;
  assign N1029 = N990 | N1028;
  assign N1030 = N1012 | N1029;
  assign N1031 = \scan_3_.curr_instr [1] | N1030;
  assign N1032 = N938 | N1031;
  assign N1033 = ~N1032;
  assign N1034 = N1011 | N1033;
  assign N1035 = \scan_3_.curr_instr [30] | \scan_3_.curr_instr [31];
  assign N1036 = \scan_3_.curr_instr [29] | N1035;
  assign N1037 = \scan_3_.curr_instr [28] | N1036;
  assign N1038 = \scan_3_.curr_instr [27] | N1037;
  assign N1039 = \scan_3_.curr_instr [26] | N1038;
  assign N1040 = \scan_3_.curr_instr [25] | N1039;
  assign N1041 = \scan_3_.curr_instr [24] | N1040;
  assign N1042 = \scan_3_.curr_instr [23] | N1041;
  assign N1043 = \scan_3_.curr_instr [22] | N1042;
  assign N1044 = \scan_3_.curr_instr [21] | N1043;
  assign N1045 = \scan_3_.curr_instr [20] | N1044;
  assign N1046 = \scan_3_.curr_instr [19] | N1045;
  assign N1047 = \scan_3_.curr_instr [18] | N1046;
  assign N1048 = \scan_3_.curr_instr [17] | N1047;
  assign N1049 = \scan_3_.curr_instr [16] | N1048;
  assign N1050 = N977 | N1049;
  assign N1051 = \scan_3_.curr_instr [14] | N1050;
  assign N1052 = N1012 | N1051;
  assign N1053 = \scan_3_.curr_instr [1] | N1052;
  assign N1054 = N938 | N1053;
  assign N1055 = ~N1054;
  assign N1056 = \scan_3_.curr_instr [30] | \scan_3_.curr_instr [31];
  assign N1057 = \scan_3_.curr_instr [29] | N1056;
  assign N1058 = \scan_3_.curr_instr [28] | N1057;
  assign N1059 = \scan_3_.curr_instr [27] | N1058;
  assign N1060 = \scan_3_.curr_instr [26] | N1059;
  assign N1061 = \scan_3_.curr_instr [25] | N1060;
  assign N1062 = \scan_3_.curr_instr [24] | N1061;
  assign N1063 = \scan_3_.curr_instr [23] | N1062;
  assign N1064 = \scan_3_.curr_instr [22] | N1063;
  assign N1065 = \scan_3_.curr_instr [21] | N1064;
  assign N1066 = \scan_3_.curr_instr [20] | N1065;
  assign N1067 = \scan_3_.curr_instr [19] | N1066;
  assign N1068 = \scan_3_.curr_instr [18] | N1067;
  assign N1069 = \scan_3_.curr_instr [17] | N1068;
  assign N1070 = \scan_3_.curr_instr [16] | N1069;
  assign N1071 = N977 | N1070;
  assign N1072 = \scan_3_.curr_instr [14] | N1071;
  assign N1073 = \scan_3_.curr_instr [13] | N1072;
  assign N1074 = \scan_3_.curr_instr [12] | N1073;
  assign N1075 = \scan_3_.curr_instr [6] | N1074;
  assign N1076 = \scan_3_.curr_instr [5] | N1075;
  assign N1077 = \scan_3_.curr_instr [4] | N1076;
  assign N1078 = \scan_3_.curr_instr [3] | N1077;
  assign N1079 = \scan_3_.curr_instr [2] | N1078;
  assign N1080 = N937 | N1079;
  assign N1081 = \scan_3_.curr_instr [0] | N1080;
  assign N1082 = ~N1081;
  assign N1083 = ~\scan_3_.curr_instr [12];
  assign N1084 = \scan_3_.curr_instr [30] | \scan_3_.curr_instr [31];
  assign N1085 = \scan_3_.curr_instr [29] | N1084;
  assign N1086 = \scan_3_.curr_instr [28] | N1085;
  assign N1087 = \scan_3_.curr_instr [27] | N1086;
  assign N1088 = \scan_3_.curr_instr [26] | N1087;
  assign N1089 = \scan_3_.curr_instr [25] | N1088;
  assign N1090 = \scan_3_.curr_instr [24] | N1089;
  assign N1091 = \scan_3_.curr_instr [23] | N1090;
  assign N1092 = \scan_3_.curr_instr [22] | N1091;
  assign N1093 = \scan_3_.curr_instr [21] | N1092;
  assign N1094 = \scan_3_.curr_instr [20] | N1093;
  assign N1095 = \scan_3_.curr_instr [19] | N1094;
  assign N1096 = \scan_3_.curr_instr [18] | N1095;
  assign N1097 = \scan_3_.curr_instr [17] | N1096;
  assign N1098 = \scan_3_.curr_instr [16] | N1097;
  assign N1099 = N977 | N1098;
  assign N1100 = \scan_3_.curr_instr [14] | N1099;
  assign N1101 = \scan_3_.curr_instr [13] | N1100;
  assign N1102 = N1083 | N1101;
  assign N1103 = \scan_3_.curr_instr [6] | N1102;
  assign N1104 = \scan_3_.curr_instr [5] | N1103;
  assign N1105 = \scan_3_.curr_instr [4] | N1104;
  assign N1106 = \scan_3_.curr_instr [3] | N1105;
  assign N1107 = \scan_3_.curr_instr [2] | N1106;
  assign N1108 = N937 | N1107;
  assign N1109 = \scan_3_.curr_instr [0] | N1108;
  assign N1110 = ~N1109;
  assign N1111 = \scan_3_.curr_instr [10] | \scan_3_.curr_instr [11];
  assign N1112 = \scan_3_.curr_instr [9] | N1111;
  assign N1113 = \scan_3_.curr_instr [8] | N1112;
  assign N1114 = N965 | N1113;
  assign N1115 = ~N1114;
  assign N1116 = \scan_3_.curr_instr [10] | \scan_3_.curr_instr [11];
  assign N1117 = N971 | N1116;
  assign N1118 = \scan_3_.curr_instr [8] | N1117;
  assign N1119 = N965 | N1118;
  assign N1120 = ~N1119;
  assign \scan_3_.is_clink_src  = N1115 | N1120;
  assign N1287 = { 1'b1, 1'b0, 1'b0 } < assembled_count_i;
  assign N1290 = ~\scan_4_.curr_instr [6];
  assign N1291 = ~\scan_4_.curr_instr [5];
  assign N1292 = ~\scan_4_.curr_instr [1];
  assign N1293 = ~\scan_4_.curr_instr [0];
  assign N1294 = N1291 | N1290;
  assign N1295 = \scan_4_.curr_instr [4] | N1294;
  assign N1296 = \scan_4_.curr_instr [3] | N1295;
  assign N1297 = \scan_4_.curr_instr [2] | N1296;
  assign N1298 = N1292 | N1297;
  assign N1299 = N1293 | N1298;
  assign N1300 = ~N1299;
  assign N1301 = ~\scan_4_.curr_instr [3];
  assign N1302 = ~\scan_4_.curr_instr [2];
  assign N1303 = N1291 | N1290;
  assign N1304 = \scan_4_.curr_instr [4] | N1303;
  assign N1305 = N1301 | N1304;
  assign N1306 = N1302 | N1305;
  assign N1307 = N1292 | N1306;
  assign N1308 = N1293 | N1307;
  assign N1309 = ~N1308;
  assign N1310 = \scan_4_.curr_instr [13] | \scan_4_.curr_instr [14];
  assign N1311 = \scan_4_.curr_instr [12] | N1310;
  assign N1312 = N1290 | N1311;
  assign N1313 = N1291 | N1312;
  assign N1314 = \scan_4_.curr_instr [4] | N1313;
  assign N1315 = \scan_4_.curr_instr [3] | N1314;
  assign N1316 = N1302 | N1315;
  assign N1317 = N1292 | N1316;
  assign N1318 = N1293 | N1317;
  assign N1319 = ~N1318;
  assign N1320 = ~\scan_4_.curr_instr [7];
  assign N1321 = \scan_4_.curr_instr [10] | \scan_4_.curr_instr [11];
  assign N1322 = \scan_4_.curr_instr [9] | N1321;
  assign N1323 = \scan_4_.curr_instr [8] | N1322;
  assign N1324 = N1320 | N1323;
  assign N1325 = ~N1324;
  assign N1326 = ~\scan_4_.curr_instr [9];
  assign N1327 = \scan_4_.curr_instr [10] | \scan_4_.curr_instr [11];
  assign N1328 = N1326 | N1327;
  assign N1329 = \scan_4_.curr_instr [8] | N1328;
  assign N1330 = N1320 | N1329;
  assign N1331 = ~N1330;
  assign \scan_4_.is_link_dest  = N1325 | N1331;
  assign N1332 = ~\scan_4_.curr_instr [15];
  assign N1333 = \scan_4_.curr_instr [18] | \scan_4_.curr_instr [19];
  assign N1334 = \scan_4_.curr_instr [17] | N1333;
  assign N1335 = \scan_4_.curr_instr [16] | N1334;
  assign N1336 = N1332 | N1335;
  assign N1337 = ~N1336;
  assign N1338 = ~\scan_4_.curr_instr [17];
  assign N1339 = \scan_4_.curr_instr [18] | \scan_4_.curr_instr [19];
  assign N1340 = N1338 | N1339;
  assign N1341 = \scan_4_.curr_instr [16] | N1340;
  assign N1342 = N1332 | N1341;
  assign N1343 = ~N1342;
  assign \scan_4_.is_link_src  = N1337 | N1343;
  assign N1344 = \scan_4_.curr_instr [11:7] == \scan_4_.curr_instr [19:15];
  assign N1345 = ~\scan_4_.curr_instr [14];
  assign N1346 = \scan_4_.curr_instr [30] | \scan_4_.curr_instr [31];
  assign N1347 = \scan_4_.curr_instr [29] | N1346;
  assign N1348 = \scan_4_.curr_instr [28] | N1347;
  assign N1349 = \scan_4_.curr_instr [27] | N1348;
  assign N1350 = \scan_4_.curr_instr [26] | N1349;
  assign N1351 = \scan_4_.curr_instr [25] | N1350;
  assign N1352 = \scan_4_.curr_instr [24] | N1351;
  assign N1353 = \scan_4_.curr_instr [23] | N1352;
  assign N1354 = \scan_4_.curr_instr [22] | N1353;
  assign N1355 = \scan_4_.curr_instr [21] | N1354;
  assign N1356 = \scan_4_.curr_instr [20] | N1355;
  assign N1357 = \scan_4_.curr_instr [19] | N1356;
  assign N1358 = \scan_4_.curr_instr [18] | N1357;
  assign N1359 = \scan_4_.curr_instr [17] | N1358;
  assign N1360 = \scan_4_.curr_instr [16] | N1359;
  assign N1361 = N1332 | N1360;
  assign N1362 = N1345 | N1361;
  assign N1363 = \scan_4_.curr_instr [13] | N1362;
  assign N1364 = \scan_4_.curr_instr [1] | N1363;
  assign N1365 = N1293 | N1364;
  assign N1366 = ~N1365;
  assign N1367 = ~\scan_4_.curr_instr [13];
  assign N1368 = \scan_4_.curr_instr [30] | \scan_4_.curr_instr [31];
  assign N1369 = \scan_4_.curr_instr [29] | N1368;
  assign N1370 = \scan_4_.curr_instr [28] | N1369;
  assign N1371 = \scan_4_.curr_instr [27] | N1370;
  assign N1372 = \scan_4_.curr_instr [26] | N1371;
  assign N1373 = \scan_4_.curr_instr [25] | N1372;
  assign N1374 = \scan_4_.curr_instr [24] | N1373;
  assign N1375 = \scan_4_.curr_instr [23] | N1374;
  assign N1376 = \scan_4_.curr_instr [22] | N1375;
  assign N1377 = \scan_4_.curr_instr [21] | N1376;
  assign N1378 = \scan_4_.curr_instr [20] | N1377;
  assign N1379 = \scan_4_.curr_instr [19] | N1378;
  assign N1380 = \scan_4_.curr_instr [18] | N1379;
  assign N1381 = \scan_4_.curr_instr [17] | N1380;
  assign N1382 = \scan_4_.curr_instr [16] | N1381;
  assign N1383 = N1332 | N1382;
  assign N1384 = N1345 | N1383;
  assign N1385 = N1367 | N1384;
  assign N1386 = \scan_4_.curr_instr [1] | N1385;
  assign N1387 = N1293 | N1386;
  assign N1388 = ~N1387;
  assign N1389 = N1366 | N1388;
  assign N1390 = \scan_4_.curr_instr [30] | \scan_4_.curr_instr [31];
  assign N1391 = \scan_4_.curr_instr [29] | N1390;
  assign N1392 = \scan_4_.curr_instr [28] | N1391;
  assign N1393 = \scan_4_.curr_instr [27] | N1392;
  assign N1394 = \scan_4_.curr_instr [26] | N1393;
  assign N1395 = \scan_4_.curr_instr [25] | N1394;
  assign N1396 = \scan_4_.curr_instr [24] | N1395;
  assign N1397 = \scan_4_.curr_instr [23] | N1396;
  assign N1398 = \scan_4_.curr_instr [22] | N1397;
  assign N1399 = \scan_4_.curr_instr [21] | N1398;
  assign N1400 = \scan_4_.curr_instr [20] | N1399;
  assign N1401 = \scan_4_.curr_instr [19] | N1400;
  assign N1402 = \scan_4_.curr_instr [18] | N1401;
  assign N1403 = \scan_4_.curr_instr [17] | N1402;
  assign N1404 = \scan_4_.curr_instr [16] | N1403;
  assign N1405 = N1332 | N1404;
  assign N1406 = \scan_4_.curr_instr [14] | N1405;
  assign N1407 = N1367 | N1406;
  assign N1408 = \scan_4_.curr_instr [1] | N1407;
  assign N1409 = N1293 | N1408;
  assign N1410 = ~N1409;
  assign N1411 = \scan_4_.curr_instr [30] | \scan_4_.curr_instr [31];
  assign N1412 = \scan_4_.curr_instr [29] | N1411;
  assign N1413 = \scan_4_.curr_instr [28] | N1412;
  assign N1414 = \scan_4_.curr_instr [27] | N1413;
  assign N1415 = \scan_4_.curr_instr [26] | N1414;
  assign N1416 = \scan_4_.curr_instr [25] | N1415;
  assign N1417 = \scan_4_.curr_instr [24] | N1416;
  assign N1418 = \scan_4_.curr_instr [23] | N1417;
  assign N1419 = \scan_4_.curr_instr [22] | N1418;
  assign N1420 = \scan_4_.curr_instr [21] | N1419;
  assign N1421 = \scan_4_.curr_instr [20] | N1420;
  assign N1422 = \scan_4_.curr_instr [19] | N1421;
  assign N1423 = \scan_4_.curr_instr [18] | N1422;
  assign N1424 = \scan_4_.curr_instr [17] | N1423;
  assign N1425 = \scan_4_.curr_instr [16] | N1424;
  assign N1426 = N1332 | N1425;
  assign N1427 = \scan_4_.curr_instr [14] | N1426;
  assign N1428 = \scan_4_.curr_instr [13] | N1427;
  assign N1429 = \scan_4_.curr_instr [12] | N1428;
  assign N1430 = \scan_4_.curr_instr [6] | N1429;
  assign N1431 = \scan_4_.curr_instr [5] | N1430;
  assign N1432 = \scan_4_.curr_instr [4] | N1431;
  assign N1433 = \scan_4_.curr_instr [3] | N1432;
  assign N1434 = \scan_4_.curr_instr [2] | N1433;
  assign N1435 = N1292 | N1434;
  assign N1436 = \scan_4_.curr_instr [0] | N1435;
  assign N1437 = ~N1436;
  assign N1438 = ~\scan_4_.curr_instr [12];
  assign N1439 = \scan_4_.curr_instr [30] | \scan_4_.curr_instr [31];
  assign N1440 = \scan_4_.curr_instr [29] | N1439;
  assign N1441 = \scan_4_.curr_instr [28] | N1440;
  assign N1442 = \scan_4_.curr_instr [27] | N1441;
  assign N1443 = \scan_4_.curr_instr [26] | N1442;
  assign N1444 = \scan_4_.curr_instr [25] | N1443;
  assign N1445 = \scan_4_.curr_instr [24] | N1444;
  assign N1446 = \scan_4_.curr_instr [23] | N1445;
  assign N1447 = \scan_4_.curr_instr [22] | N1446;
  assign N1448 = \scan_4_.curr_instr [21] | N1447;
  assign N1449 = \scan_4_.curr_instr [20] | N1448;
  assign N1450 = \scan_4_.curr_instr [19] | N1449;
  assign N1451 = \scan_4_.curr_instr [18] | N1450;
  assign N1452 = \scan_4_.curr_instr [17] | N1451;
  assign N1453 = \scan_4_.curr_instr [16] | N1452;
  assign N1454 = N1332 | N1453;
  assign N1455 = \scan_4_.curr_instr [14] | N1454;
  assign N1456 = \scan_4_.curr_instr [13] | N1455;
  assign N1457 = N1438 | N1456;
  assign N1458 = \scan_4_.curr_instr [6] | N1457;
  assign N1459 = \scan_4_.curr_instr [5] | N1458;
  assign N1460 = \scan_4_.curr_instr [4] | N1459;
  assign N1461 = \scan_4_.curr_instr [3] | N1460;
  assign N1462 = \scan_4_.curr_instr [2] | N1461;
  assign N1463 = N1292 | N1462;
  assign N1464 = \scan_4_.curr_instr [0] | N1463;
  assign N1465 = ~N1464;
  assign N1466 = \scan_4_.curr_instr [10] | \scan_4_.curr_instr [11];
  assign N1467 = \scan_4_.curr_instr [9] | N1466;
  assign N1468 = \scan_4_.curr_instr [8] | N1467;
  assign N1469 = N1320 | N1468;
  assign N1470 = ~N1469;
  assign N1471 = \scan_4_.curr_instr [10] | \scan_4_.curr_instr [11];
  assign N1472 = N1326 | N1471;
  assign N1473 = \scan_4_.curr_instr [8] | N1472;
  assign N1474 = N1320 | N1473;
  assign N1475 = ~N1474;
  assign \scan_4_.is_clink_src  = N1470 | N1475;
  assign N1642 = { 1'b1, 1'b0, 1'b1 } < assembled_count_i;
  assign N1645 = ~\scan_5_.curr_instr_opcode__6_ ;
  assign N1646 = ~\scan_5_.curr_instr_opcode__5_ ;
  assign N1647 = ~\scan_5_.curr_instr_opcode__1_ ;
  assign N1648 = ~\scan_5_.curr_instr_opcode__0_ ;
  assign N1649 = N1646 | N1645;
  assign N1650 = \scan_5_.curr_instr_opcode__4_  | N1649;
  assign N1651 = \scan_5_.curr_instr_opcode__3_  | N1650;
  assign N1652 = \scan_5_.curr_instr_opcode__2_  | N1651;
  assign N1653 = N1647 | N1652;
  assign N1654 = N1648 | N1653;
  assign N1655 = ~N1654;
  assign N1656 = ~\scan_5_.curr_instr_opcode__3_ ;
  assign N1657 = ~\scan_5_.curr_instr_opcode__2_ ;
  assign N1658 = N1646 | N1645;
  assign N1659 = \scan_5_.curr_instr_opcode__4_  | N1658;
  assign N1660 = N1656 | N1659;
  assign N1661 = N1657 | N1660;
  assign N1662 = N1647 | N1661;
  assign N1663 = N1648 | N1662;
  assign N1664 = ~N1663;
  assign N1665 = \scan_5_.curr_instr_funct3__1_  | \scan_5_.curr_instr_funct3__2_ ;
  assign N1666 = \scan_5_.curr_instr_funct3__0_  | N1665;
  assign N1667 = N1645 | N1666;
  assign N1668 = N1646 | N1667;
  assign N1669 = \scan_5_.curr_instr_opcode__4_  | N1668;
  assign N1670 = \scan_5_.curr_instr_opcode__3_  | N1669;
  assign N1671 = N1657 | N1670;
  assign N1672 = N1647 | N1671;
  assign N1673 = N1648 | N1672;
  assign N1674 = ~N1673;
  assign N1675 = ~\scan_5_.curr_instr_rd_addr__0_ ;
  assign N1676 = \scan_5_.curr_instr_rd_addr__3_  | \scan_5_.curr_instr_rd_addr__4_ ;
  assign N1677 = \scan_5_.curr_instr_rd_addr__2_  | N1676;
  assign N1678 = \scan_5_.curr_instr_rd_addr__1_  | N1677;
  assign N1679 = N1675 | N1678;
  assign N1680 = ~N1679;
  assign N1681 = ~\scan_5_.curr_instr_rd_addr__2_ ;
  assign N1682 = \scan_5_.curr_instr_rd_addr__3_  | \scan_5_.curr_instr_rd_addr__4_ ;
  assign N1683 = N1681 | N1682;
  assign N1684 = \scan_5_.curr_instr_rd_addr__1_  | N1683;
  assign N1685 = N1675 | N1684;
  assign N1686 = ~N1685;
  assign \scan_5_.is_link_dest  = N1680 | N1686;
  assign N1687 = ~\scan_5_.curr_instr_rs1_addr__0_ ;
  assign N1688 = { \scan_5_.curr_instr_rd_addr__4_ , \scan_5_.curr_instr_rd_addr__3_ , \scan_5_.curr_instr_rd_addr__2_ , \scan_5_.curr_instr_rd_addr__1_ , \scan_5_.curr_instr_rd_addr__0_  } == { 1'b0, 1'b0, 1'b0, 1'b0, \scan_5_.curr_instr_rs1_addr__0_  };
  assign N1689 = ~\scan_5_.curr_instr_funct3__2_ ;
  assign N1690 = N1689 | N1687;
  assign N1691 = \scan_5_.curr_instr_funct3__1_  | N1690;
  assign N1692 = \scan_5_.curr_instr_opcode__1_  | N1691;
  assign N1693 = N1648 | N1692;
  assign N1694 = ~N1693;
  assign N1695 = ~\scan_5_.curr_instr_funct3__1_ ;
  assign N1696 = N1689 | N1687;
  assign N1697 = N1695 | N1696;
  assign N1698 = \scan_5_.curr_instr_opcode__1_  | N1697;
  assign N1699 = N1648 | N1698;
  assign N1700 = ~N1699;
  assign N1701 = N1694 | N1700;
  assign N1702 = \scan_5_.curr_instr_funct3__2_  | N1687;
  assign N1703 = N1695 | N1702;
  assign N1704 = \scan_5_.curr_instr_opcode__1_  | N1703;
  assign N1705 = N1648 | N1704;
  assign N1706 = ~N1705;
  assign N1707 = \scan_5_.curr_instr_funct3__2_  | N1687;
  assign N1708 = \scan_5_.curr_instr_funct3__1_  | N1707;
  assign N1709 = \scan_5_.curr_instr_funct3__0_  | N1708;
  assign N1710 = \scan_5_.curr_instr_opcode__6_  | N1709;
  assign N1711 = \scan_5_.curr_instr_opcode__5_  | N1710;
  assign N1712 = \scan_5_.curr_instr_opcode__4_  | N1711;
  assign N1713 = \scan_5_.curr_instr_opcode__3_  | N1712;
  assign N1714 = \scan_5_.curr_instr_opcode__2_  | N1713;
  assign N1715 = N1647 | N1714;
  assign N1716 = \scan_5_.curr_instr_opcode__0_  | N1715;
  assign N1717 = ~N1716;
  assign N1718 = ~\scan_5_.curr_instr_funct3__0_ ;
  assign N1719 = \scan_5_.curr_instr_funct3__2_  | N1687;
  assign N1720 = \scan_5_.curr_instr_funct3__1_  | N1719;
  assign N1721 = N1718 | N1720;
  assign N1722 = \scan_5_.curr_instr_opcode__6_  | N1721;
  assign N1723 = \scan_5_.curr_instr_opcode__5_  | N1722;
  assign N1724 = \scan_5_.curr_instr_opcode__4_  | N1723;
  assign N1725 = \scan_5_.curr_instr_opcode__3_  | N1724;
  assign N1726 = \scan_5_.curr_instr_opcode__2_  | N1725;
  assign N1727 = N1647 | N1726;
  assign N1728 = \scan_5_.curr_instr_opcode__0_  | N1727;
  assign N1729 = ~N1728;
  assign N1730 = \scan_5_.curr_instr_rd_addr__3_  | \scan_5_.curr_instr_rd_addr__4_ ;
  assign N1731 = \scan_5_.curr_instr_rd_addr__2_  | N1730;
  assign N1732 = \scan_5_.curr_instr_rd_addr__1_  | N1731;
  assign N1733 = N1675 | N1732;
  assign N1734 = ~N1733;
  assign N1735 = \scan_5_.curr_instr_rd_addr__3_  | \scan_5_.curr_instr_rd_addr__4_ ;
  assign N1736 = N1681 | N1735;
  assign N1737 = \scan_5_.curr_instr_rd_addr__1_  | N1736;
  assign N1738 = N1675 | N1737;
  assign N1739 = ~N1738;
  assign \scan_5_.is_clink_src  = N1734 | N1739;

  bsg_priority_encode_00000005_0
  complete_pe
  (
    .i(complete),
    .addr_o(complete_addr),
    .v_o(any_complete)
  );


  bsg_priority_encode_00000005_1
  branch_sel_pe
  (
    .i(branch[4:0]),
    .addr_o(branch_sel),
    .v_o(any_branch)
  );


  bsg_priority_encode_00000006_0
  second_branch_pe
  (
    .i(branch),
    .addr_o(last_branch_addr),
    .v_o(any_last_branch)
  );

  assign N1866 = branch_sel != last_branch_sel;

  bsg_mux_47_00000006
  branch_decode_mux
  (
    .data_i({ decode_lo_5__br_, decode_lo_5__jal_, decode_lo_5__jalr_, decode_lo_5__call_, decode_lo_5___return_, decode_lo_5__full1_, decode_lo_5__full2_, decode_lo_5__comp_, \scan_5_.imm , decode_lo_4__br_, decode_lo_4__jal_, decode_lo_4__jalr_, decode_lo_4__call_, decode_lo_4___return_, decode_lo_4__full1_, decode_lo_4__full2_, decode_lo_4__comp_, \scan_4_.imm , decode_lo_3__br_, decode_lo_3__jal_, decode_lo_3__jalr_, decode_lo_3__call_, decode_lo_3___return_, decode_lo_3__full1_, decode_lo_3__full2_, decode_lo_3__comp_, \scan_3_.imm , decode_lo_2__br_, decode_lo_2__jal_, decode_lo_2__jalr_, decode_lo_2__call_, decode_lo_2___return_, decode_lo_2__full1_, decode_lo_2__full2_, decode_lo_2__comp_, \scan_2_.imm , decode_lo_1__br_, decode_lo_1__jal_, decode_lo_1__jalr_, decode_lo_1__call_, decode_lo_1___return_, decode_lo_1__full1_, decode_lo_1__full2_, decode_lo_1__comp_, \scan_1_.imm , decode_lo_0__br_, decode_lo_0__jal_, decode_lo_0__jalr_, decode_lo_0__call_, decode_lo_0___return_, decode_lo_0__full1_, decode_lo_0__full2_, decode_lo_0__comp_, \scan_0_.imm  }),
    .sel_i(branch_sel),
    .data_o({ branch_decode_lo_br_, branch_decode_lo_jal_, branch_decode_lo_jalr_, branch_decode_lo_call_, branch_decode_lo__return_, branch_decode_lo_full1_, branch_decode_lo_full2_, branch_decode_lo_comp_, fetch_scan_o[38:0] })
  );


  bsg_mux_47_00000006
  next_decode_mux
  (
    .data_i({ decode_lo_5__br_, decode_lo_5__jal_, decode_lo_5__jalr_, decode_lo_5__call_, decode_lo_5___return_, decode_lo_5__full1_, decode_lo_5__full2_, decode_lo_5__comp_, \scan_5_.imm , decode_lo_4__br_, decode_lo_4__jal_, decode_lo_4__jalr_, decode_lo_4__call_, decode_lo_4___return_, decode_lo_4__full1_, decode_lo_4__full2_, decode_lo_4__comp_, \scan_4_.imm , decode_lo_3__br_, decode_lo_3__jal_, decode_lo_3__jalr_, decode_lo_3__call_, decode_lo_3___return_, decode_lo_3__full1_, decode_lo_3__full2_, decode_lo_3__comp_, \scan_3_.imm , decode_lo_2__br_, decode_lo_2__jal_, decode_lo_2__jalr_, decode_lo_2__call_, decode_lo_2___return_, decode_lo_2__full1_, decode_lo_2__full2_, decode_lo_2__comp_, \scan_2_.imm , decode_lo_1__br_, decode_lo_1__jal_, decode_lo_1__jalr_, decode_lo_1__call_, decode_lo_1___return_, decode_lo_1__full1_, decode_lo_1__full2_, decode_lo_1__comp_, \scan_1_.imm , decode_lo_0__br_, decode_lo_0__jal_, decode_lo_0__jalr_, decode_lo_0__call_, decode_lo_0___return_, decode_lo_0__full1_, decode_lo_0__full2_, decode_lo_0__comp_, \scan_0_.imm  }),
    .sel_i(next_sel),
    .data_o(next_decode_lo)
  );

  assign N1873 = assembled_count_i > branch_count;
  assign N1874 = assembled_count_i > branch_count;
  assign N1875 = assembled_count_i > linear_count;
  assign N1882 = linear_count[1] | linear_count[2];
  assign N1883 = linear_count[0] | N1882;
  assign N1884 = ~N1883;
  assign N1885 = \scan_5_.curr_instr_rd_addr__3_  | \scan_5_.curr_instr_rd_addr__4_ ;
  assign N1886 = \scan_5_.curr_instr_rd_addr__2_  | N1885;
  assign N1887 = \scan_5_.curr_instr_rd_addr__1_  | N1886;
  assign N1888 = N1675 | N1887;
  assign N1889 = ~N1888;
  assign N1890 = \scan_4_.curr_instr [10] | \scan_4_.curr_instr [11];
  assign N1891 = \scan_4_.curr_instr [9] | N1890;
  assign N1892 = \scan_4_.curr_instr [8] | N1891;
  assign N1893 = N1320 | N1892;
  assign N1894 = ~N1893;
  assign N1895 = \scan_3_.curr_instr [10] | \scan_3_.curr_instr [11];
  assign N1896 = \scan_3_.curr_instr [9] | N1895;
  assign N1897 = \scan_3_.curr_instr [8] | N1896;
  assign N1898 = N965 | N1897;
  assign N1899 = ~N1898;
  assign N1900 = \scan_2_.curr_instr [10] | \scan_2_.curr_instr [11];
  assign N1901 = \scan_2_.curr_instr [9] | N1900;
  assign N1902 = \scan_2_.curr_instr [8] | N1901;
  assign N1903 = N610 | N1902;
  assign N1904 = ~N1903;
  assign N1905 = \scan_1_.curr_instr [10] | \scan_1_.curr_instr [11];
  assign N1906 = \scan_1_.curr_instr [9] | N1905;
  assign N1907 = \scan_1_.curr_instr [8] | N1906;
  assign N1908 = N334 | N1907;
  assign N1909 = ~N1908;
  assign N1910 = \scan_0_.curr_instr [10] | \scan_0_.curr_instr [11];
  assign N1911 = \scan_0_.curr_instr [9] | N1910;
  assign N1912 = \scan_0_.curr_instr [8] | N1911;
  assign N1913 = N58 | N1912;
  assign N1914 = ~N1913;
  assign linear_sel = { 1'b1, 1'b0, 1'b0 } - complete_addr;
  assign last_branch_sel = { 1'b1, 1'b0, 1'b1 } - last_branch_addr;
  assign { N1869, N1868, N1867 } = branch_sel + 1'b1;
  assign { N1865, N1864, N1863 } = branch_sel + 1'b1;
  assign { N1861, N1860, N1859 } = linear_sel + 1'b1;
  assign { N1872, N1871, N1870 } = linear_sel + 1'b1;
  assign fetch_scan_o[82:79] = linear_count + 1'b1;
  assign { N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217 } = { \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [7:7], \scan_0_.curr_instr [30:25], \scan_0_.curr_instr [11:8], 1'b0 } + { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 };
  assign { N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257 } = { \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [31:31], \scan_0_.curr_instr [19:12], \scan_0_.curr_instr [20:20], \scan_0_.curr_instr [30:21], 1'b0 } + { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 };
  assign { N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769 } = { \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [7:7], \scan_2_.curr_instr [30:25], \scan_2_.curr_instr [11:8], 1'b0 } + { 1'b1, 1'b0 };
  assign { N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809 } = { \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [31:31], \scan_2_.curr_instr [19:12], \scan_2_.curr_instr [20:20], \scan_2_.curr_instr [30:21], 1'b0 } + { 1'b1, 1'b0 };
  assign { N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124 } = { \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [7:7], \scan_3_.curr_instr [30:25], \scan_3_.curr_instr [11:8], 1'b0 } + { 1'b1, 1'b0, 1'b0 };
  assign { N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164 } = { \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [31:31], \scan_3_.curr_instr [19:12], \scan_3_.curr_instr [20:20], \scan_3_.curr_instr [30:21], 1'b0 } + { 1'b1, 1'b0, 1'b0 };
  assign { N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479 } = { \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [7:7], \scan_4_.curr_instr [30:25], \scan_4_.curr_instr [11:8], 1'b0 } + { 1'b1, 1'b1, 1'b0 };
  assign { N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533 } = { \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [6:5], \scan_1_.curr_instr [2:2], \scan_1_.curr_instr [11:10], \scan_1_.curr_instr [4:3], 1'b0 } + { 1'b1, 1'b0 };
  assign { N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494 } = { \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [12:12], \scan_1_.curr_instr [8:8], \scan_1_.curr_instr [10:9], \scan_1_.curr_instr [6:6], \scan_1_.curr_instr [7:7], \scan_1_.curr_instr [2:2], \scan_1_.curr_instr [11:11], \scan_1_.curr_instr [5:3], 1'b0 } + { 1'b1, 1'b0 };
  assign { N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519 } = { \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [31:31], \scan_4_.curr_instr [19:12], \scan_4_.curr_instr [20:20], \scan_4_.curr_instr [30:21], 1'b0 } + { 1'b1, 1'b1, 1'b0 };
  assign { N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743 } = { \scan_5_.curr_instr_rd_addr__0_ , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \scan_5_.curr_instr_rd_addr__4_ , \scan_5_.curr_instr_rd_addr__3_ , \scan_5_.curr_instr_rd_addr__2_ , \scan_5_.curr_instr_rd_addr__1_ , 1'b0 } + { 1'b1, 1'b0, 1'b0, 1'b0 };
  assign { N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888 } = { \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [6:5], \scan_2_.curr_instr [2:2], \scan_2_.curr_instr [11:10], \scan_2_.curr_instr [4:3], 1'b0 } + { 1'b1, 1'b0, 1'b0 };
  assign { N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849 } = { \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [12:12], \scan_2_.curr_instr [8:8], \scan_2_.curr_instr [10:9], \scan_2_.curr_instr [6:6], \scan_2_.curr_instr [7:7], \scan_2_.curr_instr [2:2], \scan_2_.curr_instr [11:11], \scan_2_.curr_instr [5:3], 1'b0 } + { 1'b1, 1'b0, 1'b0 };
  assign { N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757 } = { \scan_5_.curr_instr_rs1_addr__0_ , \scan_5_.curr_instr_funct3__2_ , \scan_5_.curr_instr_funct3__1_ , \scan_5_.curr_instr_funct3__0_ , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } + { 1'b1, 1'b0, 1'b0, 1'b0 };
  assign { N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243 } = { \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [6:5], \scan_3_.curr_instr [2:2], \scan_3_.curr_instr [11:10], \scan_3_.curr_instr [4:3], 1'b0 } + { 1'b1, 1'b1, 1'b0 };
  assign { N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204 } = { \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [12:12], \scan_3_.curr_instr [8:8], \scan_3_.curr_instr [10:9], \scan_3_.curr_instr [6:6], \scan_3_.curr_instr [7:7], \scan_3_.curr_instr [2:2], \scan_3_.curr_instr [11:11], \scan_3_.curr_instr [5:3], 1'b0 } + { 1'b1, 1'b1, 1'b0 };
  assign { N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598 } = { \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [6:5], \scan_4_.curr_instr [2:2], \scan_4_.curr_instr [11:10], \scan_4_.curr_instr [4:3], 1'b0 } + { 1'b1, 1'b0, 1'b0, 1'b0 };
  assign { N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559 } = { \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [12:12], \scan_4_.curr_instr [8:8], \scan_4_.curr_instr [10:9], \scan_4_.curr_instr [6:6], \scan_4_.curr_instr [7:7], \scan_4_.curr_instr [2:2], \scan_4_.curr_instr [11:11], \scan_4_.curr_instr [5:3], 1'b0 } + { 1'b1, 1'b0, 1'b0, 1'b0 };
  assign { N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814 } = { \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_opcode__6_ , \scan_5_.curr_instr_opcode__5_ , \scan_5_.curr_instr_opcode__2_ , \scan_5_.curr_instr_rd_addr__4_ , \scan_5_.curr_instr_rd_addr__3_ , \scan_5_.curr_instr_opcode__4_ , \scan_5_.curr_instr_opcode__3_ , 1'b0 } + { 1'b1, 1'b0, 1'b1, 1'b0 };
  assign { N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775 } = { \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_rd_addr__1_ , \scan_5_.curr_instr_rd_addr__3_ , \scan_5_.curr_instr_rd_addr__2_ , \scan_5_.curr_instr_opcode__6_ , \scan_5_.curr_instr_rd_addr__0_ , \scan_5_.curr_instr_opcode__2_ , \scan_5_.curr_instr_rd_addr__4_ , \scan_5_.curr_instr_opcode__5_ , \scan_5_.curr_instr_opcode__4_ , \scan_5_.curr_instr_opcode__3_ , 1'b0 } + { 1'b1, 1'b0, 1'b1, 1'b0 };
  assign \scan_0_.curr_instr  = (N0)? { fetch_instr_o[15:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fetch_instr_o[15:0] } : 1'b0;
  assign N0 = N27;
  assign N1 = N26;
  assign \scan_0_.imm  = (N2)? { N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217 } : 
                         (N297)? { N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257 } : 
                         (N300)? { \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [8:8], \scan_0_.curr_instr [10:9], \scan_0_.curr_instr [6:6], \scan_0_.curr_instr [7:7], \scan_0_.curr_instr [2:2], \scan_0_.curr_instr [11:11], \scan_0_.curr_instr [5:3], 1'b0 } : 
                         (N216)? { \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [12:12], \scan_0_.curr_instr [6:5], \scan_0_.curr_instr [2:2], \scan_0_.curr_instr [11:10], \scan_0_.curr_instr [4:3], 1'b0 } : 1'b0;
  assign N2 = \scan_0_.is_br ;
  assign \scan_1_.curr_instr  = (N3)? fetch_instr_o[31:0] : 
                                (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fetch_instr_o[31:16] } : 1'b0;
  assign N3 = N303;
  assign N4 = N302;
  assign \scan_1_.imm  = (N5)? { \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [7:7], \scan_1_.curr_instr [30:25], \scan_1_.curr_instr [11:8], 1'b0 } : 
                         (N573)? { \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [31:31], \scan_1_.curr_instr [19:12], \scan_1_.curr_instr [20:20], \scan_1_.curr_instr [30:21], 1'b0 } : 
                         (N576)? { N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494 } : 
                         (N492)? { N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533 } : 1'b0;
  assign N5 = \scan_1_.is_br ;
  assign \scan_2_.curr_instr  = (N6)? fetch_instr_o[47:16] : 
                                (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fetch_instr_o[47:32] } : 1'b0;
  assign N6 = N579;
  assign N7 = N578;
  assign \scan_2_.imm  = (N8)? { N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769 } : 
                         (N928)? { N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809 } : 
                         (N931)? { N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849 } : 
                         (N768)? { N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888 } : 1'b0;
  assign N8 = \scan_2_.is_br ;
  assign \scan_3_.curr_instr  = (N9)? fetch_instr_o[63:32] : 
                                (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fetch_instr_o[63:48] } : 1'b0;
  assign N9 = N934;
  assign N10 = N933;
  assign \scan_3_.imm  = (N11)? { N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124 } : 
                         (N1283)? { N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164 } : 
                         (N1286)? { N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204 } : 
                         (N1123)? { N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243 } : 1'b0;
  assign N11 = \scan_3_.is_br ;
  assign \scan_4_.curr_instr  = (N12)? fetch_instr_o[79:48] : 
                                (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fetch_instr_o[79:64] } : 1'b0;
  assign N12 = N1289;
  assign N13 = N1288;
  assign \scan_4_.imm  = (N14)? { N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479 } : 
                         (N1638)? { N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519 } : 
                         (N1641)? { N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559 } : 
                         (N1478)? { N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598 } : 1'b0;
  assign N14 = \scan_4_.is_br ;
  assign { \scan_5_.curr_instr_rs1_addr__0_ , \scan_5_.curr_instr_funct3__2_ , \scan_5_.curr_instr_funct3__1_ , \scan_5_.curr_instr_funct3__0_ , \scan_5_.curr_instr_rd_addr__4_ , \scan_5_.curr_instr_rd_addr__3_ , \scan_5_.curr_instr_rd_addr__2_ , \scan_5_.curr_instr_rd_addr__1_ , \scan_5_.curr_instr_rd_addr__0_ , \scan_5_.curr_instr_opcode__6_ , \scan_5_.curr_instr_opcode__5_ , \scan_5_.curr_instr_opcode__4_ , \scan_5_.curr_instr_opcode__3_ , \scan_5_.curr_instr_opcode__2_ , \scan_5_.curr_instr_opcode__1_ , \scan_5_.curr_instr_opcode__0_  } = (N15)? fetch_instr_o[79:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = N1644;
  assign N16 = N1643;
  assign \scan_5_.imm  = (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743 } : 
                         (N1854)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757 } : 
                         (N1857)? { N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775 } : 
                         (N1742)? { N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814 } : 1'b0;
  assign N17 = \scan_5_.is_br ;
  assign linear_count = (N18)? { N1861, N1860, N1859 } : 
                        (N19)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N18 = any_complete;
  assign N19 = N1858;
  assign branch_count = (N20)? { N1865, N1864, N1863 } : 
                        (N21)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N20 = any_branch;
  assign N21 = N1862;
  assign next_sel = (N20)? { N1869, N1868, N1867 } : 
                    (N21)? { N1872, N1871, N1870 } : 1'b0;
  assign fetch_scan_o[42:40] = (N18)? next_sel : 
                               (N19)? { 1'b0, 1'b0, 1'b1 } : 1'b0;
  assign fetch_scan_o[121:117] = (N22)? { branch_decode_lo_br_, branch_decode_lo_jal_, branch_decode_lo_jalr_, branch_decode_lo_call_, branch_decode_lo__return_ } : 
                                 (N23)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N22 = assembled_yumi_o;
  assign N23 = N1876;
  assign fetch_count_o = (N20)? branch_count : 
                         (N21)? linear_count : 1'b0;
  assign { N1881, N1880, N1879 } = (N24)? assembled_count_i : 
                                   (N1878)? branch_count : 1'b0;
  assign N24 = N1877;
  assign assembled_count_o = (N20)? { N1881, N1880, N1879 } : 
                             (N21)? linear_count : 1'b0;
  assign decode_lo_0__full1_ = N1915 & full1_0_;
  assign N1915 = fetch_v_o & N25;
  assign decode_lo_0__full2_ = N1916 & 1'b0;
  assign N1916 = fetch_v_o & N25;
  assign decode_lo_0__comp_ = N1917 & N1920;
  assign N1917 = fetch_v_o & N25;
  assign N1920 = N1918 & N1919;
  assign N1918 = ~full1_0_;
  assign N1919 = ~1'b0;
  assign N26 = ~decode_lo_0__full2_;
  assign N27 = decode_lo_0__full2_;
  assign \scan_0_.is_br  = decode_lo_0__full2_ & N38;
  assign \scan_0_.is_jal  = decode_lo_0__full2_ & N47;
  assign \scan_0_.is_jalr  = decode_lo_0__full2_ & N57;
  assign \scan_0_.is_link_match  = N1921 & N82;
  assign N1921 = \scan_0_.is_link_src  & \scan_0_.is_link_dest ;
  assign \scan_0_.is_call  = N1922 & \scan_0_.is_link_dest ;
  assign N1922 = \scan_0_.is_jal  | \scan_0_.is_jalr ;
  assign \scan_0_.is_return  = N1923 & N1924;
  assign N1923 = \scan_0_.is_jalr  & \scan_0_.is_link_src ;
  assign N1924 = ~\scan_0_.is_link_match ;
  assign \scan_0_.is_cbr  = decode_lo_0__comp_ & N127;
  assign \scan_0_.is_cj  = decode_lo_0__comp_ & N148;
  assign \scan_0_.is_cjr  = decode_lo_0__comp_ & N175;
  assign \scan_0_.is_cjalr  = decode_lo_0__comp_ & N203;
  assign \scan_0_.is_clink_match  = N1925 & N1914;
  assign N1925 = \scan_0_.is_clink_src  & \scan_0_.is_cjalr ;
  assign \scan_0_.is_ccall  = N1927 & \scan_0_.is_cjalr ;
  assign N1927 = N1926 | \scan_0_.is_cjalr ;
  assign N1926 = \scan_0_.is_cj  | \scan_0_.is_cjr ;
  assign \scan_0_.is_creturn  = N1929 & N1930;
  assign N1929 = N1928 & \scan_0_.is_clink_src ;
  assign N1928 = \scan_0_.is_cjr  | \scan_0_.is_cjalr ;
  assign N1930 = ~\scan_0_.is_clink_match ;
  assign N214 = \scan_0_.is_jal  | \scan_0_.is_br ;
  assign N215 = \scan_0_.is_cj  | N214;
  assign N216 = ~N215;
  assign N256 = N297;
  assign N296 = ~\scan_0_.is_br ;
  assign N297 = \scan_0_.is_jal  & N296;
  assign N298 = ~\scan_0_.is_jal ;
  assign N299 = N296 & N298;
  assign N300 = \scan_0_.is_cj  & N299;
  assign full1_0_ = N1931 & N1919;
  assign N1931 = \scan_0_.curr_instr [1] & \scan_0_.curr_instr [0];
  assign branch[0] = N1936 | \scan_0_.is_cjalr ;
  assign N1936 = N1935 | \scan_0_.is_cjr ;
  assign N1935 = N1934 | \scan_0_.is_cj ;
  assign N1934 = N1933 | \scan_0_.is_cbr ;
  assign N1933 = N1932 | \scan_0_.is_jalr ;
  assign N1932 = \scan_0_.is_br  | \scan_0_.is_jal ;
  assign complete[0] = decode_lo_0__comp_ | decode_lo_0__full2_;
  assign decode_lo_0__br_ = \scan_0_.is_br  | \scan_0_.is_cbr ;
  assign decode_lo_0__jal_ = \scan_0_.is_jal  | \scan_0_.is_cj ;
  assign decode_lo_0__jalr_ = N1937 | \scan_0_.is_cjalr ;
  assign N1937 = \scan_0_.is_jalr  | \scan_0_.is_cjr ;
  assign decode_lo_0__call_ = \scan_0_.is_call  | \scan_0_.is_ccall ;
  assign decode_lo_0___return_ = \scan_0_.is_return  | \scan_0_.is_creturn ;
  assign decode_lo_1__full1_ = N1938 & full1_1_;
  assign N1938 = fetch_v_o & N301;
  assign decode_lo_1__full2_ = N1939 & full1_0_;
  assign N1939 = fetch_v_o & N301;
  assign decode_lo_1__comp_ = N1940 & N1942;
  assign N1940 = fetch_v_o & N301;
  assign N1942 = N1941 & N1918;
  assign N1941 = ~full1_1_;
  assign N302 = ~decode_lo_1__full2_;
  assign N303 = decode_lo_1__full2_;
  assign \scan_1_.is_br  = decode_lo_1__full2_ & N314;
  assign \scan_1_.is_jal  = decode_lo_1__full2_ & N323;
  assign \scan_1_.is_jalr  = decode_lo_1__full2_ & N333;
  assign \scan_1_.is_link_match  = N1943 & N358;
  assign N1943 = \scan_1_.is_link_src  & \scan_1_.is_link_dest ;
  assign \scan_1_.is_call  = N1944 & \scan_1_.is_link_dest ;
  assign N1944 = \scan_1_.is_jal  | \scan_1_.is_jalr ;
  assign \scan_1_.is_return  = N1945 & N1946;
  assign N1945 = \scan_1_.is_jalr  & \scan_1_.is_link_src ;
  assign N1946 = ~\scan_1_.is_link_match ;
  assign \scan_1_.is_cbr  = decode_lo_1__comp_ & N403;
  assign \scan_1_.is_cj  = decode_lo_1__comp_ & N424;
  assign \scan_1_.is_cjr  = decode_lo_1__comp_ & N451;
  assign \scan_1_.is_cjalr  = decode_lo_1__comp_ & N479;
  assign \scan_1_.is_clink_match  = N1947 & N1909;
  assign N1947 = \scan_1_.is_clink_src  & \scan_1_.is_cjalr ;
  assign \scan_1_.is_ccall  = N1949 & \scan_1_.is_cjalr ;
  assign N1949 = N1948 | \scan_1_.is_cjalr ;
  assign N1948 = \scan_1_.is_cj  | \scan_1_.is_cjr ;
  assign \scan_1_.is_creturn  = N1951 & N1952;
  assign N1951 = N1950 & \scan_1_.is_clink_src ;
  assign N1950 = \scan_1_.is_cjr  | \scan_1_.is_cjalr ;
  assign N1952 = ~\scan_1_.is_clink_match ;
  assign N490 = \scan_1_.is_jal  | \scan_1_.is_br ;
  assign N491 = \scan_1_.is_cj  | N490;
  assign N492 = ~N491;
  assign N493 = N576;
  assign N572 = ~\scan_1_.is_br ;
  assign N573 = \scan_1_.is_jal  & N572;
  assign N574 = ~\scan_1_.is_jal ;
  assign N575 = N572 & N574;
  assign N576 = \scan_1_.is_cj  & N575;
  assign full1_1_ = N1953 & N1918;
  assign N1953 = \scan_1_.curr_instr [1] & \scan_1_.curr_instr [0];
  assign branch[1] = N1958 | \scan_1_.is_cjalr ;
  assign N1958 = N1957 | \scan_1_.is_cjr ;
  assign N1957 = N1956 | \scan_1_.is_cj ;
  assign N1956 = N1955 | \scan_1_.is_cbr ;
  assign N1955 = N1954 | \scan_1_.is_jalr ;
  assign N1954 = \scan_1_.is_br  | \scan_1_.is_jal ;
  assign complete[1] = decode_lo_1__comp_ | decode_lo_1__full2_;
  assign decode_lo_1__br_ = \scan_1_.is_br  | \scan_1_.is_cbr ;
  assign decode_lo_1__jal_ = \scan_1_.is_jal  | \scan_1_.is_cj ;
  assign decode_lo_1__jalr_ = N1959 | \scan_1_.is_cjalr ;
  assign N1959 = \scan_1_.is_jalr  | \scan_1_.is_cjr ;
  assign decode_lo_1__call_ = \scan_1_.is_call  | \scan_1_.is_ccall ;
  assign decode_lo_1___return_ = \scan_1_.is_return  | \scan_1_.is_creturn ;
  assign decode_lo_2__full1_ = N1960 & full1_2_;
  assign N1960 = fetch_v_o & N577;
  assign decode_lo_2__full2_ = N1961 & full1_1_;
  assign N1961 = fetch_v_o & N577;
  assign decode_lo_2__comp_ = N1962 & N1964;
  assign N1962 = fetch_v_o & N577;
  assign N1964 = N1963 & N1941;
  assign N1963 = ~full1_2_;
  assign N578 = ~decode_lo_2__full2_;
  assign N579 = decode_lo_2__full2_;
  assign \scan_2_.is_br  = decode_lo_2__full2_ & N590;
  assign \scan_2_.is_jal  = decode_lo_2__full2_ & N599;
  assign \scan_2_.is_jalr  = decode_lo_2__full2_ & N609;
  assign \scan_2_.is_link_match  = N1965 & N634;
  assign N1965 = \scan_2_.is_link_src  & \scan_2_.is_link_dest ;
  assign \scan_2_.is_call  = N1966 & \scan_2_.is_link_dest ;
  assign N1966 = \scan_2_.is_jal  | \scan_2_.is_jalr ;
  assign \scan_2_.is_return  = N1967 & N1968;
  assign N1967 = \scan_2_.is_jalr  & \scan_2_.is_link_src ;
  assign N1968 = ~\scan_2_.is_link_match ;
  assign \scan_2_.is_cbr  = decode_lo_2__comp_ & N679;
  assign \scan_2_.is_cj  = decode_lo_2__comp_ & N700;
  assign \scan_2_.is_cjr  = decode_lo_2__comp_ & N727;
  assign \scan_2_.is_cjalr  = decode_lo_2__comp_ & N755;
  assign \scan_2_.is_clink_match  = N1969 & N1904;
  assign N1969 = \scan_2_.is_clink_src  & \scan_2_.is_cjalr ;
  assign \scan_2_.is_ccall  = N1971 & \scan_2_.is_cjalr ;
  assign N1971 = N1970 | \scan_2_.is_cjalr ;
  assign N1970 = \scan_2_.is_cj  | \scan_2_.is_cjr ;
  assign \scan_2_.is_creturn  = N1973 & N1974;
  assign N1973 = N1972 & \scan_2_.is_clink_src ;
  assign N1972 = \scan_2_.is_cjr  | \scan_2_.is_cjalr ;
  assign N1974 = ~\scan_2_.is_clink_match ;
  assign N766 = \scan_2_.is_jal  | \scan_2_.is_br ;
  assign N767 = \scan_2_.is_cj  | N766;
  assign N768 = ~N767;
  assign N808 = N928;
  assign N848 = N931;
  assign N927 = ~\scan_2_.is_br ;
  assign N928 = \scan_2_.is_jal  & N927;
  assign N929 = ~\scan_2_.is_jal ;
  assign N930 = N927 & N929;
  assign N931 = \scan_2_.is_cj  & N930;
  assign full1_2_ = N1975 & N1941;
  assign N1975 = \scan_2_.curr_instr [1] & \scan_2_.curr_instr [0];
  assign branch[2] = N1980 | \scan_2_.is_cjalr ;
  assign N1980 = N1979 | \scan_2_.is_cjr ;
  assign N1979 = N1978 | \scan_2_.is_cj ;
  assign N1978 = N1977 | \scan_2_.is_cbr ;
  assign N1977 = N1976 | \scan_2_.is_jalr ;
  assign N1976 = \scan_2_.is_br  | \scan_2_.is_jal ;
  assign complete[2] = decode_lo_2__comp_ | decode_lo_2__full2_;
  assign decode_lo_2__br_ = \scan_2_.is_br  | \scan_2_.is_cbr ;
  assign decode_lo_2__jal_ = \scan_2_.is_jal  | \scan_2_.is_cj ;
  assign decode_lo_2__jalr_ = N1981 | \scan_2_.is_cjalr ;
  assign N1981 = \scan_2_.is_jalr  | \scan_2_.is_cjr ;
  assign decode_lo_2__call_ = \scan_2_.is_call  | \scan_2_.is_ccall ;
  assign decode_lo_2___return_ = \scan_2_.is_return  | \scan_2_.is_creturn ;
  assign decode_lo_3__full1_ = N1982 & full1_3_;
  assign N1982 = fetch_v_o & N932;
  assign decode_lo_3__full2_ = N1983 & full1_2_;
  assign N1983 = fetch_v_o & N932;
  assign decode_lo_3__comp_ = N1984 & N1986;
  assign N1984 = fetch_v_o & N932;
  assign N1986 = N1985 & N1963;
  assign N1985 = ~full1_3_;
  assign N933 = ~decode_lo_3__full2_;
  assign N934 = decode_lo_3__full2_;
  assign \scan_3_.is_br  = decode_lo_3__full2_ & N945;
  assign \scan_3_.is_jal  = decode_lo_3__full2_ & N954;
  assign \scan_3_.is_jalr  = decode_lo_3__full2_ & N964;
  assign \scan_3_.is_link_match  = N1987 & N989;
  assign N1987 = \scan_3_.is_link_src  & \scan_3_.is_link_dest ;
  assign \scan_3_.is_call  = N1988 & \scan_3_.is_link_dest ;
  assign N1988 = \scan_3_.is_jal  | \scan_3_.is_jalr ;
  assign \scan_3_.is_return  = N1989 & N1990;
  assign N1989 = \scan_3_.is_jalr  & \scan_3_.is_link_src ;
  assign N1990 = ~\scan_3_.is_link_match ;
  assign \scan_3_.is_cbr  = decode_lo_3__comp_ & N1034;
  assign \scan_3_.is_cj  = decode_lo_3__comp_ & N1055;
  assign \scan_3_.is_cjr  = decode_lo_3__comp_ & N1082;
  assign \scan_3_.is_cjalr  = decode_lo_3__comp_ & N1110;
  assign \scan_3_.is_clink_match  = N1991 & N1899;
  assign N1991 = \scan_3_.is_clink_src  & \scan_3_.is_cjalr ;
  assign \scan_3_.is_ccall  = N1993 & \scan_3_.is_cjalr ;
  assign N1993 = N1992 | \scan_3_.is_cjalr ;
  assign N1992 = \scan_3_.is_cj  | \scan_3_.is_cjr ;
  assign \scan_3_.is_creturn  = N1995 & N1996;
  assign N1995 = N1994 & \scan_3_.is_clink_src ;
  assign N1994 = \scan_3_.is_cjr  | \scan_3_.is_cjalr ;
  assign N1996 = ~\scan_3_.is_clink_match ;
  assign N1121 = \scan_3_.is_jal  | \scan_3_.is_br ;
  assign N1122 = \scan_3_.is_cj  | N1121;
  assign N1123 = ~N1122;
  assign N1163 = N1283;
  assign N1203 = N1286;
  assign N1282 = ~\scan_3_.is_br ;
  assign N1283 = \scan_3_.is_jal  & N1282;
  assign N1284 = ~\scan_3_.is_jal ;
  assign N1285 = N1282 & N1284;
  assign N1286 = \scan_3_.is_cj  & N1285;
  assign full1_3_ = N1997 & N1963;
  assign N1997 = \scan_3_.curr_instr [1] & \scan_3_.curr_instr [0];
  assign branch[3] = N2002 | \scan_3_.is_cjalr ;
  assign N2002 = N2001 | \scan_3_.is_cjr ;
  assign N2001 = N2000 | \scan_3_.is_cj ;
  assign N2000 = N1999 | \scan_3_.is_cbr ;
  assign N1999 = N1998 | \scan_3_.is_jalr ;
  assign N1998 = \scan_3_.is_br  | \scan_3_.is_jal ;
  assign complete[3] = decode_lo_3__comp_ | decode_lo_3__full2_;
  assign decode_lo_3__br_ = \scan_3_.is_br  | \scan_3_.is_cbr ;
  assign decode_lo_3__jal_ = \scan_3_.is_jal  | \scan_3_.is_cj ;
  assign decode_lo_3__jalr_ = N2003 | \scan_3_.is_cjalr ;
  assign N2003 = \scan_3_.is_jalr  | \scan_3_.is_cjr ;
  assign decode_lo_3__call_ = \scan_3_.is_call  | \scan_3_.is_ccall ;
  assign decode_lo_3___return_ = \scan_3_.is_return  | \scan_3_.is_creturn ;
  assign decode_lo_4__full1_ = N2004 & full1_4_;
  assign N2004 = fetch_v_o & N1287;
  assign decode_lo_4__full2_ = N2005 & full1_3_;
  assign N2005 = fetch_v_o & N1287;
  assign decode_lo_4__comp_ = N2006 & N2008;
  assign N2006 = fetch_v_o & N1287;
  assign N2008 = N2007 & N1985;
  assign N2007 = ~full1_4_;
  assign N1288 = ~decode_lo_4__full2_;
  assign N1289 = decode_lo_4__full2_;
  assign \scan_4_.is_br  = decode_lo_4__full2_ & N1300;
  assign \scan_4_.is_jal  = decode_lo_4__full2_ & N1309;
  assign \scan_4_.is_jalr  = decode_lo_4__full2_ & N1319;
  assign \scan_4_.is_link_match  = N2009 & N1344;
  assign N2009 = \scan_4_.is_link_src  & \scan_4_.is_link_dest ;
  assign \scan_4_.is_call  = N2010 & \scan_4_.is_link_dest ;
  assign N2010 = \scan_4_.is_jal  | \scan_4_.is_jalr ;
  assign \scan_4_.is_return  = N2011 & N2012;
  assign N2011 = \scan_4_.is_jalr  & \scan_4_.is_link_src ;
  assign N2012 = ~\scan_4_.is_link_match ;
  assign \scan_4_.is_cbr  = decode_lo_4__comp_ & N1389;
  assign \scan_4_.is_cj  = decode_lo_4__comp_ & N1410;
  assign \scan_4_.is_cjr  = decode_lo_4__comp_ & N1437;
  assign \scan_4_.is_cjalr  = decode_lo_4__comp_ & N1465;
  assign \scan_4_.is_clink_match  = N2013 & N1894;
  assign N2013 = \scan_4_.is_clink_src  & \scan_4_.is_cjalr ;
  assign \scan_4_.is_ccall  = N2015 & \scan_4_.is_cjalr ;
  assign N2015 = N2014 | \scan_4_.is_cjalr ;
  assign N2014 = \scan_4_.is_cj  | \scan_4_.is_cjr ;
  assign \scan_4_.is_creturn  = N2017 & N2018;
  assign N2017 = N2016 & \scan_4_.is_clink_src ;
  assign N2016 = \scan_4_.is_cjr  | \scan_4_.is_cjalr ;
  assign N2018 = ~\scan_4_.is_clink_match ;
  assign N1476 = \scan_4_.is_jal  | \scan_4_.is_br ;
  assign N1477 = \scan_4_.is_cj  | N1476;
  assign N1478 = ~N1477;
  assign N1518 = N1638;
  assign N1558 = N1641;
  assign N1637 = ~\scan_4_.is_br ;
  assign N1638 = \scan_4_.is_jal  & N1637;
  assign N1639 = ~\scan_4_.is_jal ;
  assign N1640 = N1637 & N1639;
  assign N1641 = \scan_4_.is_cj  & N1640;
  assign full1_4_ = N2019 & N1985;
  assign N2019 = \scan_4_.curr_instr [1] & \scan_4_.curr_instr [0];
  assign branch[4] = N2024 | \scan_4_.is_cjalr ;
  assign N2024 = N2023 | \scan_4_.is_cjr ;
  assign N2023 = N2022 | \scan_4_.is_cj ;
  assign N2022 = N2021 | \scan_4_.is_cbr ;
  assign N2021 = N2020 | \scan_4_.is_jalr ;
  assign N2020 = \scan_4_.is_br  | \scan_4_.is_jal ;
  assign complete[4] = decode_lo_4__comp_ | decode_lo_4__full2_;
  assign decode_lo_4__br_ = \scan_4_.is_br  | \scan_4_.is_cbr ;
  assign decode_lo_4__jal_ = \scan_4_.is_jal  | \scan_4_.is_cj ;
  assign decode_lo_4__jalr_ = N2025 | \scan_4_.is_cjalr ;
  assign N2025 = \scan_4_.is_jalr  | \scan_4_.is_cjr ;
  assign decode_lo_4__call_ = \scan_4_.is_call  | \scan_4_.is_ccall ;
  assign decode_lo_4___return_ = \scan_4_.is_return  | \scan_4_.is_creturn ;
  assign decode_lo_5__full1_ = N2026 & full1_5_;
  assign N2026 = fetch_v_o & N1642;
  assign decode_lo_5__full2_ = N2027 & full1_4_;
  assign N2027 = fetch_v_o & N1642;
  assign decode_lo_5__comp_ = N2028 & N2030;
  assign N2028 = fetch_v_o & N1642;
  assign N2030 = N2029 & N2007;
  assign N2029 = ~full1_5_;
  assign N1643 = ~decode_lo_5__full2_;
  assign N1644 = decode_lo_5__full2_;
  assign \scan_5_.is_br  = decode_lo_5__full2_ & N1655;
  assign \scan_5_.is_jal  = decode_lo_5__full2_ & N1664;
  assign \scan_5_.is_jalr  = decode_lo_5__full2_ & N1674;
  assign \scan_5_.is_link_match  = N2031 & N1688;
  assign N2031 = \scan_5_.curr_instr_rs1_addr__0_  & \scan_5_.is_link_dest ;
  assign \scan_5_.is_call  = N2032 & \scan_5_.is_link_dest ;
  assign N2032 = \scan_5_.is_jal  | \scan_5_.is_jalr ;
  assign \scan_5_.is_return  = N2033 & N2034;
  assign N2033 = \scan_5_.is_jalr  & \scan_5_.curr_instr_rs1_addr__0_ ;
  assign N2034 = ~\scan_5_.is_link_match ;
  assign \scan_5_.is_cbr  = decode_lo_5__comp_ & N1701;
  assign \scan_5_.is_cj  = decode_lo_5__comp_ & N1706;
  assign \scan_5_.is_cjr  = decode_lo_5__comp_ & N1717;
  assign \scan_5_.is_cjalr  = decode_lo_5__comp_ & N1729;
  assign \scan_5_.is_clink_match  = N2035 & N1889;
  assign N2035 = \scan_5_.is_clink_src  & \scan_5_.is_cjalr ;
  assign \scan_5_.is_ccall  = N2037 & \scan_5_.is_cjalr ;
  assign N2037 = N2036 | \scan_5_.is_cjalr ;
  assign N2036 = \scan_5_.is_cj  | \scan_5_.is_cjr ;
  assign \scan_5_.is_creturn  = N2039 & N2040;
  assign N2039 = N2038 & \scan_5_.is_clink_src ;
  assign N2038 = \scan_5_.is_cjr  | \scan_5_.is_cjalr ;
  assign N2040 = ~\scan_5_.is_clink_match ;
  assign N1740 = \scan_5_.is_jal  | \scan_5_.is_br ;
  assign N1741 = \scan_5_.is_cj  | N1740;
  assign N1742 = ~N1741;
  assign N1756 = N1854;
  assign N1774 = N1857;
  assign N1853 = ~\scan_5_.is_br ;
  assign N1854 = \scan_5_.is_jal  & N1853;
  assign N1855 = ~\scan_5_.is_jal ;
  assign N1856 = N1853 & N1855;
  assign N1857 = \scan_5_.is_cj  & N1856;
  assign full1_5_ = N2041 & N2007;
  assign N2041 = \scan_5_.curr_instr_opcode__1_  & \scan_5_.curr_instr_opcode__0_ ;
  assign branch[5] = N2046 | \scan_5_.is_cjalr ;
  assign N2046 = N2045 | \scan_5_.is_cjr ;
  assign N2045 = N2044 | \scan_5_.is_cj ;
  assign N2044 = N2043 | \scan_5_.is_cbr ;
  assign N2043 = N2042 | \scan_5_.is_jalr ;
  assign N2042 = \scan_5_.is_br  | \scan_5_.is_jal ;
  assign decode_lo_5__br_ = \scan_5_.is_br  | \scan_5_.is_cbr ;
  assign decode_lo_5__jal_ = \scan_5_.is_jal  | \scan_5_.is_cj ;
  assign decode_lo_5__jalr_ = N2047 | \scan_5_.is_cjalr ;
  assign N2047 = \scan_5_.is_jalr  | \scan_5_.is_cjr ;
  assign decode_lo_5__call_ = \scan_5_.is_call  | \scan_5_.is_ccall ;
  assign decode_lo_5___return_ = \scan_5_.is_return  | \scan_5_.is_creturn ;
  assign N1858 = ~any_complete;
  assign N1862 = ~any_branch;
  assign double_branch = any_branch & N1866;
  assign assembled_startup = N2049 & N1884;
  assign N2049 = N1862 & N2048;
  assign N2048 = ~fetch_taken_i;
  assign assembled_catchup = N2051 & N2052;
  assign N2051 = N2050 & N1873;
  assign N2050 = any_branch & N2048;
  assign N2052 = ~double_branch;
  assign assembled_rebase = N2054 & double_branch;
  assign N2054 = N2053 & N1874;
  assign N2053 = any_branch & N2048;
  assign assembled_linear = N1862 & N1875;
  assign N1876 = ~assembled_yumi_o;
  assign fetch_startup_o = assembled_yumi_o & assembled_startup;
  assign fetch_catchup_o = assembled_yumi_o & assembled_catchup;
  assign fetch_rebase_o = assembled_yumi_o & assembled_rebase;
  assign fetch_linear_o = assembled_yumi_o & assembled_linear;
  assign N1877 = assembled_rebase | fetch_taken_i;
  assign N1878 = ~N1877;

endmodule



module bsg_dff_reset_en_width_p3
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [2:0] data_i;
  output [2:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [2:0] data_o;
  wire N0,N1,N2;
  reg data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bp_fe_controller_00
(
  clk_i,
  reset_i,
  pc_gen_init_done_i,
  fe_cmd_i,
  fe_cmd_v_i,
  fe_cmd_yumi_o,
  fe_queue_o,
  fe_queue_v_o,
  fe_queue_ready_and_i,
  redirect_v_o,
  redirect_pc_o,
  redirect_npc_o,
  redirect_instr_o,
  redirect_resume_o,
  redirect_br_v_o,
  redirect_br_taken_o,
  redirect_br_ntaken_o,
  redirect_br_nonbr_o,
  redirect_br_metadata_fwd_o,
  attaboy_v_o,
  attaboy_force_o,
  attaboy_pc_o,
  attaboy_taken_o,
  attaboy_ntaken_o,
  attaboy_br_metadata_fwd_o,
  attaboy_yumi_i,
  next_pc_i,
  ovr_i,
  tl_flush_o,
  tv_we_i,
  itlb_miss_tl_i,
  instr_page_fault_tl_i,
  instr_access_fault_tl_i,
  icache_miss_tv_i,
  tv_flush_o,
  fetch_v_i,
  fetch_pc_i,
  fetch_instr_i,
  fetch_count_i,
  fetch_partial_i,
  fetch_br_metadata_fwd_i,
  fetch_yumi_o,
  itlb_r_v_o,
  itlb_w_v_o,
  itlb_w_vtag_o,
  itlb_w_entry_o,
  itlb_fence_v_o,
  icache_v_o,
  icache_force_o,
  icache_pkt_o,
  icache_yumi_i,
  shadow_priv_w_o,
  shadow_priv_o,
  shadow_translation_en_w_o,
  shadow_translation_en_o
);

  input [113:0] fe_cmd_i;
  output [173:0] fe_queue_o;
  output [38:0] redirect_pc_o;
  output [38:0] redirect_npc_o;
  output [15:0] redirect_instr_o;
  output [48:0] redirect_br_metadata_fwd_o;
  output [38:0] attaboy_pc_o;
  output [48:0] attaboy_br_metadata_fwd_o;
  input [38:0] next_pc_i;
  input [38:0] fetch_pc_i;
  input [79:0] fetch_instr_i;
  input [2:0] fetch_count_i;
  input [48:0] fetch_br_metadata_fwd_i;
  output [26:0] itlb_w_vtag_o;
  output [35:0] itlb_w_entry_o;
  output [71:0] icache_pkt_o;
  output [1:0] shadow_priv_o;
  input clk_i;
  input reset_i;
  input pc_gen_init_done_i;
  input fe_cmd_v_i;
  input fe_queue_ready_and_i;
  input attaboy_yumi_i;
  input ovr_i;
  input tv_we_i;
  input itlb_miss_tl_i;
  input instr_page_fault_tl_i;
  input instr_access_fault_tl_i;
  input icache_miss_tv_i;
  input fetch_v_i;
  input fetch_partial_i;
  input icache_yumi_i;
  output fe_cmd_yumi_o;
  output fe_queue_v_o;
  output redirect_v_o;
  output redirect_resume_o;
  output redirect_br_v_o;
  output redirect_br_taken_o;
  output redirect_br_ntaken_o;
  output redirect_br_nonbr_o;
  output attaboy_v_o;
  output attaboy_force_o;
  output attaboy_taken_o;
  output attaboy_ntaken_o;
  output tl_flush_o;
  output tv_flush_o;
  output fetch_yumi_o;
  output itlb_r_v_o;
  output itlb_w_v_o;
  output itlb_fence_v_o;
  output icache_v_o;
  output icache_force_o;
  output shadow_priv_w_o;
  output shadow_translation_en_w_o;
  output shadow_translation_en_o;
  wire [173:0] fe_queue_o;
  wire [38:0] redirect_pc_o,redirect_npc_o,attaboy_pc_o;
  wire [15:0] redirect_instr_o;
  wire [48:0] redirect_br_metadata_fwd_o,attaboy_br_metadata_fwd_o;
  wire [26:0] itlb_w_vtag_o;
  wire [35:0] itlb_w_entry_o;
  wire [71:0] icache_pkt_o;
  wire [1:0] shadow_priv_o,state_r,state_n;
  wire fe_cmd_yumi_o,fe_queue_v_o,redirect_v_o,redirect_resume_o,redirect_br_v_o,
  redirect_br_taken_o,redirect_br_ntaken_o,redirect_br_nonbr_o,attaboy_v_o,
  attaboy_force_o,attaboy_taken_o,attaboy_ntaken_o,tl_flush_o,tv_flush_o,fetch_yumi_o,
  itlb_r_v_o,itlb_w_v_o,itlb_fence_v_o,icache_v_o,icache_force_o,shadow_priv_w_o,
  shadow_translation_en_w_o,shadow_translation_en_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,
  fe_cmd_i_17_,fe_queue_o_173_,fe_queue_o_172_,fe_queue_o_171_,fe_queue_o_170_,
  fe_queue_o_169_,fe_queue_o_168_,fe_queue_o_167_,fe_queue_o_166_,fe_queue_o_165_,
  fe_queue_o_164_,fe_queue_o_163_,fe_queue_o_162_,fe_queue_o_161_,fe_queue_o_160_,
  fe_queue_o_159_,fe_queue_o_158_,fe_queue_o_157_,fe_queue_o_156_,fe_queue_o_155_,
  fe_queue_o_154_,fe_queue_o_153_,fe_queue_o_152_,fe_queue_o_151_,fe_queue_o_150_,
  fe_queue_o_149_,fe_queue_o_148_,fe_queue_o_147_,fe_queue_o_146_,fe_queue_o_145_,
  fe_queue_o_144_,fe_queue_o_143_,fe_queue_o_142_,fe_queue_o_141_,fe_queue_o_140_,
  fe_queue_o_139_,fe_queue_o_138_,fe_queue_o_137_,fe_queue_o_136_,fe_queue_o_135_,
  fe_queue_o_134_,fe_queue_o_133_,fe_queue_o_132_,fe_queue_o_131_,fe_queue_o_130_,
  fe_queue_o_129_,fe_queue_o_128_,fe_queue_o_127_,fe_queue_o_126_,fe_queue_o_125_,
  fe_queue_o_124_,fe_queue_o_123_,fe_queue_o_122_,fe_queue_o_121_,fe_queue_o_120_,
  fe_queue_o_119_,fe_queue_o_118_,fe_queue_o_117_,fe_queue_o_116_,fe_queue_o_115_,
  fe_queue_o_114_,fe_queue_o_113_,fe_queue_o_112_,fe_queue_o_111_,fe_queue_o_110_,
  fe_queue_o_109_,fe_queue_o_108_,fe_queue_o_107_,fe_queue_o_106_,fe_queue_o_105_,
  fe_queue_o_104_,fe_queue_o_103_,fe_queue_o_102_,fe_queue_o_101_,fe_queue_o_100_,
  fe_queue_o_99_,fe_queue_o_98_,fe_queue_o_97_,fe_queue_o_96_,fe_queue_o_95_,
  fe_queue_o_94_,fe_queue_o_93_,fe_queue_o_92_,fe_queue_o_91_,fe_queue_o_90_,fe_queue_o_89_,
  fe_queue_o_88_,fe_queue_o_87_,fe_queue_o_86_,fe_queue_o_85_,fe_queue_o_84_,
  fe_queue_o_83_,fe_queue_o_82_,fe_queue_o_81_,fe_queue_o_80_,fe_queue_o_79_,
  fe_queue_o_78_,fe_queue_o_77_,fe_queue_o_76_,fe_queue_o_75_,fe_queue_o_74_,fe_queue_o_73_,
  fe_queue_o_72_,fe_queue_o_71_,fe_queue_o_70_,fe_queue_o_69_,fe_queue_o_68_,
  fe_queue_o_67_,fe_queue_o_66_,fe_queue_o_65_,fe_queue_o_64_,fe_queue_o_63_,
  fe_queue_o_62_,fe_queue_o_61_,fe_queue_o_60_,fe_queue_o_59_,fe_queue_o_58_,fe_queue_o_57_,
  fe_queue_o_56_,fe_queue_o_55_,fe_queue_o_54_,fe_queue_o_53_,fe_queue_o_52_,
  fe_queue_o_51_,fe_queue_o_50_,fe_queue_o_49_,fe_queue_o_48_,fe_queue_o_47_,
  fe_queue_o_46_,fe_queue_o_45_,fe_queue_o_44_,fe_queue_o_43_,fe_queue_o_42_,fe_queue_o_41_,
  fe_queue_o_40_,fe_queue_o_39_,fe_queue_o_38_,fe_queue_o_37_,fe_queue_o_36_,
  fe_queue_o_35_,fe_queue_o_34_,fe_queue_o_33_,fe_queue_o_32_,fe_queue_o_31_,
  fe_queue_o_30_,fe_queue_o_29_,fe_queue_o_28_,fe_queue_o_27_,fe_queue_o_26_,fe_queue_o_25_,
  fe_queue_o_24_,fe_queue_o_23_,fe_queue_o_22_,fe_queue_o_21_,fe_queue_o_20_,
  fe_queue_o_19_,fe_queue_o_18_,fe_queue_o_17_,fe_queue_o_16_,fe_queue_o_15_,
  fe_queue_o_14_,fe_queue_o_13_,fe_queue_o_12_,fe_queue_o_11_,fe_queue_o_10_,fe_queue_o_9_,
  fe_queue_o_8_,fe_queue_o_7_,fe_queue_o_6_,attaboy_br_metadata_fwd_o_48_,
  attaboy_br_metadata_fwd_o_47_,itlb_w_entry_o_35_,icache_pkt_o_71_,icache_pkt_o_70_,
  icache_pkt_o_69_,icache_pkt_o_68_,icache_pkt_o_67_,icache_pkt_o_66_,icache_pkt_o_65_,
  icache_pkt_o_64_,icache_pkt_o_63_,icache_pkt_o_62_,icache_pkt_o_61_,icache_pkt_o_60_,
  icache_pkt_o_59_,icache_pkt_o_58_,icache_pkt_o_57_,icache_pkt_o_56_,
  icache_pkt_o_55_,icache_pkt_o_54_,icache_pkt_o_53_,icache_pkt_o_52_,icache_pkt_o_51_,
  icache_pkt_o_50_,icache_pkt_o_49_,icache_pkt_o_48_,icache_pkt_o_47_,icache_pkt_o_46_,
  icache_pkt_o_45_,icache_pkt_o_44_,icache_pkt_o_43_,icache_pkt_o_42_,
  icache_pkt_o_41_,icache_pkt_o_40_,icache_pkt_o_39_,icache_pkt_o_38_,icache_pkt_o_37_,
  icache_pkt_o_36_,icache_pkt_o_35_,icache_pkt_o_34_,icache_pkt_o_33_,pc_redirect_v,
  icache_fill_response_v,icache_fence_v,state_reset_v,itlb_fill_response_v,itlb_fence_v,
  wait_v,br_miss_v,eret_v,interrupt_v,trap_v,translation_v,cmd_nonattaboy_v,
  cmd_immediate_v,cmd_complex_v,N11,N12,N13,N14,N15,N16,N17,N18,N19,_0_net_,
  itlb_miss_tv_r,instr_page_fault_tv_r,instr_access_fault_tv_r,if2_exception_v,N20,
  fetch_instr_v,fetch_exception_v,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,
  N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,
  N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,
  N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,
  N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,
  N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,
  N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143;
  reg state_r_1_sv2v_reg,state_r_0_sv2v_reg;
  assign state_r[1] = state_r_1_sv2v_reg;
  assign state_r[0] = state_r_0_sv2v_reg;
  assign icache_pkt_o[2] = 1'b0;
  assign icache_pkt_o[3] = 1'b0;
  assign icache_pkt_o[4] = 1'b0;
  assign icache_pkt_o[5] = 1'b0;
  assign icache_pkt_o[6] = 1'b0;
  assign icache_pkt_o[7] = 1'b0;
  assign icache_pkt_o[8] = 1'b0;
  assign icache_pkt_o[9] = 1'b0;
  assign icache_pkt_o[10] = 1'b0;
  assign icache_pkt_o[11] = 1'b0;
  assign icache_pkt_o[12] = 1'b0;
  assign icache_pkt_o[13] = 1'b0;
  assign icache_pkt_o[14] = 1'b0;
  assign icache_pkt_o[15] = 1'b0;
  assign icache_pkt_o[16] = 1'b0;
  assign icache_pkt_o[17] = 1'b0;
  assign icache_pkt_o[18] = 1'b0;
  assign icache_pkt_o[19] = 1'b0;
  assign icache_pkt_o[20] = 1'b0;
  assign icache_pkt_o[21] = 1'b0;
  assign icache_pkt_o[22] = 1'b0;
  assign icache_pkt_o[23] = 1'b0;
  assign icache_pkt_o[24] = 1'b0;
  assign icache_pkt_o[25] = 1'b0;
  assign icache_pkt_o[26] = 1'b0;
  assign icache_pkt_o[27] = 1'b0;
  assign icache_pkt_o[28] = 1'b0;
  assign icache_pkt_o[29] = 1'b0;
  assign icache_pkt_o[30] = 1'b0;
  assign icache_pkt_o[31] = 1'b0;
  assign icache_pkt_o[32] = 1'b0;
  assign fe_cmd_i_17_ = fe_cmd_i[17];
  assign shadow_translation_en_o = fe_cmd_i_17_;
  assign fe_queue_o_173_ = fetch_pc_i[38];
  assign fe_queue_o[173] = fe_queue_o_173_;
  assign fe_queue_o_172_ = fetch_pc_i[37];
  assign fe_queue_o[172] = fe_queue_o_172_;
  assign fe_queue_o_171_ = fetch_pc_i[36];
  assign fe_queue_o[171] = fe_queue_o_171_;
  assign fe_queue_o_170_ = fetch_pc_i[35];
  assign fe_queue_o[170] = fe_queue_o_170_;
  assign fe_queue_o_169_ = fetch_pc_i[34];
  assign fe_queue_o[169] = fe_queue_o_169_;
  assign fe_queue_o_168_ = fetch_pc_i[33];
  assign fe_queue_o[168] = fe_queue_o_168_;
  assign fe_queue_o_167_ = fetch_pc_i[32];
  assign fe_queue_o[167] = fe_queue_o_167_;
  assign fe_queue_o_166_ = fetch_pc_i[31];
  assign fe_queue_o[166] = fe_queue_o_166_;
  assign fe_queue_o_165_ = fetch_pc_i[30];
  assign fe_queue_o[165] = fe_queue_o_165_;
  assign fe_queue_o_164_ = fetch_pc_i[29];
  assign fe_queue_o[164] = fe_queue_o_164_;
  assign fe_queue_o_163_ = fetch_pc_i[28];
  assign fe_queue_o[163] = fe_queue_o_163_;
  assign fe_queue_o_162_ = fetch_pc_i[27];
  assign fe_queue_o[162] = fe_queue_o_162_;
  assign fe_queue_o_161_ = fetch_pc_i[26];
  assign fe_queue_o[161] = fe_queue_o_161_;
  assign fe_queue_o_160_ = fetch_pc_i[25];
  assign fe_queue_o[160] = fe_queue_o_160_;
  assign fe_queue_o_159_ = fetch_pc_i[24];
  assign fe_queue_o[159] = fe_queue_o_159_;
  assign fe_queue_o_158_ = fetch_pc_i[23];
  assign fe_queue_o[158] = fe_queue_o_158_;
  assign fe_queue_o_157_ = fetch_pc_i[22];
  assign fe_queue_o[157] = fe_queue_o_157_;
  assign fe_queue_o_156_ = fetch_pc_i[21];
  assign fe_queue_o[156] = fe_queue_o_156_;
  assign fe_queue_o_155_ = fetch_pc_i[20];
  assign fe_queue_o[155] = fe_queue_o_155_;
  assign fe_queue_o_154_ = fetch_pc_i[19];
  assign fe_queue_o[154] = fe_queue_o_154_;
  assign fe_queue_o_153_ = fetch_pc_i[18];
  assign fe_queue_o[153] = fe_queue_o_153_;
  assign fe_queue_o_152_ = fetch_pc_i[17];
  assign fe_queue_o[152] = fe_queue_o_152_;
  assign fe_queue_o_151_ = fetch_pc_i[16];
  assign fe_queue_o[151] = fe_queue_o_151_;
  assign fe_queue_o_150_ = fetch_pc_i[15];
  assign fe_queue_o[150] = fe_queue_o_150_;
  assign fe_queue_o_149_ = fetch_pc_i[14];
  assign fe_queue_o[149] = fe_queue_o_149_;
  assign fe_queue_o_148_ = fetch_pc_i[13];
  assign fe_queue_o[148] = fe_queue_o_148_;
  assign fe_queue_o_147_ = fetch_pc_i[12];
  assign fe_queue_o[147] = fe_queue_o_147_;
  assign fe_queue_o_146_ = fetch_pc_i[11];
  assign fe_queue_o[146] = fe_queue_o_146_;
  assign fe_queue_o_145_ = fetch_pc_i[10];
  assign fe_queue_o[145] = fe_queue_o_145_;
  assign fe_queue_o_144_ = fetch_pc_i[9];
  assign fe_queue_o[144] = fe_queue_o_144_;
  assign fe_queue_o_143_ = fetch_pc_i[8];
  assign fe_queue_o[143] = fe_queue_o_143_;
  assign fe_queue_o_142_ = fetch_pc_i[7];
  assign fe_queue_o[142] = fe_queue_o_142_;
  assign fe_queue_o_141_ = fetch_pc_i[6];
  assign fe_queue_o[141] = fe_queue_o_141_;
  assign fe_queue_o_140_ = fetch_pc_i[5];
  assign fe_queue_o[140] = fe_queue_o_140_;
  assign fe_queue_o_139_ = fetch_pc_i[4];
  assign fe_queue_o[139] = fe_queue_o_139_;
  assign fe_queue_o_138_ = fetch_pc_i[3];
  assign fe_queue_o[138] = fe_queue_o_138_;
  assign fe_queue_o_137_ = fetch_pc_i[2];
  assign fe_queue_o[137] = fe_queue_o_137_;
  assign fe_queue_o_136_ = fetch_pc_i[1];
  assign fe_queue_o[136] = fe_queue_o_136_;
  assign fe_queue_o_135_ = fetch_pc_i[0];
  assign fe_queue_o[135] = fe_queue_o_135_;
  assign fe_queue_o_134_ = fetch_instr_i[79];
  assign fe_queue_o[134] = fe_queue_o_134_;
  assign fe_queue_o_133_ = fetch_instr_i[78];
  assign fe_queue_o[133] = fe_queue_o_133_;
  assign fe_queue_o_132_ = fetch_instr_i[77];
  assign fe_queue_o[132] = fe_queue_o_132_;
  assign fe_queue_o_131_ = fetch_instr_i[76];
  assign fe_queue_o[131] = fe_queue_o_131_;
  assign fe_queue_o_130_ = fetch_instr_i[75];
  assign fe_queue_o[130] = fe_queue_o_130_;
  assign fe_queue_o_129_ = fetch_instr_i[74];
  assign fe_queue_o[129] = fe_queue_o_129_;
  assign fe_queue_o_128_ = fetch_instr_i[73];
  assign fe_queue_o[128] = fe_queue_o_128_;
  assign fe_queue_o_127_ = fetch_instr_i[72];
  assign fe_queue_o[127] = fe_queue_o_127_;
  assign fe_queue_o_126_ = fetch_instr_i[71];
  assign fe_queue_o[126] = fe_queue_o_126_;
  assign fe_queue_o_125_ = fetch_instr_i[70];
  assign fe_queue_o[125] = fe_queue_o_125_;
  assign fe_queue_o_124_ = fetch_instr_i[69];
  assign fe_queue_o[124] = fe_queue_o_124_;
  assign fe_queue_o_123_ = fetch_instr_i[68];
  assign fe_queue_o[123] = fe_queue_o_123_;
  assign fe_queue_o_122_ = fetch_instr_i[67];
  assign fe_queue_o[122] = fe_queue_o_122_;
  assign fe_queue_o_121_ = fetch_instr_i[66];
  assign fe_queue_o[121] = fe_queue_o_121_;
  assign fe_queue_o_120_ = fetch_instr_i[65];
  assign fe_queue_o[120] = fe_queue_o_120_;
  assign fe_queue_o_119_ = fetch_instr_i[64];
  assign fe_queue_o[119] = fe_queue_o_119_;
  assign fe_queue_o_118_ = fetch_instr_i[63];
  assign fe_queue_o[118] = fe_queue_o_118_;
  assign fe_queue_o_117_ = fetch_instr_i[62];
  assign fe_queue_o[117] = fe_queue_o_117_;
  assign fe_queue_o_116_ = fetch_instr_i[61];
  assign fe_queue_o[116] = fe_queue_o_116_;
  assign fe_queue_o_115_ = fetch_instr_i[60];
  assign fe_queue_o[115] = fe_queue_o_115_;
  assign fe_queue_o_114_ = fetch_instr_i[59];
  assign fe_queue_o[114] = fe_queue_o_114_;
  assign fe_queue_o_113_ = fetch_instr_i[58];
  assign fe_queue_o[113] = fe_queue_o_113_;
  assign fe_queue_o_112_ = fetch_instr_i[57];
  assign fe_queue_o[112] = fe_queue_o_112_;
  assign fe_queue_o_111_ = fetch_instr_i[56];
  assign fe_queue_o[111] = fe_queue_o_111_;
  assign fe_queue_o_110_ = fetch_instr_i[55];
  assign fe_queue_o[110] = fe_queue_o_110_;
  assign fe_queue_o_109_ = fetch_instr_i[54];
  assign fe_queue_o[109] = fe_queue_o_109_;
  assign fe_queue_o_108_ = fetch_instr_i[53];
  assign fe_queue_o[108] = fe_queue_o_108_;
  assign fe_queue_o_107_ = fetch_instr_i[52];
  assign fe_queue_o[107] = fe_queue_o_107_;
  assign fe_queue_o_106_ = fetch_instr_i[51];
  assign fe_queue_o[106] = fe_queue_o_106_;
  assign fe_queue_o_105_ = fetch_instr_i[50];
  assign fe_queue_o[105] = fe_queue_o_105_;
  assign fe_queue_o_104_ = fetch_instr_i[49];
  assign fe_queue_o[104] = fe_queue_o_104_;
  assign fe_queue_o_103_ = fetch_instr_i[48];
  assign fe_queue_o[103] = fe_queue_o_103_;
  assign fe_queue_o_102_ = fetch_instr_i[47];
  assign fe_queue_o[102] = fe_queue_o_102_;
  assign fe_queue_o_101_ = fetch_instr_i[46];
  assign fe_queue_o[101] = fe_queue_o_101_;
  assign fe_queue_o_100_ = fetch_instr_i[45];
  assign fe_queue_o[100] = fe_queue_o_100_;
  assign fe_queue_o_99_ = fetch_instr_i[44];
  assign fe_queue_o[99] = fe_queue_o_99_;
  assign fe_queue_o_98_ = fetch_instr_i[43];
  assign fe_queue_o[98] = fe_queue_o_98_;
  assign fe_queue_o_97_ = fetch_instr_i[42];
  assign fe_queue_o[97] = fe_queue_o_97_;
  assign fe_queue_o_96_ = fetch_instr_i[41];
  assign fe_queue_o[96] = fe_queue_o_96_;
  assign fe_queue_o_95_ = fetch_instr_i[40];
  assign fe_queue_o[95] = fe_queue_o_95_;
  assign fe_queue_o_94_ = fetch_instr_i[39];
  assign fe_queue_o[94] = fe_queue_o_94_;
  assign fe_queue_o_93_ = fetch_instr_i[38];
  assign fe_queue_o[93] = fe_queue_o_93_;
  assign fe_queue_o_92_ = fetch_instr_i[37];
  assign fe_queue_o[92] = fe_queue_o_92_;
  assign fe_queue_o_91_ = fetch_instr_i[36];
  assign fe_queue_o[91] = fe_queue_o_91_;
  assign fe_queue_o_90_ = fetch_instr_i[35];
  assign fe_queue_o[90] = fe_queue_o_90_;
  assign fe_queue_o_89_ = fetch_instr_i[34];
  assign fe_queue_o[89] = fe_queue_o_89_;
  assign fe_queue_o_88_ = fetch_instr_i[33];
  assign fe_queue_o[88] = fe_queue_o_88_;
  assign fe_queue_o_87_ = fetch_instr_i[32];
  assign fe_queue_o[87] = fe_queue_o_87_;
  assign fe_queue_o_86_ = fetch_instr_i[31];
  assign fe_queue_o[86] = fe_queue_o_86_;
  assign fe_queue_o_85_ = fetch_instr_i[30];
  assign fe_queue_o[85] = fe_queue_o_85_;
  assign fe_queue_o_84_ = fetch_instr_i[29];
  assign fe_queue_o[84] = fe_queue_o_84_;
  assign fe_queue_o_83_ = fetch_instr_i[28];
  assign fe_queue_o[83] = fe_queue_o_83_;
  assign fe_queue_o_82_ = fetch_instr_i[27];
  assign fe_queue_o[82] = fe_queue_o_82_;
  assign fe_queue_o_81_ = fetch_instr_i[26];
  assign fe_queue_o[81] = fe_queue_o_81_;
  assign fe_queue_o_80_ = fetch_instr_i[25];
  assign fe_queue_o[80] = fe_queue_o_80_;
  assign fe_queue_o_79_ = fetch_instr_i[24];
  assign fe_queue_o[79] = fe_queue_o_79_;
  assign fe_queue_o_78_ = fetch_instr_i[23];
  assign fe_queue_o[78] = fe_queue_o_78_;
  assign fe_queue_o_77_ = fetch_instr_i[22];
  assign fe_queue_o[77] = fe_queue_o_77_;
  assign fe_queue_o_76_ = fetch_instr_i[21];
  assign fe_queue_o[76] = fe_queue_o_76_;
  assign fe_queue_o_75_ = fetch_instr_i[20];
  assign fe_queue_o[75] = fe_queue_o_75_;
  assign fe_queue_o_74_ = fetch_instr_i[19];
  assign fe_queue_o[74] = fe_queue_o_74_;
  assign fe_queue_o_73_ = fetch_instr_i[18];
  assign fe_queue_o[73] = fe_queue_o_73_;
  assign fe_queue_o_72_ = fetch_instr_i[17];
  assign fe_queue_o[72] = fe_queue_o_72_;
  assign fe_queue_o_71_ = fetch_instr_i[16];
  assign fe_queue_o[71] = fe_queue_o_71_;
  assign fe_queue_o_70_ = fetch_instr_i[15];
  assign fe_queue_o[70] = fe_queue_o_70_;
  assign fe_queue_o_69_ = fetch_instr_i[14];
  assign fe_queue_o[69] = fe_queue_o_69_;
  assign fe_queue_o_68_ = fetch_instr_i[13];
  assign fe_queue_o[68] = fe_queue_o_68_;
  assign fe_queue_o_67_ = fetch_instr_i[12];
  assign fe_queue_o[67] = fe_queue_o_67_;
  assign fe_queue_o_66_ = fetch_instr_i[11];
  assign fe_queue_o[66] = fe_queue_o_66_;
  assign fe_queue_o_65_ = fetch_instr_i[10];
  assign fe_queue_o[65] = fe_queue_o_65_;
  assign fe_queue_o_64_ = fetch_instr_i[9];
  assign fe_queue_o[64] = fe_queue_o_64_;
  assign fe_queue_o_63_ = fetch_instr_i[8];
  assign fe_queue_o[63] = fe_queue_o_63_;
  assign fe_queue_o_62_ = fetch_instr_i[7];
  assign fe_queue_o[62] = fe_queue_o_62_;
  assign fe_queue_o_61_ = fetch_instr_i[6];
  assign fe_queue_o[61] = fe_queue_o_61_;
  assign fe_queue_o_60_ = fetch_instr_i[5];
  assign fe_queue_o[60] = fe_queue_o_60_;
  assign fe_queue_o_59_ = fetch_instr_i[4];
  assign fe_queue_o[59] = fe_queue_o_59_;
  assign fe_queue_o_58_ = fetch_instr_i[3];
  assign fe_queue_o[58] = fe_queue_o_58_;
  assign fe_queue_o_57_ = fetch_instr_i[2];
  assign fe_queue_o[57] = fe_queue_o_57_;
  assign fe_queue_o_56_ = fetch_instr_i[1];
  assign fe_queue_o[56] = fe_queue_o_56_;
  assign fe_queue_o_55_ = fetch_instr_i[0];
  assign fe_queue_o[55] = fe_queue_o_55_;
  assign fe_queue_o_54_ = fetch_br_metadata_fwd_i[48];
  assign fe_queue_o[54] = fe_queue_o_54_;
  assign fe_queue_o_53_ = fetch_br_metadata_fwd_i[47];
  assign fe_queue_o[53] = fe_queue_o_53_;
  assign fe_queue_o_52_ = fetch_br_metadata_fwd_i[46];
  assign fe_queue_o[52] = fe_queue_o_52_;
  assign fe_queue_o_51_ = fetch_br_metadata_fwd_i[45];
  assign fe_queue_o[51] = fe_queue_o_51_;
  assign fe_queue_o_50_ = fetch_br_metadata_fwd_i[44];
  assign fe_queue_o[50] = fe_queue_o_50_;
  assign fe_queue_o_49_ = fetch_br_metadata_fwd_i[43];
  assign fe_queue_o[49] = fe_queue_o_49_;
  assign fe_queue_o_48_ = fetch_br_metadata_fwd_i[42];
  assign fe_queue_o[48] = fe_queue_o_48_;
  assign fe_queue_o_47_ = fetch_br_metadata_fwd_i[41];
  assign fe_queue_o[47] = fe_queue_o_47_;
  assign fe_queue_o_46_ = fetch_br_metadata_fwd_i[40];
  assign fe_queue_o[46] = fe_queue_o_46_;
  assign fe_queue_o_45_ = fetch_br_metadata_fwd_i[39];
  assign fe_queue_o[45] = fe_queue_o_45_;
  assign fe_queue_o_44_ = fetch_br_metadata_fwd_i[38];
  assign fe_queue_o[44] = fe_queue_o_44_;
  assign fe_queue_o_43_ = fetch_br_metadata_fwd_i[37];
  assign fe_queue_o[43] = fe_queue_o_43_;
  assign fe_queue_o_42_ = fetch_br_metadata_fwd_i[36];
  assign fe_queue_o[42] = fe_queue_o_42_;
  assign fe_queue_o_41_ = fetch_br_metadata_fwd_i[35];
  assign fe_queue_o[41] = fe_queue_o_41_;
  assign fe_queue_o_40_ = fetch_br_metadata_fwd_i[34];
  assign fe_queue_o[40] = fe_queue_o_40_;
  assign fe_queue_o_39_ = fetch_br_metadata_fwd_i[33];
  assign fe_queue_o[39] = fe_queue_o_39_;
  assign fe_queue_o_38_ = fetch_br_metadata_fwd_i[32];
  assign fe_queue_o[38] = fe_queue_o_38_;
  assign fe_queue_o_37_ = fetch_br_metadata_fwd_i[31];
  assign fe_queue_o[37] = fe_queue_o_37_;
  assign fe_queue_o_36_ = fetch_br_metadata_fwd_i[30];
  assign fe_queue_o[36] = fe_queue_o_36_;
  assign fe_queue_o_35_ = fetch_br_metadata_fwd_i[29];
  assign fe_queue_o[35] = fe_queue_o_35_;
  assign fe_queue_o_34_ = fetch_br_metadata_fwd_i[28];
  assign fe_queue_o[34] = fe_queue_o_34_;
  assign fe_queue_o_33_ = fetch_br_metadata_fwd_i[27];
  assign fe_queue_o[33] = fe_queue_o_33_;
  assign fe_queue_o_32_ = fetch_br_metadata_fwd_i[26];
  assign fe_queue_o[32] = fe_queue_o_32_;
  assign fe_queue_o_31_ = fetch_br_metadata_fwd_i[25];
  assign fe_queue_o[31] = fe_queue_o_31_;
  assign fe_queue_o_30_ = fetch_br_metadata_fwd_i[24];
  assign fe_queue_o[30] = fe_queue_o_30_;
  assign fe_queue_o_29_ = fetch_br_metadata_fwd_i[23];
  assign fe_queue_o[29] = fe_queue_o_29_;
  assign fe_queue_o_28_ = fetch_br_metadata_fwd_i[22];
  assign fe_queue_o[28] = fe_queue_o_28_;
  assign fe_queue_o_27_ = fetch_br_metadata_fwd_i[21];
  assign fe_queue_o[27] = fe_queue_o_27_;
  assign fe_queue_o_26_ = fetch_br_metadata_fwd_i[20];
  assign fe_queue_o[26] = fe_queue_o_26_;
  assign fe_queue_o_25_ = fetch_br_metadata_fwd_i[19];
  assign fe_queue_o[25] = fe_queue_o_25_;
  assign fe_queue_o_24_ = fetch_br_metadata_fwd_i[18];
  assign fe_queue_o[24] = fe_queue_o_24_;
  assign fe_queue_o_23_ = fetch_br_metadata_fwd_i[17];
  assign fe_queue_o[23] = fe_queue_o_23_;
  assign fe_queue_o_22_ = fetch_br_metadata_fwd_i[16];
  assign fe_queue_o[22] = fe_queue_o_22_;
  assign fe_queue_o_21_ = fetch_br_metadata_fwd_i[15];
  assign fe_queue_o[21] = fe_queue_o_21_;
  assign fe_queue_o_20_ = fetch_br_metadata_fwd_i[14];
  assign fe_queue_o[20] = fe_queue_o_20_;
  assign fe_queue_o_19_ = fetch_br_metadata_fwd_i[13];
  assign fe_queue_o[19] = fe_queue_o_19_;
  assign fe_queue_o_18_ = fetch_br_metadata_fwd_i[12];
  assign fe_queue_o[18] = fe_queue_o_18_;
  assign fe_queue_o_17_ = fetch_br_metadata_fwd_i[11];
  assign fe_queue_o[17] = fe_queue_o_17_;
  assign fe_queue_o_16_ = fetch_br_metadata_fwd_i[10];
  assign fe_queue_o[16] = fe_queue_o_16_;
  assign fe_queue_o_15_ = fetch_br_metadata_fwd_i[9];
  assign fe_queue_o[15] = fe_queue_o_15_;
  assign fe_queue_o_14_ = fetch_br_metadata_fwd_i[8];
  assign fe_queue_o[14] = fe_queue_o_14_;
  assign fe_queue_o_13_ = fetch_br_metadata_fwd_i[7];
  assign fe_queue_o[13] = fe_queue_o_13_;
  assign fe_queue_o_12_ = fetch_br_metadata_fwd_i[6];
  assign fe_queue_o[12] = fe_queue_o_12_;
  assign fe_queue_o_11_ = fetch_br_metadata_fwd_i[5];
  assign fe_queue_o[11] = fe_queue_o_11_;
  assign fe_queue_o_10_ = fetch_br_metadata_fwd_i[4];
  assign fe_queue_o[10] = fe_queue_o_10_;
  assign fe_queue_o_9_ = fetch_br_metadata_fwd_i[3];
  assign fe_queue_o[9] = fe_queue_o_9_;
  assign fe_queue_o_8_ = fetch_br_metadata_fwd_i[2];
  assign fe_queue_o[8] = fe_queue_o_8_;
  assign fe_queue_o_7_ = fetch_br_metadata_fwd_i[1];
  assign fe_queue_o[7] = fe_queue_o_7_;
  assign fe_queue_o_6_ = fetch_br_metadata_fwd_i[0];
  assign fe_queue_o[6] = fe_queue_o_6_;
  assign redirect_npc_o[38] = fe_cmd_i[113];
  assign itlb_w_vtag_o[26] = redirect_npc_o[38];
  assign attaboy_pc_o[38] = redirect_npc_o[38];
  assign redirect_npc_o[37] = fe_cmd_i[112];
  assign itlb_w_vtag_o[25] = redirect_npc_o[37];
  assign attaboy_pc_o[37] = redirect_npc_o[37];
  assign redirect_npc_o[36] = fe_cmd_i[111];
  assign itlb_w_vtag_o[24] = redirect_npc_o[36];
  assign attaboy_pc_o[36] = redirect_npc_o[36];
  assign redirect_npc_o[35] = fe_cmd_i[110];
  assign itlb_w_vtag_o[23] = redirect_npc_o[35];
  assign attaboy_pc_o[35] = redirect_npc_o[35];
  assign redirect_npc_o[34] = fe_cmd_i[109];
  assign itlb_w_vtag_o[22] = redirect_npc_o[34];
  assign attaboy_pc_o[34] = redirect_npc_o[34];
  assign redirect_npc_o[33] = fe_cmd_i[108];
  assign itlb_w_vtag_o[21] = redirect_npc_o[33];
  assign attaboy_pc_o[33] = redirect_npc_o[33];
  assign redirect_npc_o[32] = fe_cmd_i[107];
  assign itlb_w_vtag_o[20] = redirect_npc_o[32];
  assign attaboy_pc_o[32] = redirect_npc_o[32];
  assign redirect_npc_o[31] = fe_cmd_i[106];
  assign itlb_w_vtag_o[19] = redirect_npc_o[31];
  assign attaboy_pc_o[31] = redirect_npc_o[31];
  assign redirect_npc_o[30] = fe_cmd_i[105];
  assign itlb_w_vtag_o[18] = redirect_npc_o[30];
  assign attaboy_pc_o[30] = redirect_npc_o[30];
  assign redirect_npc_o[29] = fe_cmd_i[104];
  assign itlb_w_vtag_o[17] = redirect_npc_o[29];
  assign attaboy_pc_o[29] = redirect_npc_o[29];
  assign redirect_npc_o[28] = fe_cmd_i[103];
  assign itlb_w_vtag_o[16] = redirect_npc_o[28];
  assign attaboy_pc_o[28] = redirect_npc_o[28];
  assign redirect_npc_o[27] = fe_cmd_i[102];
  assign itlb_w_vtag_o[15] = redirect_npc_o[27];
  assign attaboy_pc_o[27] = redirect_npc_o[27];
  assign redirect_npc_o[26] = fe_cmd_i[101];
  assign itlb_w_vtag_o[14] = redirect_npc_o[26];
  assign attaboy_pc_o[26] = redirect_npc_o[26];
  assign redirect_npc_o[25] = fe_cmd_i[100];
  assign itlb_w_vtag_o[13] = redirect_npc_o[25];
  assign attaboy_pc_o[25] = redirect_npc_o[25];
  assign redirect_npc_o[24] = fe_cmd_i[99];
  assign itlb_w_vtag_o[12] = redirect_npc_o[24];
  assign attaboy_pc_o[24] = redirect_npc_o[24];
  assign redirect_npc_o[23] = fe_cmd_i[98];
  assign itlb_w_vtag_o[11] = redirect_npc_o[23];
  assign attaboy_pc_o[23] = redirect_npc_o[23];
  assign redirect_npc_o[22] = fe_cmd_i[97];
  assign itlb_w_vtag_o[10] = redirect_npc_o[22];
  assign attaboy_pc_o[22] = redirect_npc_o[22];
  assign redirect_npc_o[21] = fe_cmd_i[96];
  assign itlb_w_vtag_o[9] = redirect_npc_o[21];
  assign attaboy_pc_o[21] = redirect_npc_o[21];
  assign redirect_npc_o[20] = fe_cmd_i[95];
  assign itlb_w_vtag_o[8] = redirect_npc_o[20];
  assign attaboy_pc_o[20] = redirect_npc_o[20];
  assign redirect_npc_o[19] = fe_cmd_i[94];
  assign itlb_w_vtag_o[7] = redirect_npc_o[19];
  assign attaboy_pc_o[19] = redirect_npc_o[19];
  assign redirect_npc_o[18] = fe_cmd_i[93];
  assign itlb_w_vtag_o[6] = redirect_npc_o[18];
  assign attaboy_pc_o[18] = redirect_npc_o[18];
  assign redirect_npc_o[17] = fe_cmd_i[92];
  assign itlb_w_vtag_o[5] = redirect_npc_o[17];
  assign attaboy_pc_o[17] = redirect_npc_o[17];
  assign redirect_npc_o[16] = fe_cmd_i[91];
  assign itlb_w_vtag_o[4] = redirect_npc_o[16];
  assign attaboy_pc_o[16] = redirect_npc_o[16];
  assign redirect_npc_o[15] = fe_cmd_i[90];
  assign itlb_w_vtag_o[3] = redirect_npc_o[15];
  assign attaboy_pc_o[15] = redirect_npc_o[15];
  assign redirect_npc_o[14] = fe_cmd_i[89];
  assign itlb_w_vtag_o[2] = redirect_npc_o[14];
  assign attaboy_pc_o[14] = redirect_npc_o[14];
  assign redirect_npc_o[13] = fe_cmd_i[88];
  assign itlb_w_vtag_o[1] = redirect_npc_o[13];
  assign attaboy_pc_o[13] = redirect_npc_o[13];
  assign redirect_npc_o[12] = fe_cmd_i[87];
  assign itlb_w_vtag_o[0] = redirect_npc_o[12];
  assign attaboy_pc_o[12] = redirect_npc_o[12];
  assign redirect_npc_o[11] = fe_cmd_i[86];
  assign attaboy_pc_o[11] = redirect_npc_o[11];
  assign redirect_npc_o[10] = fe_cmd_i[85];
  assign attaboy_pc_o[10] = redirect_npc_o[10];
  assign redirect_npc_o[9] = fe_cmd_i[84];
  assign attaboy_pc_o[9] = redirect_npc_o[9];
  assign redirect_npc_o[8] = fe_cmd_i[83];
  assign attaboy_pc_o[8] = redirect_npc_o[8];
  assign redirect_npc_o[7] = fe_cmd_i[82];
  assign attaboy_pc_o[7] = redirect_npc_o[7];
  assign redirect_npc_o[6] = fe_cmd_i[81];
  assign attaboy_pc_o[6] = redirect_npc_o[6];
  assign redirect_npc_o[5] = fe_cmd_i[80];
  assign attaboy_pc_o[5] = redirect_npc_o[5];
  assign redirect_npc_o[4] = fe_cmd_i[79];
  assign attaboy_pc_o[4] = redirect_npc_o[4];
  assign redirect_npc_o[3] = fe_cmd_i[78];
  assign attaboy_pc_o[3] = redirect_npc_o[3];
  assign redirect_npc_o[2] = fe_cmd_i[77];
  assign attaboy_pc_o[2] = redirect_npc_o[2];
  assign redirect_npc_o[1] = fe_cmd_i[76];
  assign attaboy_pc_o[1] = redirect_npc_o[1];
  assign redirect_npc_o[0] = fe_cmd_i[75];
  assign attaboy_pc_o[0] = redirect_npc_o[0];
  assign redirect_br_metadata_fwd_o[48] = fe_cmd_i[68];
  assign itlb_w_entry_o[32] = redirect_br_metadata_fwd_o[48];
  assign attaboy_br_metadata_fwd_o[46] = redirect_br_metadata_fwd_o[48];
  assign redirect_br_metadata_fwd_o[47] = fe_cmd_i[67];
  assign itlb_w_entry_o[31] = redirect_br_metadata_fwd_o[47];
  assign attaboy_br_metadata_fwd_o[45] = redirect_br_metadata_fwd_o[47];
  assign redirect_br_metadata_fwd_o[46] = fe_cmd_i[66];
  assign itlb_w_entry_o[30] = redirect_br_metadata_fwd_o[46];
  assign attaboy_br_metadata_fwd_o[44] = redirect_br_metadata_fwd_o[46];
  assign redirect_br_metadata_fwd_o[45] = fe_cmd_i[65];
  assign itlb_w_entry_o[29] = redirect_br_metadata_fwd_o[45];
  assign attaboy_br_metadata_fwd_o[43] = redirect_br_metadata_fwd_o[45];
  assign redirect_br_metadata_fwd_o[44] = fe_cmd_i[64];
  assign itlb_w_entry_o[28] = redirect_br_metadata_fwd_o[44];
  assign attaboy_br_metadata_fwd_o[42] = redirect_br_metadata_fwd_o[44];
  assign redirect_br_metadata_fwd_o[43] = fe_cmd_i[63];
  assign itlb_w_entry_o[27] = redirect_br_metadata_fwd_o[43];
  assign attaboy_br_metadata_fwd_o[41] = redirect_br_metadata_fwd_o[43];
  assign redirect_br_metadata_fwd_o[42] = fe_cmd_i[62];
  assign itlb_w_entry_o[26] = redirect_br_metadata_fwd_o[42];
  assign attaboy_br_metadata_fwd_o[40] = redirect_br_metadata_fwd_o[42];
  assign redirect_br_metadata_fwd_o[41] = fe_cmd_i[61];
  assign itlb_w_entry_o[25] = redirect_br_metadata_fwd_o[41];
  assign attaboy_br_metadata_fwd_o[39] = redirect_br_metadata_fwd_o[41];
  assign redirect_br_metadata_fwd_o[40] = fe_cmd_i[60];
  assign itlb_w_entry_o[24] = redirect_br_metadata_fwd_o[40];
  assign attaboy_br_metadata_fwd_o[38] = redirect_br_metadata_fwd_o[40];
  assign redirect_br_metadata_fwd_o[39] = fe_cmd_i[59];
  assign itlb_w_entry_o[23] = redirect_br_metadata_fwd_o[39];
  assign attaboy_br_metadata_fwd_o[37] = redirect_br_metadata_fwd_o[39];
  assign redirect_br_metadata_fwd_o[38] = fe_cmd_i[58];
  assign itlb_w_entry_o[22] = redirect_br_metadata_fwd_o[38];
  assign attaboy_br_metadata_fwd_o[36] = redirect_br_metadata_fwd_o[38];
  assign redirect_br_metadata_fwd_o[37] = fe_cmd_i[57];
  assign itlb_w_entry_o[21] = redirect_br_metadata_fwd_o[37];
  assign attaboy_br_metadata_fwd_o[35] = redirect_br_metadata_fwd_o[37];
  assign redirect_br_metadata_fwd_o[36] = fe_cmd_i[56];
  assign itlb_w_entry_o[20] = redirect_br_metadata_fwd_o[36];
  assign attaboy_br_metadata_fwd_o[34] = redirect_br_metadata_fwd_o[36];
  assign redirect_br_metadata_fwd_o[35] = fe_cmd_i[55];
  assign itlb_w_entry_o[19] = redirect_br_metadata_fwd_o[35];
  assign attaboy_br_metadata_fwd_o[33] = redirect_br_metadata_fwd_o[35];
  assign redirect_br_metadata_fwd_o[34] = fe_cmd_i[54];
  assign itlb_w_entry_o[18] = redirect_br_metadata_fwd_o[34];
  assign attaboy_br_metadata_fwd_o[32] = redirect_br_metadata_fwd_o[34];
  assign redirect_br_metadata_fwd_o[33] = fe_cmd_i[53];
  assign itlb_w_entry_o[17] = redirect_br_metadata_fwd_o[33];
  assign attaboy_br_metadata_fwd_o[31] = redirect_br_metadata_fwd_o[33];
  assign redirect_br_metadata_fwd_o[32] = fe_cmd_i[52];
  assign itlb_w_entry_o[16] = redirect_br_metadata_fwd_o[32];
  assign attaboy_br_metadata_fwd_o[30] = redirect_br_metadata_fwd_o[32];
  assign redirect_br_metadata_fwd_o[31] = fe_cmd_i[51];
  assign itlb_w_entry_o[15] = redirect_br_metadata_fwd_o[31];
  assign attaboy_br_metadata_fwd_o[29] = redirect_br_metadata_fwd_o[31];
  assign redirect_br_metadata_fwd_o[30] = fe_cmd_i[50];
  assign itlb_w_entry_o[14] = redirect_br_metadata_fwd_o[30];
  assign attaboy_br_metadata_fwd_o[28] = redirect_br_metadata_fwd_o[30];
  assign redirect_br_metadata_fwd_o[29] = fe_cmd_i[49];
  assign itlb_w_entry_o[13] = redirect_br_metadata_fwd_o[29];
  assign attaboy_br_metadata_fwd_o[27] = redirect_br_metadata_fwd_o[29];
  assign redirect_br_metadata_fwd_o[28] = fe_cmd_i[48];
  assign itlb_w_entry_o[12] = redirect_br_metadata_fwd_o[28];
  assign attaboy_br_metadata_fwd_o[26] = redirect_br_metadata_fwd_o[28];
  assign redirect_br_metadata_fwd_o[27] = fe_cmd_i[47];
  assign itlb_w_entry_o[11] = redirect_br_metadata_fwd_o[27];
  assign attaboy_br_metadata_fwd_o[25] = redirect_br_metadata_fwd_o[27];
  assign redirect_br_metadata_fwd_o[26] = fe_cmd_i[46];
  assign itlb_w_entry_o[10] = redirect_br_metadata_fwd_o[26];
  assign attaboy_br_metadata_fwd_o[24] = redirect_br_metadata_fwd_o[26];
  assign redirect_br_metadata_fwd_o[25] = fe_cmd_i[45];
  assign itlb_w_entry_o[9] = redirect_br_metadata_fwd_o[25];
  assign attaboy_br_metadata_fwd_o[23] = redirect_br_metadata_fwd_o[25];
  assign redirect_br_metadata_fwd_o[24] = fe_cmd_i[44];
  assign itlb_w_entry_o[8] = redirect_br_metadata_fwd_o[24];
  assign attaboy_br_metadata_fwd_o[22] = redirect_br_metadata_fwd_o[24];
  assign redirect_br_metadata_fwd_o[23] = fe_cmd_i[43];
  assign itlb_w_entry_o[7] = redirect_br_metadata_fwd_o[23];
  assign attaboy_br_metadata_fwd_o[21] = redirect_br_metadata_fwd_o[23];
  assign redirect_br_metadata_fwd_o[22] = fe_cmd_i[42];
  assign itlb_w_entry_o[6] = redirect_br_metadata_fwd_o[22];
  assign attaboy_br_metadata_fwd_o[20] = redirect_br_metadata_fwd_o[22];
  assign redirect_br_metadata_fwd_o[21] = fe_cmd_i[41];
  assign itlb_w_entry_o[5] = redirect_br_metadata_fwd_o[21];
  assign attaboy_br_metadata_fwd_o[19] = redirect_br_metadata_fwd_o[21];
  assign redirect_br_metadata_fwd_o[20] = fe_cmd_i[40];
  assign itlb_w_entry_o[4] = redirect_br_metadata_fwd_o[20];
  assign attaboy_br_metadata_fwd_o[18] = redirect_br_metadata_fwd_o[20];
  assign redirect_br_metadata_fwd_o[19] = fe_cmd_i[39];
  assign itlb_w_entry_o[3] = redirect_br_metadata_fwd_o[19];
  assign attaboy_br_metadata_fwd_o[17] = redirect_br_metadata_fwd_o[19];
  assign redirect_br_metadata_fwd_o[18] = fe_cmd_i[38];
  assign itlb_w_entry_o[2] = redirect_br_metadata_fwd_o[18];
  assign attaboy_br_metadata_fwd_o[16] = redirect_br_metadata_fwd_o[18];
  assign redirect_br_metadata_fwd_o[17] = fe_cmd_i[37];
  assign itlb_w_entry_o[1] = redirect_br_metadata_fwd_o[17];
  assign attaboy_br_metadata_fwd_o[15] = redirect_br_metadata_fwd_o[17];
  assign redirect_br_metadata_fwd_o[16] = fe_cmd_i[36];
  assign itlb_w_entry_o[0] = redirect_br_metadata_fwd_o[16];
  assign attaboy_br_metadata_fwd_o[14] = redirect_br_metadata_fwd_o[16];
  assign redirect_br_metadata_fwd_o[15] = fe_cmd_i[35];
  assign attaboy_br_metadata_fwd_o[13] = redirect_br_metadata_fwd_o[15];
  assign redirect_br_metadata_fwd_o[14] = fe_cmd_i[34];
  assign attaboy_br_metadata_fwd_o[12] = redirect_br_metadata_fwd_o[14];
  assign redirect_br_metadata_fwd_o[13] = fe_cmd_i[33];
  assign attaboy_br_metadata_fwd_o[11] = redirect_br_metadata_fwd_o[13];
  assign redirect_br_metadata_fwd_o[12] = fe_cmd_i[32];
  assign attaboy_br_metadata_fwd_o[10] = redirect_br_metadata_fwd_o[12];
  assign redirect_br_metadata_fwd_o[11] = fe_cmd_i[31];
  assign attaboy_br_metadata_fwd_o[9] = redirect_br_metadata_fwd_o[11];
  assign redirect_br_metadata_fwd_o[10] = fe_cmd_i[30];
  assign attaboy_br_metadata_fwd_o[8] = redirect_br_metadata_fwd_o[10];
  assign redirect_br_metadata_fwd_o[9] = fe_cmd_i[29];
  assign attaboy_br_metadata_fwd_o[7] = redirect_br_metadata_fwd_o[9];
  assign redirect_br_metadata_fwd_o[8] = fe_cmd_i[28];
  assign attaboy_br_metadata_fwd_o[6] = redirect_br_metadata_fwd_o[8];
  assign redirect_br_metadata_fwd_o[7] = fe_cmd_i[27];
  assign attaboy_br_metadata_fwd_o[5] = redirect_br_metadata_fwd_o[7];
  assign redirect_br_metadata_fwd_o[6] = fe_cmd_i[26];
  assign attaboy_br_metadata_fwd_o[4] = redirect_br_metadata_fwd_o[6];
  assign redirect_br_metadata_fwd_o[5] = fe_cmd_i[25];
  assign attaboy_br_metadata_fwd_o[3] = redirect_br_metadata_fwd_o[5];
  assign redirect_br_metadata_fwd_o[4] = fe_cmd_i[24];
  assign attaboy_br_metadata_fwd_o[2] = redirect_br_metadata_fwd_o[4];
  assign redirect_br_metadata_fwd_o[3] = fe_cmd_i[23];
  assign attaboy_br_metadata_fwd_o[1] = redirect_br_metadata_fwd_o[3];
  assign redirect_br_metadata_fwd_o[2] = fe_cmd_i[22];
  assign attaboy_br_metadata_fwd_o[0] = redirect_br_metadata_fwd_o[2];
  assign redirect_br_metadata_fwd_o[1] = fe_cmd_i[21];
  assign redirect_br_metadata_fwd_o[0] = fe_cmd_i[20];
  assign attaboy_br_metadata_fwd_o_48_ = fe_cmd_i[70];
  assign itlb_w_entry_o[34] = attaboy_br_metadata_fwd_o_48_;
  assign attaboy_br_metadata_fwd_o[48] = attaboy_br_metadata_fwd_o_48_;
  assign attaboy_br_metadata_fwd_o_47_ = fe_cmd_i[69];
  assign itlb_w_entry_o[33] = attaboy_br_metadata_fwd_o_47_;
  assign attaboy_br_metadata_fwd_o[47] = attaboy_br_metadata_fwd_o_47_;
  assign itlb_w_entry_o_35_ = fe_cmd_i[71];
  assign itlb_w_entry_o[35] = itlb_w_entry_o_35_;
  assign icache_pkt_o_71_ = next_pc_i[38];
  assign icache_pkt_o[71] = icache_pkt_o_71_;
  assign icache_pkt_o_70_ = next_pc_i[37];
  assign icache_pkt_o[70] = icache_pkt_o_70_;
  assign icache_pkt_o_69_ = next_pc_i[36];
  assign icache_pkt_o[69] = icache_pkt_o_69_;
  assign icache_pkt_o_68_ = next_pc_i[35];
  assign icache_pkt_o[68] = icache_pkt_o_68_;
  assign icache_pkt_o_67_ = next_pc_i[34];
  assign icache_pkt_o[67] = icache_pkt_o_67_;
  assign icache_pkt_o_66_ = next_pc_i[33];
  assign icache_pkt_o[66] = icache_pkt_o_66_;
  assign icache_pkt_o_65_ = next_pc_i[32];
  assign icache_pkt_o[65] = icache_pkt_o_65_;
  assign icache_pkt_o_64_ = next_pc_i[31];
  assign icache_pkt_o[64] = icache_pkt_o_64_;
  assign icache_pkt_o_63_ = next_pc_i[30];
  assign icache_pkt_o[63] = icache_pkt_o_63_;
  assign icache_pkt_o_62_ = next_pc_i[29];
  assign icache_pkt_o[62] = icache_pkt_o_62_;
  assign icache_pkt_o_61_ = next_pc_i[28];
  assign icache_pkt_o[61] = icache_pkt_o_61_;
  assign icache_pkt_o_60_ = next_pc_i[27];
  assign icache_pkt_o[60] = icache_pkt_o_60_;
  assign icache_pkt_o_59_ = next_pc_i[26];
  assign icache_pkt_o[59] = icache_pkt_o_59_;
  assign icache_pkt_o_58_ = next_pc_i[25];
  assign icache_pkt_o[58] = icache_pkt_o_58_;
  assign icache_pkt_o_57_ = next_pc_i[24];
  assign icache_pkt_o[57] = icache_pkt_o_57_;
  assign icache_pkt_o_56_ = next_pc_i[23];
  assign icache_pkt_o[56] = icache_pkt_o_56_;
  assign icache_pkt_o_55_ = next_pc_i[22];
  assign icache_pkt_o[55] = icache_pkt_o_55_;
  assign icache_pkt_o_54_ = next_pc_i[21];
  assign icache_pkt_o[54] = icache_pkt_o_54_;
  assign icache_pkt_o_53_ = next_pc_i[20];
  assign icache_pkt_o[53] = icache_pkt_o_53_;
  assign icache_pkt_o_52_ = next_pc_i[19];
  assign icache_pkt_o[52] = icache_pkt_o_52_;
  assign icache_pkt_o_51_ = next_pc_i[18];
  assign icache_pkt_o[51] = icache_pkt_o_51_;
  assign icache_pkt_o_50_ = next_pc_i[17];
  assign icache_pkt_o[50] = icache_pkt_o_50_;
  assign icache_pkt_o_49_ = next_pc_i[16];
  assign icache_pkt_o[49] = icache_pkt_o_49_;
  assign icache_pkt_o_48_ = next_pc_i[15];
  assign icache_pkt_o[48] = icache_pkt_o_48_;
  assign icache_pkt_o_47_ = next_pc_i[14];
  assign icache_pkt_o[47] = icache_pkt_o_47_;
  assign icache_pkt_o_46_ = next_pc_i[13];
  assign icache_pkt_o[46] = icache_pkt_o_46_;
  assign icache_pkt_o_45_ = next_pc_i[12];
  assign icache_pkt_o[45] = icache_pkt_o_45_;
  assign icache_pkt_o_44_ = next_pc_i[11];
  assign icache_pkt_o[44] = icache_pkt_o_44_;
  assign icache_pkt_o_43_ = next_pc_i[10];
  assign icache_pkt_o[43] = icache_pkt_o_43_;
  assign icache_pkt_o_42_ = next_pc_i[9];
  assign icache_pkt_o[42] = icache_pkt_o_42_;
  assign icache_pkt_o_41_ = next_pc_i[8];
  assign icache_pkt_o[41] = icache_pkt_o_41_;
  assign icache_pkt_o_40_ = next_pc_i[7];
  assign icache_pkt_o[40] = icache_pkt_o_40_;
  assign icache_pkt_o_39_ = next_pc_i[6];
  assign icache_pkt_o[39] = icache_pkt_o_39_;
  assign icache_pkt_o_38_ = next_pc_i[5];
  assign icache_pkt_o[38] = icache_pkt_o_38_;
  assign icache_pkt_o_37_ = next_pc_i[4];
  assign icache_pkt_o[37] = icache_pkt_o_37_;
  assign icache_pkt_o_36_ = next_pc_i[3];
  assign icache_pkt_o[36] = icache_pkt_o_36_;
  assign icache_pkt_o_35_ = next_pc_i[2];
  assign icache_pkt_o[35] = icache_pkt_o_35_;
  assign icache_pkt_o_34_ = next_pc_i[1];
  assign icache_pkt_o[34] = icache_pkt_o_34_;
  assign icache_pkt_o_33_ = next_pc_i[0];
  assign icache_pkt_o[33] = icache_pkt_o_33_;
  assign shadow_priv_o[1] = fe_cmd_i[16];
  assign shadow_priv_o[0] = fe_cmd_i[15];
  assign N15 = fe_cmd_i[3:1] > 1'b0;
  assign N17 = redirect_br_metadata_fwd_o[19:17] > 1'b0;

  bsg_dff_reset_en_width_p3
  exception_reg
  (
    .clk_i(clk_i),
    .reset_i(_0_net_),
    .en_i(tv_we_i),
    .data_i({ itlb_miss_tl_i, instr_page_fault_tl_i, instr_access_fault_tl_i }),
    .data_o({ itlb_miss_tv_r, instr_page_fault_tv_r, instr_access_fault_tv_r })
  );

  assign N20 = fetch_count_i > 1'b0;
  assign N33 = N103 & N71;
  assign N34 = state_r[1] | N71;
  assign N36 = state_r[1] & state_r[0];
  assign N37 = N103 | state_r[0];
  assign N71 = ~state_r[0];
  assign N72 = N71 | state_r[1];
  assign N73 = ~fe_cmd_i[18];
  assign N74 = N73 | fe_cmd_i[19];
  assign N75 = ~N74;
  assign N76 = ~fe_cmd_i[19];
  assign N77 = fe_cmd_i[18] | N76;
  assign N78 = ~N77;
  assign N79 = fe_cmd_i[18] | fe_cmd_i[19];
  assign N80 = ~N79;
  assign N81 = ~attaboy_br_metadata_fwd_o_48_;
  assign N82 = N81 | itlb_w_entry_o_35_;
  assign N83 = attaboy_br_metadata_fwd_o_47_ | N82;
  assign N84 = ~N83;
  assign N85 = ~attaboy_br_metadata_fwd_o_47_;
  assign N86 = N81 | itlb_w_entry_o_35_;
  assign N87 = N85 | N86;
  assign N88 = ~N87;
  assign N89 = attaboy_br_metadata_fwd_o_48_ | itlb_w_entry_o_35_;
  assign N90 = N85 | N89;
  assign N91 = ~N90;
  assign N92 = attaboy_br_metadata_fwd_o_48_ | itlb_w_entry_o_35_;
  assign N93 = attaboy_br_metadata_fwd_o_47_ | N92;
  assign N94 = ~N93;
  assign N95 = ~itlb_w_entry_o_35_;
  assign N96 = attaboy_br_metadata_fwd_o_48_ | N95;
  assign N97 = N85 | N96;
  assign N98 = ~N97;
  assign N99 = ~fe_cmd_i[73];
  assign N100 = N99 | fe_cmd_i[74];
  assign N101 = fe_cmd_i[72] | N100;
  assign N102 = ~N101;
  assign N103 = ~state_r[1];
  assign N104 = state_r[0] | N103;
  assign N105 = ~N104;
  assign N106 = ~fe_cmd_i[74];
  assign N107 = fe_cmd_i[73] | N106;
  assign N108 = fe_cmd_i[72] | N107;
  assign N109 = ~N108;
  assign N110 = N99 | N106;
  assign N111 = fe_cmd_i[72] | N110;
  assign N112 = ~N111;
  assign N113 = ~fe_cmd_i[72];
  assign N114 = fe_cmd_i[73] | fe_cmd_i[74];
  assign N115 = N113 | N114;
  assign N116 = ~N115;
  assign N117 = N113 | N100;
  assign N118 = ~N117;
  assign N119 = fe_cmd_i[73] & fe_cmd_i[74];
  assign N120 = fe_cmd_i[72] & N119;
  assign N121 = N113 | N107;
  assign N122 = ~N121;
  assign N123 = fe_cmd_i[72] | N114;
  assign N124 = ~N123;
  assign redirect_pc_o = redirect_npc_o - { redirect_resume_o, 1'b0 };
  assign redirect_instr_o = (N0)? { fe_cmd_i[19:18], fe_cmd_i_17_, shadow_priv_o, fe_cmd_i[14:4] } : 
                            (N1)? redirect_br_metadata_fwd_o[35:20] : 1'b0;
  assign N0 = itlb_fill_response_v;
  assign N1 = N12;
  assign redirect_resume_o = (N0)? N15 : 
                             (N19)? N17 : 
                             (N14)? 1'b0 : 1'b0;
  assign fe_queue_o[2:0] = (N2)? { 1'b1, 1'b0, 1'b0 } : 
                           (N26)? { 1'b0, 1'b0, 1'b0 } : 
                           (N29)? { 1'b0, 1'b0, 1'b1 } : 
                           (N32)? { 1'b0, 1'b1, 1'b0 } : 
                           (N24)? { 1'b0, 1'b1, 1'b1 } : 1'b0;
  assign N2 = fetch_instr_v;
  assign fe_queue_o[5:3] = (N2)? fetch_count_i : 
                           (N3)? { 1'b0, 1'b0, fetch_partial_i } : 1'b0;
  assign N3 = N141;
  assign { N51, N50 } = (N4)? { 1'b0, 1'b1 } : 
                        (N5)? state_r : 1'b0;
  assign N4 = fetch_exception_v;
  assign N5 = N49;
  assign N52 = (N6)? 1'b1 : 
               (N62)? icache_fence_v : 
               (N46)? 1'b1 : 1'b0;
  assign N6 = cmd_immediate_v;
  assign N53 = (N6)? 1'b1 : 
               (N62)? 1'b1 : 
               (N46)? ovr_i : 1'b0;
  assign N54 = (N6)? icache_yumi_i : 
               (N62)? 1'b0 : 
               (N46)? icache_yumi_i : 1'b0;
  assign N55 = (N6)? icache_yumi_i : 
               (N62)? 1'b0 : 
               (N46)? N48 : 1'b0;
  assign N56 = (N6)? 1'b0 : 
               (N62)? itlb_fill_response_v : 
               (N46)? 1'b0 : 1'b0;
  assign N57 = (N6)? 1'b0 : 
               (N62)? itlb_fence_v : 
               (N46)? 1'b0 : 1'b0;
  assign N58 = (N6)? 1'b0 : 
               (N62)? N47 : 
               (N46)? 1'b0 : 1'b0;
  assign { N60, N59 } = (N62)? { 1'b1, 1'b1 } : 
                        (N46)? { N51, N50 } : 1'b0;
  assign fe_cmd_yumi_o = (N7)? N39 : 
                         (N8)? N42 : 
                         (N9)? icache_yumi_i : 
                         (N10)? N55 : 1'b0;
  assign N7 = N33;
  assign N8 = N35;
  assign N9 = N36;
  assign N10 = N38;
  assign state_n = (N7)? { 1'b1, 1'b1 } : 
                   (N8)? { 1'b1, 1'b0 } : 
                   (N9)? { 1'b1, 1'b0 } : 
                   (N10)? { N60, N59 } : 1'b0;
  assign tl_flush_o = (N7)? 1'b0 : 
                      (N8)? 1'b1 : 
                      (N9)? 1'b0 : 
                      (N10)? N58 : 1'b0;
  assign tv_flush_o = (N7)? 1'b0 : 
                      (N8)? 1'b1 : 
                      (N9)? 1'b0 : 
                      (N10)? N53 : 1'b0;
  assign icache_v_o = (N7)? 1'b0 : 
                      (N8)? 1'b0 : 
                      (N9)? fe_cmd_v_i : 
                      (N10)? N52 : 1'b0;
  assign itlb_r_v_o = (N7)? 1'b0 : 
                      (N8)? 1'b0 : 
                      (N9)? icache_yumi_i : 
                      (N10)? N54 : 1'b0;
  assign icache_force_o = (N7)? 1'b0 : 
                          (N8)? 1'b0 : 
                          (N9)? 1'b0 : 
                          (N10)? N53 : 1'b0;
  assign itlb_w_v_o = (N7)? 1'b0 : 
                      (N8)? 1'b0 : 
                      (N9)? 1'b0 : 
                      (N10)? N56 : 1'b0;
  assign itlb_fence_v_o = (N7)? 1'b0 : 
                          (N8)? 1'b0 : 
                          (N9)? 1'b0 : 
                          (N10)? N57 : 1'b0;
  assign pc_redirect_v = fe_cmd_v_i & N116;
  assign icache_fill_response_v = fe_cmd_v_i & N118;
  assign icache_fence_v = fe_cmd_v_i & N109;
  assign state_reset_v = fe_cmd_v_i & N124;
  assign itlb_fill_response_v = fe_cmd_v_i & N122;
  assign itlb_fence_v = fe_cmd_v_i & N112;
  assign wait_v = fe_cmd_v_i & N120;
  assign br_miss_v = pc_redirect_v & N84;
  assign eret_v = pc_redirect_v & N94;
  assign interrupt_v = pc_redirect_v & N91;
  assign trap_v = pc_redirect_v & N88;
  assign translation_v = pc_redirect_v & N98;
  assign redirect_br_taken_o = br_miss_v & N75;
  assign redirect_br_ntaken_o = br_miss_v & N78;
  assign redirect_br_nonbr_o = br_miss_v & N80;
  assign attaboy_v_o = fe_cmd_v_i & N102;
  assign cmd_nonattaboy_v = fe_cmd_v_i & N101;
  assign cmd_immediate_v = fe_cmd_v_i & N126;
  assign N126 = N125 | wait_v;
  assign N125 = pc_redirect_v | icache_fill_response_v;
  assign cmd_complex_v = fe_cmd_v_i & N129;
  assign N129 = N128 | itlb_fence_v;
  assign N128 = N127 | icache_fence_v;
  assign N127 = state_reset_v | itlb_fill_response_v;
  assign redirect_v_o = N72 & cmd_nonattaboy_v;
  assign redirect_br_v_o = N72 & br_miss_v;
  assign attaboy_force_o = ~fe_queue_ready_and_i;
  assign attaboy_taken_o = attaboy_v_o & itlb_w_entry_o_35_;
  assign attaboy_ntaken_o = attaboy_v_o & N95;
  assign shadow_priv_w_o = N131 | eret_v;
  assign N131 = N130 | interrupt_v;
  assign N130 = state_reset_v | trap_v;
  assign shadow_translation_en_w_o = N134 | translation_v;
  assign N134 = N133 | eret_v;
  assign N133 = N132 | interrupt_v;
  assign N132 = state_reset_v | trap_v;
  assign N11 = N105 & icache_fence_v;
  assign icache_pkt_o[1] = N11;
  assign icache_pkt_o[0] = ~icache_fill_response_v;
  assign N12 = ~itlb_fill_response_v;
  assign N13 = icache_fill_response_v | itlb_fill_response_v;
  assign N14 = ~N13;
  assign N16 = N19;
  assign N18 = ~itlb_fill_response_v;
  assign N19 = icache_fill_response_v & N18;
  assign _0_net_ = reset_i | tv_flush_o;
  assign if2_exception_v = N136 | icache_miss_tv_i;
  assign N136 = N135 | instr_access_fault_tv_r;
  assign N135 = itlb_miss_tv_r | instr_page_fault_tv_r;
  assign fetch_instr_v = N138 & N20;
  assign N138 = N137 & fetch_v_i;
  assign N137 = N105 & fe_queue_ready_and_i;
  assign fetch_exception_v = N140 & N141;
  assign N140 = N139 & if2_exception_v;
  assign N139 = N105 & fe_queue_ready_and_i;
  assign N141 = ~fetch_instr_v;
  assign fetch_yumi_o = N142 & fetch_v_i;
  assign N142 = N105 & fe_queue_ready_and_i;
  assign fe_queue_v_o = fetch_instr_v | fetch_exception_v;
  assign N21 = itlb_miss_tv_r | fetch_instr_v;
  assign N22 = instr_page_fault_tv_r | N21;
  assign N23 = instr_access_fault_tv_r | N22;
  assign N24 = ~N23;
  assign N25 = ~fetch_instr_v;
  assign N26 = itlb_miss_tv_r & N25;
  assign N27 = ~itlb_miss_tv_r;
  assign N28 = N25 & N27;
  assign N29 = instr_page_fault_tv_r & N28;
  assign N30 = ~instr_page_fault_tv_r;
  assign N31 = N28 & N30;
  assign N32 = instr_access_fault_tv_r & N31;
  assign N35 = ~N34;
  assign N38 = ~N37;
  assign N39 = fe_cmd_v_i & N143;
  assign N143 = ~state_reset_v;
  assign N40 = state_reset_v & pc_gen_init_done_i;
  assign N41 = ~N40;
  assign N42 = attaboy_v_o & attaboy_yumi_i;
  assign N43 = ~cmd_nonattaboy_v;
  assign N44 = ~icache_yumi_i;
  assign N45 = cmd_complex_v | cmd_immediate_v;
  assign N46 = ~N45;
  assign N47 = itlb_fill_response_v | itlb_fence_v;
  assign N48 = attaboy_v_o & attaboy_yumi_i;
  assign N49 = ~fetch_exception_v;
  assign N61 = ~cmd_immediate_v;
  assign N62 = cmd_complex_v & N61;
  assign N63 = N41 & N33;
  assign N64 = N43 & N35;
  assign N65 = N63 | N64;
  assign N66 = N44 & N36;
  assign N67 = N65 | N66;
  assign N68 = cmd_immediate_v & N38;
  assign N69 = N67 | N68;
  assign N70 = ~N69;

  always @(posedge clk_i) begin
    if(reset_i) begin
      state_r_1_sv2v_reg <= 1'b0;
      state_r_0_sv2v_reg <= 1'b0;
    end else if(N70) begin
      state_r_1_sv2v_reg <= state_n[1];
      state_r_0_sv2v_reg <= state_n[0];
    end 
  end


endmodule



module bp_fe_top
(
  clk_i,
  reset_i,
  cfg_bus_i,
  fe_cmd_i,
  fe_cmd_v_i,
  fe_cmd_yumi_o,
  fe_queue_o,
  fe_queue_v_o,
  fe_queue_ready_and_i,
  cache_req_o,
  cache_req_v_o,
  cache_req_yumi_i,
  cache_req_lock_i,
  cache_req_metadata_o,
  cache_req_metadata_v_o,
  cache_req_id_i,
  cache_req_critical_i,
  cache_req_last_i,
  cache_req_credits_full_i,
  cache_req_credits_empty_i,
  data_mem_pkt_i,
  data_mem_pkt_v_i,
  data_mem_pkt_yumi_o,
  data_mem_o,
  tag_mem_pkt_i,
  tag_mem_pkt_v_i,
  tag_mem_pkt_yumi_o,
  tag_mem_o,
  stat_mem_pkt_i,
  stat_mem_pkt_v_i,
  stat_mem_pkt_yumi_o,
  stat_mem_o
);

  input [60:0] cfg_bus_i;
  input [113:0] fe_cmd_i;
  output [173:0] fe_queue_o;
  output [116:0] cache_req_o;
  output [3:0] cache_req_metadata_o;
  input [0:0] cache_req_id_i;
  input [142:0] data_mem_pkt_i;
  output [511:0] data_mem_o;
  input [34:0] tag_mem_pkt_i;
  output [22:0] tag_mem_o;
  input [10:0] stat_mem_pkt_i;
  output [14:0] stat_mem_o;
  input clk_i;
  input reset_i;
  input fe_cmd_v_i;
  input fe_queue_ready_and_i;
  input cache_req_yumi_i;
  input cache_req_lock_i;
  input cache_req_critical_i;
  input cache_req_last_i;
  input cache_req_credits_full_i;
  input cache_req_credits_empty_i;
  input data_mem_pkt_v_i;
  input tag_mem_pkt_v_i;
  input stat_mem_pkt_v_i;
  output fe_cmd_yumi_o;
  output fe_queue_v_o;
  output cache_req_v_o;
  output cache_req_metadata_v_o;
  output data_mem_pkt_yumi_o;
  output tag_mem_pkt_yumi_o;
  output stat_mem_pkt_yumi_o;
  wire [173:0] fe_queue_o;
  wire [116:0] cache_req_o;
  wire [3:0] cache_req_metadata_o;
  wire [511:0] data_mem_o;
  wire [22:0] tag_mem_o;
  wire [14:0] stat_mem_o;
  wire fe_cmd_yumi_o,fe_queue_v_o,cache_req_v_o,cache_req_metadata_v_o,
  data_mem_pkt_yumi_o,tag_mem_pkt_yumi_o,stat_mem_pkt_yumi_o,shadow_priv_w,
  shadow_translation_en_w,shadow_translation_en_n,shadow_translation_en_r,pc_gen_init_done_lo,
  attaboy_v_li,attaboy_force_li,attaboy_taken_li,attaboy_ntaken_li,attaboy_yumi_lo,
  redirect_v_li,redirect_br_v_li,redirect_br_taken_li,redirect_br_ntaken_li,
  redirect_br_nonbr_li,icache_yumi_lo,ovr_lo,icache_tv_we,icache_hit_v_lo,icache_miss_v_lo,
  icache_hit_yumi_li,if2_hit_v_lo,if2_miss_v_lo,if2_yumi_li,fetch_startup_lo,
  fetch_catchup_lo,fetch_rebase_lo,fetch_linear_lo,fetch_yumi_li,fetch_taken_li,tv_flush_lo,
  itlb_fence_v_li,itlb_w_v_li,itlb_r_v_li,ptag_v_lo,ptag_miss_lo,ptag_uncached_lo,
  ptag_nonidem_lo,ptag_dram_lo,instr_access_fault_lo,instr_page_fault_lo,
  icache_v_li,icache_force_li,tl_flush_lo,icache_fence_v_lo,icache_yumi_li,
  redirect_resume_li,assembled_v_lo,assembled_partial_lo,assembled_yumi_li,fetch_v_lo,
  fetch_partial_lo,N0,N1,N2,N3,N4;
  wire [1:0] shadow_priv_n,shadow_priv_r;
  wire [38:0] attaboy_pc_li,redirect_pc_li,redirect_npc_li,next_pc_lo,if2_pc_lo,fetch_pc_lo,
  assembled_pc_lo;
  wire [48:0] attaboy_br_metadata_fwd_li,redirect_br_metadata_fwd_li,if2_br_metadata_fwd_lo,
  assembled_br_metadata_fwd_lo,fetch_br_metadata_fwd_lo;
  wire [63:0] icache_data_lo,if2_data_lo;
  wire [2:0] fetch_count_lo,assembled_count_lo,assembled_count_li;
  wire [124:0] fetch_scan_lo;
  wire [26:0] itlb_w_vtag_li;
  wire [35:0] itlb_w_tlb_entry_li;
  wire [27:0] ptag_lo;
  wire [71:0] icache_pkt_li;
  wire [15:0] redirect_instr_li;
  wire [79:0] assembled_instr_lo,fetch_instr_lo;

  bsg_dff_reset_en_bypass_width_p2
  shadow_priv_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(shadow_priv_w),
    .data_i(shadow_priv_n),
    .data_o(shadow_priv_r)
  );


  bsg_dff_reset_en_bypass_width_p1
  shadow_translation_en_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(shadow_translation_en_w),
    .data_i(shadow_translation_en_n),
    .data_o(shadow_translation_en_r)
  );


  bp_fe_pc_gen_00
  pc_gen
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .init_done_o(pc_gen_init_done_lo),
    .attaboy_v_i(attaboy_v_li),
    .attaboy_force_i(attaboy_force_li),
    .attaboy_pc_i(attaboy_pc_li),
    .attaboy_br_metadata_fwd_i(attaboy_br_metadata_fwd_li),
    .attaboy_taken_i(attaboy_taken_li),
    .attaboy_ntaken_i(attaboy_ntaken_li),
    .attaboy_yumi_o(attaboy_yumi_lo),
    .redirect_v_i(redirect_v_li),
    .redirect_pc_i(redirect_pc_li),
    .redirect_npc_i(redirect_npc_li),
    .redirect_br_v_i(redirect_br_v_li),
    .redirect_br_metadata_fwd_i(redirect_br_metadata_fwd_li),
    .redirect_br_taken_i(redirect_br_taken_li),
    .redirect_br_ntaken_i(redirect_br_ntaken_li),
    .redirect_br_nonbr_i(redirect_br_nonbr_li),
    .next_pc_o(next_pc_lo),
    .icache_yumi_i(icache_yumi_lo),
    .ovr_o(ovr_lo),
    .icache_tv_we_i(icache_tv_we),
    .icache_hit_v_i(icache_hit_v_lo),
    .icache_miss_v_i(icache_miss_v_lo),
    .icache_hit_yumi_o(icache_hit_yumi_li),
    .icache_data_i(icache_data_lo),
    .if2_hit_v_o(if2_hit_v_lo),
    .if2_miss_v_o(if2_miss_v_lo),
    .if2_pc_o(if2_pc_lo),
    .if2_data_o(if2_data_lo),
    .if2_br_metadata_fwd_o(if2_br_metadata_fwd_lo),
    .if2_yumi_i(if2_yumi_li),
    .fetch_yumi_i(fetch_yumi_li),
    .fetch_scan_i(fetch_scan_lo),
    .fetch_pc_i(fetch_pc_lo),
    .fetch_count_i(fetch_count_lo),
    .fetch_startup_i(fetch_startup_lo),
    .fetch_catchup_i(fetch_catchup_lo),
    .fetch_rebase_i(fetch_rebase_lo),
    .fetch_linear_i(fetch_linear_lo),
    .fetch_taken_o(fetch_taken_li)
  );


  bp_mmu_00_00000008_00000002_00000001_1
  immu
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .flush_i(tv_flush_lo),
    .fence_i(itlb_fence_v_li),
    .priv_mode_i(shadow_priv_r),
    .trans_en_i(shadow_translation_en_r),
    .sum_i(1'b0),
    .mxr_i(1'b0),
    .uncached_mode_i(N1),
    .nonspec_mode_i(N4),
    .hio_mask_i(cfg_bus_i[9:3]),
    .w_v_i(itlb_w_v_li),
    .w_vtag_i(itlb_w_vtag_li),
    .w_entry_i(itlb_w_tlb_entry_li),
    .r_v_i(itlb_r_v_li),
    .r_instr_i(1'b1),
    .r_load_i(1'b0),
    .r_store_i(1'b0),
    .r_eaddr_i({ next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo[38:38], next_pc_lo }),
    .r_size_i({ 1'b1, 1'b0 }),
    .r_cbo_i(1'b0),
    .r_ptw_i(1'b0),
    .r_v_o(ptag_v_lo),
    .r_ptag_o(ptag_lo),
    .r_instr_miss_o(ptag_miss_lo),
    .r_uncached_o(ptag_uncached_lo),
    .r_nonidem_o(ptag_nonidem_lo),
    .r_dram_o(ptag_dram_lo),
    .r_instr_access_fault_o(instr_access_fault_lo),
    .r_instr_page_fault_o(instr_page_fault_lo)
  );


  bp_fe_icache_00
  icache
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .cfg_bus_i(cfg_bus_i),
    .icache_pkt_i(icache_pkt_li),
    .v_i(icache_v_li),
    .force_i(icache_force_li),
    .yumi_o(icache_yumi_lo),
    .tl_flush_i(tl_flush_lo),
    .ptag_i(ptag_lo),
    .ptag_v_i(ptag_v_lo),
    .ptag_uncached_i(ptag_uncached_lo),
    .ptag_nonidem_i(ptag_nonidem_lo),
    .ptag_dram_i(ptag_dram_lo),
    .tv_flush_i(tv_flush_lo),
    .tv_we_o(icache_tv_we),
    .data_o(icache_data_lo),
    .hit_v_o(icache_hit_v_lo),
    .miss_v_o(icache_miss_v_lo),
    .fence_v_o(icache_fence_v_lo),
    .yumi_i(icache_yumi_li),
    .cache_req_o(cache_req_o),
    .cache_req_v_o(cache_req_v_o),
    .cache_req_yumi_i(cache_req_yumi_i),
    .cache_req_lock_i(cache_req_lock_i),
    .cache_req_metadata_o(cache_req_metadata_o),
    .cache_req_metadata_v_o(cache_req_metadata_v_o),
    .cache_req_id_i(cache_req_id_i[0]),
    .cache_req_critical_i(cache_req_critical_i),
    .cache_req_last_i(cache_req_last_i),
    .cache_req_credits_full_i(cache_req_credits_full_i),
    .cache_req_credits_empty_i(cache_req_credits_empty_i),
    .data_mem_pkt_v_i(data_mem_pkt_v_i),
    .data_mem_pkt_i(data_mem_pkt_i),
    .data_mem_pkt_yumi_o(data_mem_pkt_yumi_o),
    .data_mem_o(data_mem_o),
    .tag_mem_pkt_v_i(tag_mem_pkt_v_i),
    .tag_mem_pkt_i(tag_mem_pkt_i),
    .tag_mem_pkt_yumi_o(tag_mem_pkt_yumi_o),
    .tag_mem_o(tag_mem_o),
    .stat_mem_pkt_v_i(stat_mem_pkt_v_i),
    .stat_mem_pkt_i(stat_mem_pkt_i),
    .stat_mem_pkt_yumi_o(stat_mem_pkt_yumi_o),
    .stat_mem_o(stat_mem_o)
  );


  bp_fe_realigner_00
  realigner
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .if2_hit_v_i(if2_hit_v_lo),
    .if2_miss_v_i(if2_miss_v_lo),
    .if2_pc_i(if2_pc_lo),
    .if2_data_i(if2_data_lo),
    .if2_br_metadata_fwd_i(if2_br_metadata_fwd_lo),
    .if2_yumi_o(if2_yumi_li),
    .redirect_v_i(redirect_v_li),
    .redirect_pc_i(redirect_pc_li),
    .redirect_instr_i(redirect_instr_li),
    .redirect_br_metadata_fwd_i(redirect_br_metadata_fwd_li),
    .redirect_resume_i(redirect_resume_li),
    .assembled_v_o(assembled_v_lo),
    .assembled_pc_o(assembled_pc_lo),
    .assembled_instr_o(assembled_instr_lo),
    .assembled_br_metadata_fwd_o(assembled_br_metadata_fwd_lo),
    .assembled_count_o(assembled_count_lo),
    .assembled_partial_o(assembled_partial_lo),
    .assembled_count_i(assembled_count_li),
    .assembled_yumi_i(assembled_yumi_li)
  );


  bp_fe_scan_00
  scan
  (
    .assembled_v_i(assembled_v_lo),
    .assembled_pc_i(assembled_pc_lo),
    .assembled_instr_i(assembled_instr_lo),
    .assembled_br_metadata_fwd_i(assembled_br_metadata_fwd_lo),
    .assembled_count_i(assembled_count_lo),
    .assembled_partial_i(assembled_partial_lo),
    .assembled_count_o(assembled_count_li),
    .assembled_yumi_o(assembled_yumi_li),
    .fetch_v_o(fetch_v_lo),
    .fetch_pc_o(fetch_pc_lo),
    .fetch_instr_o(fetch_instr_lo),
    .fetch_br_metadata_fwd_o(fetch_br_metadata_fwd_lo),
    .fetch_count_o(fetch_count_lo),
    .fetch_partial_o(fetch_partial_lo),
    .fetch_scan_o(fetch_scan_lo),
    .fetch_startup_o(fetch_startup_lo),
    .fetch_catchup_o(fetch_catchup_lo),
    .fetch_rebase_o(fetch_rebase_lo),
    .fetch_linear_o(fetch_linear_lo),
    .fetch_taken_i(fetch_taken_li),
    .fetch_yumi_i(fetch_yumi_li)
  );


  bp_fe_controller_00
  controller
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .pc_gen_init_done_i(pc_gen_init_done_lo),
    .fe_cmd_i(fe_cmd_i),
    .fe_cmd_v_i(fe_cmd_v_i),
    .fe_cmd_yumi_o(fe_cmd_yumi_o),
    .fe_queue_o(fe_queue_o),
    .fe_queue_v_o(fe_queue_v_o),
    .fe_queue_ready_and_i(fe_queue_ready_and_i),
    .redirect_v_o(redirect_v_li),
    .redirect_pc_o(redirect_pc_li),
    .redirect_npc_o(redirect_npc_li),
    .redirect_instr_o(redirect_instr_li),
    .redirect_resume_o(redirect_resume_li),
    .redirect_br_v_o(redirect_br_v_li),
    .redirect_br_taken_o(redirect_br_taken_li),
    .redirect_br_ntaken_o(redirect_br_ntaken_li),
    .redirect_br_nonbr_o(redirect_br_nonbr_li),
    .redirect_br_metadata_fwd_o(redirect_br_metadata_fwd_li),
    .attaboy_v_o(attaboy_v_li),
    .attaboy_force_o(attaboy_force_li),
    .attaboy_pc_o(attaboy_pc_li),
    .attaboy_taken_o(attaboy_taken_li),
    .attaboy_ntaken_o(attaboy_ntaken_li),
    .attaboy_br_metadata_fwd_o(attaboy_br_metadata_fwd_li),
    .attaboy_yumi_i(attaboy_yumi_lo),
    .next_pc_i(next_pc_lo),
    .ovr_i(ovr_lo),
    .tl_flush_o(tl_flush_lo),
    .tv_we_i(icache_tv_we),
    .itlb_miss_tl_i(ptag_miss_lo),
    .instr_page_fault_tl_i(instr_page_fault_lo),
    .instr_access_fault_tl_i(instr_access_fault_lo),
    .icache_miss_tv_i(icache_miss_v_lo),
    .tv_flush_o(tv_flush_lo),
    .fetch_v_i(fetch_v_lo),
    .fetch_pc_i(fetch_pc_lo),
    .fetch_instr_i(fetch_instr_lo),
    .fetch_count_i(fetch_count_lo),
    .fetch_partial_i(fetch_partial_lo),
    .fetch_br_metadata_fwd_i(fetch_br_metadata_fwd_lo),
    .fetch_yumi_o(fetch_yumi_li),
    .itlb_r_v_o(itlb_r_v_li),
    .itlb_w_v_o(itlb_w_v_li),
    .itlb_w_vtag_o(itlb_w_vtag_li),
    .itlb_w_entry_o(itlb_w_tlb_entry_li),
    .itlb_fence_v_o(itlb_fence_v_li),
    .icache_v_o(icache_v_li),
    .icache_force_o(icache_force_li),
    .icache_pkt_o(icache_pkt_li),
    .icache_yumi_i(icache_yumi_lo),
    .shadow_priv_w_o(shadow_priv_w),
    .shadow_priv_o(shadow_priv_n),
    .shadow_translation_en_w_o(shadow_translation_en_w),
    .shadow_translation_en_o(shadow_translation_en_n)
  );

  assign N0 = cfg_bus_i[16] | cfg_bus_i[17];
  assign N1 = ~N0;
  assign N2 = ~cfg_bus_i[17];
  assign N3 = cfg_bus_i[16] | N2;
  assign N4 = ~N3;
  assign icache_yumi_li = icache_hit_yumi_li | icache_fence_v_lo;

endmodule

