`ifndef BSG_DEFINES_V
`define BSG_DEFINES_V

`define BSG_MAX(x,y) (((x)>(y)) ? (x) : (y))
`define BSG_MIN(x,y) (((x)<(y)) ? (x) : (y))

`define BSG_SIGN_EXTEND(sig, width) \
  ({{`BSG_MAX(width-$bits(sig),0){sig[$bits(sig)-1]}}, sig[0+:`BSG_MIN(width, $bits(sig))]})
`define BSG_ZERO_EXTEND(sig, width) \
  ({{`BSG_MAX(width-$bits(sig),0){1'b0}}, sig[0+:`BSG_MIN(width, $bits(sig))]})

// place this macro at the end of a verilog module file if that module has invalid parameters
// that must be specified by the user. this will prevent that module from becoming a top-level
// module per the discussion here: https://github.com/SymbiFlow/sv-tests/issues/1160 and the
// SystemVerilog Standard

//    "Top-level modules are modules that are included in the SystemVerilog
//    source text, but do not appear in any module instantiation statement, as
//    described in 23.3.2. This applies even if the module instantiation appears
//    in a generate block that is not itself instantiated (see 27.3). A design
//    shall contain at least one top-level module. A top-level module is
//    implicitly instantiated once, and its instance name is the same as the
//    module name. Such an instance is called a top-level instance."
//  

`define BSG_ABSTRACT_MODULE(fn) \
    /*verilator lint_off DECLFILENAME*/ \
    /*verilator lint_off PINMISSING*/ \
    module fn``__abstract(); if (0) begin : abstract fn not_used(); end endmodule \
    /*verilator lint_on PINMISSING*/ \
    /*verilator lint_on DECLFILENAME*/

// macro for defining invalid parameter; with the abstract module declaration
// it should be sufficient to omit the "inv" but we include this for tool portability
// if later we find that all tools are compatible, we can remove the use of this from BaseJump STL

`ifdef XCELIUM // Bare default parameters are incompatible as of 20.09.012
               // = "inv" causes type inference mismatch as of 20.09.012
`define BSG_INV_PARAM(param) param = -1
`elsif YOSYS // Bare default parameters are incompatible as of 0.9
`define BSG_INV_PARAM(param) param = "inv"
`else // VIVADO, DC, VERILATOR, GENUS, SURELOG
`define BSG_INV_PARAM(param) param
`endif


// maps 1 --> 1 instead of to 0
`define BSG_SAFE_CLOG2(x) ( (((x)==1) || ((x)==0))? 1 : $clog2((x)))
`define BSG_IS_POW2(x) ( (1 << $clog2(x)) == (x))
`define BSG_WIDTH(x) ($clog2(x+1))
`define BSG_SAFE_MINUS(x, y) (((x)<(y))) ? 0 : ((x)-(y))

// calculate ceil(x/y) 
`define BSG_CDIV(x,y) (((x)+(y)-1)/(y))

`ifdef SYNTHESIS
`define BSG_UNDEFINED_IN_SIM(val) (val)
`else
`define BSG_UNDEFINED_IN_SIM(val) ('X)
`endif

`ifdef VERILATOR
`define BSG_HIDE_FROM_VERILATOR(val)
`else
`define BSG_HIDE_FROM_VERILATOR(val) val
`endif

`ifdef SYNTHESIS
`define BSG_DISCONNECTED_IN_SIM(val) (val)
`elsif VERILATOR
`define BSG_DISCONNECTED_IN_SIM(val) (val)
`else
`define BSG_DISCONNECTED_IN_SIM(val) ('z)
`endif

// Ufortunately per the Xilinx forums, Xilinx does not define
// any variable that indicates that Vivado Synthesis is running
// so as a result we identify Vivado merely as the exclusion of
// Synopsys Design Compiler (DC). Support beyond DC and Vivado
// will require modification of this macro.

`ifdef SYNTHESIS
  `ifdef DC
  `define BSG_VIVADO_SYNTH_FAILS
  `elsif CDS_TOOL_DEFINE
  `define BSG_VIVADO_SYNTH_FAILS
  `elsif SURELOG
  `define BSG_VIVADO_SYNTH_FAILS
  `elsif YOSYS
  `define BSG_VIVADO_SYNTH_FAILS
  `else
  `define BSG_VIVADO_SYNTH_FAILS this_module_is_not_synthesizeable_in_vivado
  `endif
`else
`define BSG_VIVADO_SYNTH_FAILS
`endif

// macro for denoting that a code snippet is unsynthesiable

`ifdef SYNTHESIS
  `define BSG_HIDE_FROM_SYNTHESIS
`endif

`define BSG_STRINGIFY(x) `"x`"


// For the modules that must be hardened, add this macro at the top.
`ifdef SYNTHESIS
`define BSG_SYNTH_MUST_HARDEN this_module_must_be_hardened
`else
`define BSG_SYNTH_MUST_HARDEN
`endif


// using C-style shifts instead of a[i] allows the parameter of BSG_GET_BIT to be a parameter subrange                                                                                                                                                                               
// e.g., parameter[4:1][1], which DC 2016.12 does not allow                                                                                                                                                                                                                          

`define BSG_GET_BIT(X,NUM) (((X)>>(NUM))&1'b1)

// This version of countones works in synthesis, but only up to 64 bits                                                                                                                                                                                                              
// we do a funny thing where we propagate X's in simulation if it is more than 64 bits                                                                                                                                                                                               
// and in synthesis, go ahead and ignore the high bits                                                                                                                                                                      

`define BSG_COUNTONES_SYNTH(y) (($bits(y) < 65) ? 1'b0 : `BSG_UNDEFINED_IN_SIM(1'b0)) + (`BSG_GET_BIT(y,0) +`BSG_GET_BIT(y,1) +`BSG_GET_BIT(y,2) +`BSG_GET_BIT(y,3) +`BSG_GET_BIT(y,4) +`BSG_GET_BIT(y,5) +`BSG_GET_BIT(y,6)+`BSG_GET_BIT(y,7) +`BSG_GET_BIT(y,8)+`BSG_GET_BIT(y,9) \
                                                                                       +`BSG_GET_BIT(y,10)+`BSG_GET_BIT(y,11)+`BSG_GET_BIT(y,12)+`BSG_GET_BIT(y,13)+`BSG_GET_BIT(y,14)+`BSG_GET_BIT(y,15)+`BSG_GET_BIT(y,16)+`BSG_GET_BIT(y,17)+`BSG_GET_BIT(y,18)+`BSG_GET_BIT(y,19) \
                                                                                       +`BSG_GET_BIT(y,20)+`BSG_GET_BIT(y,21)+`BSG_GET_BIT(y,22)+`BSG_GET_BIT(y,23)+`BSG_GET_BIT(y,24)+`BSG_GET_BIT(y,25)+`BSG_GET_BIT(y,26)+`BSG_GET_BIT(y,27)+`BSG_GET_BIT(y,28)+`BSG_GET_BIT(y,29) \
                                                                                       +`BSG_GET_BIT(y,30)+`BSG_GET_BIT(y,31)+`BSG_GET_BIT(y,32)+`BSG_GET_BIT(y,33)+`BSG_GET_BIT(y,34)+`BSG_GET_BIT(y,35)+`BSG_GET_BIT(y,36)+`BSG_GET_BIT(y,37)+`BSG_GET_BIT(y,38)+`BSG_GET_BIT(y,39) \
                                                                                       +`BSG_GET_BIT(y,40)+`BSG_GET_BIT(y,41)+`BSG_GET_BIT(y,42)+`BSG_GET_BIT(y,43)+`BSG_GET_BIT(y,44)+`BSG_GET_BIT(y,45)+`BSG_GET_BIT(y,46)+`BSG_GET_BIT(y,47)+`BSG_GET_BIT(y,48)+`BSG_GET_BIT(y,49) \
                                                                                       +`BSG_GET_BIT(y,50)+`BSG_GET_BIT(y,51)+`BSG_GET_BIT(y,52)+`BSG_GET_BIT(y,53)+`BSG_GET_BIT(y,54)+`BSG_GET_BIT(y,55)+`BSG_GET_BIT(y,56)+`BSG_GET_BIT(y,57)+`BSG_GET_BIT(y,58)+`BSG_GET_BIT(y,59) \
                                                                                       +`BSG_GET_BIT(y,60)+`BSG_GET_BIT(y,61)+`BSG_GET_BIT(y,62)+`BSG_GET_BIT(y,63))

// nullify rpgroups
`ifndef rpgroup
`define rpgroup(x)
`endif

// verilog preprocessing -> if defined(A) && defined(B) then define C
`define BSG_DEFIF_A_AND_B(A,B,C) \
    `undef C \
    `ifdef A \
        `ifdef B \
            `define C \
        `endif \
    `endif

// verilog preprocessing -> if defined(A) && !defined(B) then define C
`define BSG_DEFIF_A_AND_NOT_B(A,B,C) \
    `undef C \
    `ifdef A \
        `ifndef B \
            `define C \
        `endif \
    `endif

// verilog preprocessing -> if !defined(A) && defined(B) then define C
`define BSG_DEFIF_NOT_A_AND_B(A,B,C) `BSG_DEFIF_A_AND_NOT_B(B,A,C)

// verilog preprocessing -> if !defined(A) && !defined(B) then define C
`define BSG_DEFIF_NOT_A_AND_NOT_B(A,B,C) \
    `undef C \
    `ifndef A \
        `ifndef B \
            `define C \
        `endif \
    `endif

// verilog preprocessing -> if defined(A) || defined(B) then define C
`define BSG_DEFIF_A_OR_B(A,B,C) \
    `undef C \
    `ifdef A \
        `define C \
    `endif \
    `ifdef B \
        `define C \
    `endif

// verilog preprocessing -> if defined(A) || !defined(B) then define C
`define BSG_DEFIF_A_OR_NOT_B(A,B,C) \
    `undef C \
    `ifdef A \
        `define C \
    `endif \
    `ifndef B \
        `define C \
    `endif

// verilog preprocessing -> if !defined(A) || defined(B) then define C
`define BSG_DEFIF_NOT_A_OR_B(A,B,C) `BSG_DEFIF_A_OR_NOT_B(B,A,C)

// verilog preprocessing -> if !defined(A) || !defined(B) then define C
`define BSG_DEFIF_NOT_A_OR_NOT_B(A,B,C) \
    `undef C \
    `ifndef A \
        `define C \
    `endif \
    `ifndef B \
        `define C \
    `endif

`endif
// MBT 7/7/2016
//
// 1 read-port, 1 write-port ram
//
// reads are synchronous
//
// NOTE: Users of BaseJump STL should not instantiate this module directly
// they should use bsg_mem_1r1w_sync_mask_write_bit.


//`include "bsg_defines.sv"

module bsg_mem_1r1w_sync_mask_write_bit_synth #(parameter `BSG_INV_PARAM(width_p)
						, parameter `BSG_INV_PARAM(els_p)
						, parameter read_write_same_addr_p=0
						, parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
                                                , parameter latch_last_read_p=0
                                                , parameter disable_collision_warning_p=1
                                        )
   (input   clk_i
    , input reset_i

    , input                     w_v_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0]       w_mask_i
    , input [addr_width_lp-1:0] w_addr_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0]       w_data_i

    // currently unused
    , input                      r_v_i
    , input [addr_width_lp-1:0]  r_addr_i

    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r_data_o
    );

   wire                   unused = reset_i;

   if (width_p == 0)
    begin: z
      wire unused0 = &{clk_i, w_v_i, w_mask_i, w_addr_i, r_v_i, r_addr_i};
      assign r_data_o = '0;
    end
   else
    begin: nz

   logic [width_p-1:0]    mem [els_p-1:0];
   logic read_en;
   logic [width_p-1:0] data_out;

   // this treats the ram as an array of registers for which the
   // read addr is latched on the clock, the write
   // is done on the clock edge, and actually multiplexing
   // of the registers for reading is done after the clock edge.

   // logically, this means that reads happen in time after
   // the writes, and "simultaneous" reads and writes to the
   // register file are allowed -- IF read_write_same_addr is set.

   // note that this behavior is generally incompatible with
   // hardened 1r1w rams, so it's better not to take advantage
   // of it if not necessary

   // we explicitly 'X out the read address if valid is not set
   // to avoid accidental use of data when the valid signal was not
   // asserted. without this, the output of the register file would
   // "auto-update" based on new writes to the ram, a spooky behavior
   // that would never correspond to that of a hardened ram.

   logic [addr_width_lp-1:0] r_addr_r;

   assign read_en = r_v_i;
   assign data_out = mem[r_addr_r];


   always_ff @(posedge clk_i)
     begin
        if (r_v_i)
          r_addr_r <= r_addr_i;

`ifndef BSG_HIDE_FROM_SYNTHESIS
        else
          r_addr_r <= 'X;

        // if addresses match and this is forbidden, then nuke the read address

        if (r_addr_i == w_addr_i && w_v_i && r_v_i && !read_write_same_addr_p)
          begin
             if (!disable_collision_warning_p)
               begin
                 $error("X'ing matched read address %x (%m)",r_addr_i);
               end
             r_addr_r <= 'X;
          end
`endif

     end

  if (latch_last_read_p)
    begin: llr
      logic read_en_r; 

      bsg_dff #(
        .width_p(1)
      ) read_en_dff (
        .clk_i(clk_i)
        ,.data_i(read_en)
        ,.data_o(read_en_r)
      );

      bsg_dff_en_bypass #(
        .width_p(width_p)
      ) dff_bypass (
        .clk_i(clk_i)
        ,.en_i(read_en_r)
        ,.data_i(data_out)
        ,.data_o(r_data_o)
      );
    end
  else
    begin: no_llr
      assign r_data_o = data_out;
    end

   genvar                       i;
   for (i = 0; i < width_p; i=i+1)
     begin
	always_ff @(posedge clk_i)

	  if (w_v_i && w_mask_i[i])
            mem[w_addr_i][i] <= w_data_i[i];
     end
  end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_1r1w_sync_mask_write_bit_synth)
// MBT 7/7/2016
//
// 1 read-port, 1 write-port ram
//
// reads are synchronous
//
// NOTE: Users of BaseJump STL should not instantiate this module directly
// they should use bsg_mem_1r1w_sync_mask_write_bit.


//`include "bsg_defines.sv"

module bsg_mem_1r1w_sync_mask_write_byte_synth #(parameter `BSG_INV_PARAM(width_p)
						, parameter `BSG_INV_PARAM(els_p)
						, parameter read_write_same_addr_p=0
						, parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
                                                , parameter latch_last_read_p=0
                                                , parameter write_mask_width_lp = width_p>>3
						, parameter harden_p=0
                                                , parameter disable_collision_warning_p=1
                                        )
   (input   clk_i
    , input reset_i

    , input                     w_v_i
    // for each bit set in the mask, a byte is written
    , input [`BSG_SAFE_MINUS(write_mask_width_lp, 1):0] w_mask_i
    , input [addr_width_lp-1:0] w_addr_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0]       w_data_i

    // currently unused
    , input                      r_v_i
    , input [addr_width_lp-1:0]  r_addr_i

    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r_data_o
    );

   wire                   unused = reset_i;

   if (width_p == 0)
    begin: z
      wire unused0 = &{clk_i, w_v_i, w_mask_i, w_addr_i, r_v_i, r_addr_i};
      assign r_data_o = '0;
    end
   else
    begin: nz

  for(genvar i=0; i<write_mask_width_lp; i=i+1)
  begin: bk
    bsg_mem_1r1w_sync #( .width_p      (8)
                        ,.els_p        (els_p)
                        ,.addr_width_lp(addr_width_lp)
                        ,.latch_last_read_p(latch_last_read_p)
			,.verbose_if_synth_p(0) // don't print out details of ram if breaks into synth srams
                      ) mem_1r1w_sync
                      ( .clk_i  (clk_i)
                       ,.reset_i(reset_i)
                       ,.w_v_i    (w_v_i & w_mask_i[i])
                       ,.w_data_i (w_data_i[(i*8)+:8])
                       ,.w_addr_i (w_addr_i)
                       ,.r_v_i    (r_v_i)
                       ,.r_addr_i (r_addr_i)
                       ,.r_data_o (r_data_o[(i*8)+:8])
                      );
  end
   end

endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_1r1w_sync_mask_write_byte_synth)

// MBT 7/7/2016
//
// 1 read-port, 1 write-port ram
//
// reads are synchronous
//
// although we could merge this with normal bsg_mem_1r1w
// and select with a parameter, we do not do this because
// it's typically a very big change to the instantiating code
// to move to/from sync/async, and we want to reflect this.
//
// NOTE: Users of BaseJump STL should not instantiate this module directly
// they should use bsg_mem_1r1w_sync.

//`include "bsg_defines.sv"

module bsg_mem_1r1w_sync_synth #(parameter `BSG_INV_PARAM(width_p)
				 , parameter `BSG_INV_PARAM(els_p)
				 , parameter read_write_same_addr_p=0
				 , parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
                                 , parameter latch_last_read_p=0
                 , parameter verbose_p=1
				 )
   (input   clk_i
    , input reset_i

    , input                     w_v_i
    , input [addr_width_lp-1:0] w_addr_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0]       w_data_i

    // currently unused
    , input                      r_v_i
    , input [addr_width_lp-1:0]  r_addr_i

    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r_data_o
    );

   wire                   unused = reset_i;

   if (width_p == 0 || els_p == 0)
    begin: z
      wire unused0 = &{clk_i, w_v_i, w_addr_i, r_v_i, r_addr_i};
      assign r_data_o = '0;
    end
   else
    begin: nz

   logic [width_p-1:0]    mem [els_p-1:0];
   logic read_en;
   logic [width_p-1:0] data_out;

   // this treats the ram as an array of registers for which the
   // read addr is latched on the clock, the write
   // is done on the clock edge, and actually multiplexing
   // of the registers for reading is done after the clock edge.

   // logically, this means that reads happen in time after
   // the writes, and "simultaneous" reads and writes to the
   // register file are allowed -- IF read_write_same_addr is set.

   // note that this behavior is generally incompatible with
   // hardened 1r1w rams, so it's better not to take advantage
   // of it if not necessary

   // we explicitly 'X out the read address if valid is not set
   // to avoid accidental use of data when the valid signal was not
   // asserted. without this, the output of the register file would
   // "auto-update" based on new writes to the ram, a spooky behavior
   // that would never correspond to that of a hardened ram.

   logic [addr_width_lp-1:0] r_addr_r;
   wire [addr_width_lp-1:0] r_addr_li = (els_p > 1) ? r_addr_i:'0;
   wire [addr_width_lp-1:0] w_addr_li = (els_p > 1) ? w_addr_i:'0;

   assign read_en = r_v_i;
   assign data_out = mem[r_addr_r];

   always_ff @(posedge clk_i)
     if (r_v_i)
       r_addr_r <= r_addr_li;
     else
       r_addr_r <= 'X;

  if (latch_last_read_p)
    begin: llr
      logic read_en_r; 

      bsg_dff #(
        .width_p(1)
      ) read_en_dff (
        .clk_i(clk_i)
        ,.data_i(read_en)
        ,.data_o(read_en_r)
      );

      bsg_dff_en_bypass #(
        .width_p(width_p)
      ) dff_bypass (
        .clk_i(clk_i)
        ,.en_i(read_en_r)
        ,.data_i(data_out)
        ,.data_o(r_data_o)
      );
    end
  else
    begin: no_llr
      assign r_data_o = data_out;
    end

   always_ff @(posedge clk_i)
     if (w_v_i)
       mem[w_addr_li] <= w_data_i;

   end

`ifndef BSG_HIDE_FROM_SYNTHESIS
   initial
     begin
        if (verbose_p)
      $display("## %L: instantiating width_p=%d, els_p=%d (%m)",width_p,els_p);
     end
`endif

endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_1r1w_sync_synth)// MBT
//
// 1 read-port, 1 write-port ram
//
// reads are asynchronous
//
// for synthesizable internal version, we omit assertions
// these should be placed in the outer wrapper
//

//`include "bsg_defines.sv"

module bsg_mem_1r1w_synth #(parameter `BSG_INV_PARAM(width_p)
			    ,parameter `BSG_INV_PARAM(els_p)
			    ,parameter read_write_same_addr_p=0
			    ,parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p))
(
  input w_clk_i
  ,input w_reset_i

  ,input w_v_i
  ,input [addr_width_lp-1:0] w_addr_i
  ,input [`BSG_SAFE_MINUS(width_p, 1):0] w_data_i

  // currently unused
  ,input r_v_i
  ,input [addr_width_lp-1:0]  r_addr_i

  ,output logic [`BSG_SAFE_MINUS(width_p, 1):0] r_data_o
);

  wire unused0 = w_reset_i;
  wire unused1 = r_v_i;

  if (width_p == 0 || els_p == 0)
   begin: z
     wire unused2 = &{w_clk_i, w_addr_i, w_data_i, r_addr_i};
     assign r_data_o = '0;
   end
  else
   begin: nz

  logic [width_p-1:0] mem [els_p-1:0];

  wire [addr_width_lp-1:0] r_addr_li = (els_p > 0) ? r_addr_i:'0;
  wire [addr_width_lp-1:0] w_addr_li = (els_p > 0) ? w_addr_i:'0;

  // this implementation ignores the r_v_i
  assign r_data_o = mem[r_addr_li];

  always_ff @(posedge w_clk_i) begin
    if (w_v_i) begin
      mem[w_addr_li] <= w_data_i;
    end
  end
   end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_1r1w_synth)
// MBT 11/9/2014
//
// Synchronous 1-port ram.
// Only one read or one write may be done per cycle.
//
// NOTE: Users of BaseJump STL should not instantiate this module directly
// they should use bsg_mem_1rw_sync_mask_write_bit.
//

//`include "bsg_defines.sv"

module bsg_mem_1rw_sync_mask_write_bit_synth
  #(parameter `BSG_INV_PARAM(width_p)
    , parameter `BSG_INV_PARAM(els_p)
    , parameter latch_last_read_p=0
    , parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
   )
   (input   clk_i
    , input reset_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0] data_i
    , input [addr_width_lp-1:0] addr_i
    , input v_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0] w_mask_i
    , input w_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0]  data_o
    );

   wire unused = reset_i;

   if (width_p == 0 || els_p == 0)
    begin: z
      wire unused0 = &{clk_i, data_i, addr_i, v_i, w_mask_i, w_i};
      assign data_o = '0;
    end
   else
    begin: nz

   logic [addr_width_lp-1:0] addr_r;
   logic [width_p-1:0] mem [els_p-1:0];
   logic read_en;
   
   wire [addr_width_lp-1:0] addr_li = (els_p>1) ? addr_i:'0;
   
   assign read_en = v_i & ~w_i;

   always_ff @(posedge clk_i)
     if (read_en)
       addr_r <= addr_li;
     else
       addr_r <= 'X;

   logic [width_p-1:0] data_out;

   assign data_out = mem[addr_r];

   if (latch_last_read_p)
     begin: llr
      logic read_en_r; 

      bsg_dff #(
        .width_p(1)
      ) read_en_dff (
        .clk_i(clk_i)
        ,.data_i(read_en)
        ,.data_o(read_en_r)
      );

      bsg_dff_en_bypass #(
        .width_p(width_p)
      ) dff_bypass (
        .clk_i(clk_i)
        ,.en_i(read_en_r)
        ,.data_i(data_out)
        ,.data_o(data_o)
      );
     end
   else
     begin: no_llr
       assign data_o = data_out;
     end



// The Verilator and non-Verilator models are functionally equivalent. However, Verilator
//   cannot handle an array of non-blocking assignments in a for loop. It would be nice to 
//   see if these two models synthesize the same, because we can then reduce to the Verilator
//   model and avoid double maintenence. One could also add this feature to Verilator...
//   (Identified in Verilator 4.011)
`ifdef VERILATOR
   logic [width_p-1:0] data_n;

   for (genvar i = 0; i < width_p; i++)
     begin : rof1
       assign data_n[i] = w_mask_i[i] ? data_i[i] : mem[addr_li][i];
     end // rof1

   always_ff @(posedge clk_i)
     if (v_i & w_i)
       mem[addr_li] <= data_n;

`else
 
// this code does not map correctly with Xilinx Ultrascale FPGAs 
// in Vivado, substitute this file with hard/ultrascale_plus/bsg_mem/bsg_mem_1rw_sync_mask_write_bit.sv
      
`BSG_VIVADO_SYNTH_FAILS
      
   always_ff @(posedge clk_i)
     if (v_i & w_i)
       for (integer i = 0; i < width_p; i=i+1)
         if (w_mask_i[i])
           mem[addr_li][i] <= data_i[i];
`endif
   end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_1rw_sync_mask_write_bit_synth)
// NOTE: Users of BaseJump STL should not instantiate this module directly
// they should use bsg_mem_1r1w_sync_mask_write_byte.

//`include "bsg_defines.sv"

module bsg_mem_1rw_sync_mask_write_byte_synth
  #(parameter `BSG_INV_PARAM(els_p)
    , parameter addr_width_lp = `BSG_SAFE_CLOG2(els_p)
    , parameter latch_last_read_p=0

    , parameter `BSG_INV_PARAM(data_width_p )
    , parameter write_mask_width_lp = data_width_p>>3
  )
  ( input clk_i
   ,input reset_i

   ,input v_i
   ,input w_i

   ,input [addr_width_lp-1:0]       addr_i
   ,input [`BSG_SAFE_MINUS(data_width_p, 1):0]        data_i
    // for each bit set in the mask, a byte is written
   ,input [`BSG_SAFE_MINUS(write_mask_width_lp, 1):0] write_mask_i

   ,output [`BSG_SAFE_MINUS(data_width_p, 1):0] data_o
  );

  genvar i;

  if (data_width_p == 0 || els_p == 0)
   begin: z
     wire unused0 = &{clk_i, reset_i, v_i, w_i, addr_i, data_i, write_mask_i};
     assign data_o = '0;
   end
  else
   begin: nz

  for(i=0; i<write_mask_width_lp; i=i+1)
  begin: bk
    bsg_mem_1rw_sync #( .width_p      (8)
                        ,.els_p        (els_p)
                        ,.addr_width_lp(addr_width_lp)
                        ,.latch_last_read_p(latch_last_read_p)
			,.verbose_if_synth_p(0) // don't print out details of ram if breaks into synth srams
                      ) mem_1rw_sync
                      ( .clk_i  (clk_i)
                       ,.reset_i(reset_i)
                       ,.data_i (data_i[(i*8)+:8])
                       ,.addr_i (addr_i)
                       ,.v_i    (v_i & (w_i ? write_mask_i[i] : 1'b1))
                       ,.w_i    (w_i & write_mask_i[i])
                       ,.data_o (data_o[(i*8)+:8])
                      );
  end
   end

endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_1rw_sync_mask_write_byte_synth)
// MBT 11/9/2014
//
// Synchronous 1-port ram.
// Only one read or one write may be done per cycle.
//
// NOTE: Users of BaseJump STL should not instantiate this module directly
// they should use bsg_mem_1rw_sync.

//`include "bsg_defines.sv"

module bsg_mem_1rw_sync_synth
  #(parameter `BSG_INV_PARAM(width_p)
    , parameter `BSG_INV_PARAM(els_p)
    , parameter latch_last_read_p=0
    , parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
    , parameter verbose_p=1
   )
   (input   clk_i
	 	, input v_i
		, input reset_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0] data_i
    , input [addr_width_lp-1:0] addr_i
    , input w_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0]  data_o
    );

  wire unused = reset_i;

  if (width_p == 0 || els_p == 0)
   begin: z
     wire unused0 = &{clk_i, v_i, data_i, addr_i, w_i};
     assign data_o = '0;
   end
  else
   begin: nz

    logic [addr_width_lp-1:0] addr_r;
    logic [width_p-1:0]    mem [els_p-1:0];
    logic read_en;
    logic [width_p-1:0] data_out;

    wire [addr_width_lp-1:0] addr_li = (els_p>0) ? addr_i:'0;

    assign read_en = v_i & ~w_i;
    assign data_out = mem[addr_r];

    always_ff @ (posedge clk_i) 
      if (read_en)
        addr_r <= addr_li;
      else
        addr_r <= 'X;

    if (latch_last_read_p)
      begin: llr
        logic read_en_r; 

        bsg_dff #(
          .width_p(1)
        ) read_en_dff (
          .clk_i(clk_i)
          ,.data_i(read_en)
          ,.data_o(read_en_r)
        );

        bsg_dff_en_bypass #(
          .width_p(width_p)
        ) dff_bypass (
          .clk_i(clk_i)
          ,.en_i(read_en_r)
          ,.data_i(data_out)
          ,.data_o(data_o)
        );
      end
    else
      begin: no_llr
        assign data_o = data_out;
      end


    always_ff @(posedge clk_i)
      if (v_i & w_i) 
        mem[addr_li] <= data_i;
   end // non_zero_width
`ifndef BSG_HIDE_FROM_SYNTHESIS
   initial
     begin
        if (verbose_p)
	  $display("## %L: instantiating width_p=%d, els_p=%d (%m)",width_p,els_p);
     end
   

   always_ff @(negedge clk_i)
     if (v_i)
       assert ( (v_i !== 1'b1) || (reset_i === 'X) || (reset_i === 1'b1) || (addr_i < els_p) || (els_p <= 1))
         else $error("Invalid address %x to %m of size %x (reset_i = %b, v_i = %b, clk_i = %b)\n", addr_i, els_p, reset_i, v_i, clk_i);
`endif

endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_1rw_sync_synth)
// MBT 7/7/2016
//
// 2 read-port, 1 write-port ram
//
// reads are synchronous
//
// although we could merge this with normal bsg_mem_1r1w
// and select with a parameter, we do not do this because
// it's typically a very big change to the instantiating code
// to move to/from sync/async, and we want to reflect this.
//
// NOTE: Users of BaseJump STL should not instantiate this module directly
// they should use bsg_mem_2r1w_sync.

//`include "bsg_defines.sv"

module bsg_mem_2r1w_sync_synth #(parameter `BSG_INV_PARAM(width_p)
				 , parameter `BSG_INV_PARAM(els_p)
				 , parameter read_write_same_addr_p=0
				 , parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
				 )
   (input   clk_i
    , input reset_i

    , input                     w_v_i
    , input [addr_width_lp-1:0] w_addr_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0]       w_data_i

    // currently unused
    , input                      r0_v_i
    , input [addr_width_lp-1:0]  r0_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r0_data_o

    , input                      r1_v_i
    , input [addr_width_lp-1:0]  r1_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r1_data_o
    );

   wire                   unused = reset_i;

   if (width_p == 0)
    begin: z
      wire unused0 = &{clk_i, w_v_i, w_addr_i, w_data_i, r0_v_i, r0_addr_i, r1_v_i, r1_addr_i};
      assign r0_data_o = '0;
      assign r1_data_o = '0;
    end
   else
    begin: nz

   logic [width_p-1:0]    mem [els_p-1:0];

   // keep consistent with bsg_ip_cores/bsg_mem/bsg_mem_2r1w_sync.sv
   // keep consistent with bsg_ip_cores/hard/bsg_mem/bsg_mem_2r1w_sync.sv
   
   // this treats the ram as an array of registers for which the
   // read addr is latched on the clock, the write
   // is done on the clock edge, and actually multiplexing
   // of the registers for reading is done after the clock edge.

   // logically, this means that reads happen in time after
   // the writes, and "simultaneous" reads and writes to the
   // register file are allowed -- IF read_write_same_addr is set.

   // note that this behavior is generally incompatible with
   // hardened 1r1w rams, so it's better not to take advantage
   // of it if not necessary

   // we explicitly 'X out the read address if valid is not set
   // to avoid accidental use of data when the valid signal was not
   // asserted. without this, the output of the register file would
   // "auto-update" based on new writes to the ram, a spooky behavior
   // that would never correspond to that of a hardened ram.
   
   //the read logic, register the input
   logic [addr_width_lp-1:0]  r0_addr_r, r1_addr_r;

   always_ff @(posedge clk_i)
     if (r0_v_i)
       r0_addr_r <= r0_addr_i;
     else
       r0_addr_r <= 'X;

   always_ff @(posedge clk_i)
     if (r1_v_i)
       r1_addr_r <= r1_addr_i;
     else
       r1_addr_r <= 'X;

   assign r0_data_o = mem[ r0_addr_r ];
   assign r1_data_o = mem[ r1_addr_r ];

   //the write logic, the memory is treated as dff array
   always_ff @(posedge clk_i)
     if (w_v_i)
       mem[w_addr_i] <= w_data_i;

   end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_2r1w_sync_synth)
// MBT 4/1/2014
//
// 2 read-port, 1 write-port ram
//
// reads are asynchronous
//
// this file should not be directly instantiated by end programmers
// use bsg_mem_2r1w instead
//

//`include "bsg_defines.sv"

module bsg_mem_2r1w_synth #(parameter `BSG_INV_PARAM(width_p)
			    , parameter `BSG_INV_PARAM(els_p)
			    , parameter read_write_same_addr_p=0
			    , parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
			    )
   (input   w_clk_i
    , input w_reset_i

    , input                     w_v_i
    , input [addr_width_lp-1:0] w_addr_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0]       w_data_i

    , input                      r0_v_i
    , input [addr_width_lp-1:0]  r0_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r0_data_o

    , input                      r1_v_i
    , input [addr_width_lp-1:0]  r1_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r1_data_o

    );

   wire                   unused = w_reset_i;

   if (width_p == 0 || els_p == 0)
    begin: z
      wire unused0 = &{w_clk_i, w_v_i, w_addr_i, w_data_i, r0_v_i, r0_addr_i, r1_v_i, r1_addr_i};
      assign r0_data_o = '0;
      assign r1_data_o = '0;
    end
   else
    begin: nz

   logic [width_p-1:0]    mem [els_p-1:0];

   // this implementation ignores the r_v_i
   wire [addr_width_lp-1:0]  r0_addr_li = (els_p>1) ? r0_addr_i:'0;
   wire [addr_width_lp-1:0]  r1_addr_li = (els_p>1) ? r1_addr_i:'0;

   assign r1_data_o = mem[r1_addr_li];
   assign r0_data_o = mem[r0_addr_li];
   
   wire [addr_width_lp-1:0]  w_addr_li = (els_p>1) ? w_addr_i:'0;

   always_ff @(posedge w_clk_i)
     if (w_v_i)
       begin
          mem[w_addr_li] <= w_data_i;
       end
   end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_2r1w_synth)

//`include "bsg_defines.sv"

module bsg_mem_2rw_sync_mask_write_bit_synth #( parameter `BSG_INV_PARAM(width_p )
                         , parameter `BSG_INV_PARAM(els_p )
                         , parameter read_write_same_addr_p = 0
                         , parameter disable_collision_warning_p = 0
                         , parameter addr_width_lp = `BSG_SAFE_CLOG2(els_p)
                         , parameter harden_p = 1
                         )
  ( input                      clk_i
  , input                      reset_i

  , input [width_p-1:0]        a_data_i
  , input [width_p-1:0]        a_w_mask_i
  , input [addr_width_lp-1:0]  a_addr_i
  , input                      a_v_i
  , input                      a_w_i

  , input [width_p-1:0]        b_data_i
  , input [width_p-1:0]        b_w_mask_i
  , input [addr_width_lp-1:0]  b_addr_i
  , input                      b_v_i
  , input                      b_w_i

  , output logic [width_p-1:0] a_data_o
  , output logic [width_p-1:0] b_data_o
  );

   wire                   unused = reset_i;

   if (width_p == 0)
    begin: z
      wire unused0 = &{clk_i, a_data_i, a_w_mask_i, a_addr_i, a_v_i, a_w_i};
      wire unused1 = &{clk_i, b_data_i, b_w_mask_i, b_addr_i, b_v_i, b_w_i};
      assign a_data_o = '0;
      assign b_data_o = '0;
    end
   else
    begin: nz

   logic [width_p-1:0]    mem [els_p-1:0];

   // this treats the ram as an array of registers for which the
   // read addr is latched on the clock, the write
   // is done on the clock edge, and actually multiplexing
   // of the registers for reading is done after the clock edge.

   // logically, this means that reads happen in time after
   // the writes, and "simultaneous" reads and writes to the
   // register file are allowed -- IF read_write_same_addr is set.

   // note that this behavior is generally incompatible with
   // hardened 1r1w rams, so it's better not to take advantage
   // of it if not necessary

   // we explicitly 'X out the read address if valid is not set
   // to avoid accidental use of data when the valid signal was not
   // asserted. without this, the output of the register file would
   // "auto-update" based on new writes to the ram, a spooky behavior
   // that would never correspond to that of a hardened ram.

   logic [addr_width_lp-1:0] a_addr_r, b_addr_r;

   always_ff @(posedge clk_i)
     begin
        if (a_v_i)
            a_addr_r <= a_addr_i;
        else
            a_addr_r <= 'X;
          
        if (b_v_i)
            b_addr_r <= b_addr_i;
        else
            b_addr_r <= 'X;

`ifndef BSG_HIDE_FROM_SYNTHESIS
        // if addresses match and this is forbidden, then nuke the read address

        if (a_addr_i == b_addr_i && a_v_i && b_v_i && (a_w_i || b_w_i) && !read_write_same_addr_p)
          begin
             if (!disable_collision_warning_p)
               begin
                 $error("X'ing matched read addresses %x %x (%m)",a_addr_i, b_addr_i);
               end
             a_addr_r <= 'X;
             b_addr_r <= 'X;
          end
`endif

     end

   assign a_data_o = mem[a_addr_r];
   assign b_data_o = mem[b_addr_r];


   genvar                       i;
   for (i = 0; i < width_p; i=i+1)
     begin
	always_ff @(posedge clk_i)
      begin

	  if (a_v_i & a_w_i && a_w_mask_i[i])
            mem[a_addr_i][i] <= a_data_i[i];
	  if (b_v_i & b_w_i && b_w_mask_i[i])
            mem[b_addr_i][i] <= b_data_i[i];
      end
     end
  end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_2rw_sync_mask_write_bit_synth)

//`include "bsg_defines.sv"

module bsg_mem_2rw_sync_mask_write_byte_synth #( parameter `BSG_INV_PARAM(width_p )
                         , parameter `BSG_INV_PARAM(els_p )
                         , parameter read_write_same_addr_p=0
                         , parameter addr_width_lp = `BSG_SAFE_CLOG2(els_p)
                         , parameter harden_p = 1
                         , parameter disable_collision_warning_p=0     
                         , parameter write_mask_width_lp=(width_p>>3)              
                         )
  ( input                      clk_i
  , input                      reset_i

  , input [width_p-1:0]        a_data_i
  , input [write_mask_width_lp-1:0] a_w_mask_i
  , input [addr_width_lp-1:0]  a_addr_i
  , input                      a_v_i
  , input                      a_w_i

  , input [width_p-1:0]        b_data_i
  , input [write_mask_width_lp-1:0] b_w_mask_i
  , input [addr_width_lp-1:0]  b_addr_i
  , input                      b_v_i
  , input                      b_w_i

  , output logic [width_p-1:0] a_data_o
  , output logic [width_p-1:0] b_data_o
  );

   wire                   unused = reset_i;

   if (width_p == 0)
    begin: z
      wire unused0 = &{clk_i, a_data_i, a_w_mask_i, a_addr_i, a_v_i, a_w_i};
      wire unused1 = &{clk_i, b_data_i, b_w_mask_i, b_addr_i, b_v_i, b_w_i};
      assign a_data_o = '0;
      assign b_data_o = '0;
    end
   else
    begin: nz

  genvar i;
  for(i=0; i<write_mask_width_lp; i=i+1)
  begin: bk
    bsg_mem_2rw_sync #( .width_p      (8)
                        ,.els_p        (els_p)
                        ,.addr_width_lp(addr_width_lp)
                        ,.disable_collision_warning_p(disable_collision_warning_p)
                        ,.harden_p(harden_p)
                      ) mem_2rw_sync
                      ( .clk_i  (clk_i)
                       ,.reset_i(reset_i)
                       ,.a_data_i (a_data_i[(i*8)+:8])
                       ,.a_addr_i (a_addr_i)
                       ,.a_v_i    (a_v_i & (a_w_i ? a_w_mask_i[i] : 1'b1))
                       ,.a_w_i    (a_w_i & a_w_mask_i[i])
                       ,.a_data_o (a_data_o[(i*8)+:8])
                       ,.b_data_i (b_data_i[(i*8)+:8])
                       ,.b_addr_i (b_addr_i)
                       ,.b_v_i    (b_v_i & (b_w_i ? b_w_mask_i[i] : 1'b1))
                       ,.b_w_i    (b_w_i & b_w_mask_i[i])
                       ,.b_data_o (b_data_o[(i*8)+:8])
                      );
  end
    end

endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_2rw_sync_mask_write_byte_synth)


//`include "bsg_defines.sv"

module bsg_mem_2rw_sync_synth #( parameter `BSG_INV_PARAM(width_p )
                         , parameter `BSG_INV_PARAM(els_p )
                         , parameter read_write_same_addr_p=0
                         , parameter addr_width_lp = `BSG_SAFE_CLOG2(els_p)
                         , parameter harden_p = 1
                         , parameter disable_collision_warning_p=0                   
                         )
  ( input                      clk_i
  , input                      reset_i

  , input [width_p-1:0]        a_data_i
  , input [addr_width_lp-1:0]  a_addr_i
  , input                      a_v_i
  , input                      a_w_i

  , input [width_p-1:0]        b_data_i
  , input [addr_width_lp-1:0]  b_addr_i
  , input                      b_v_i
  , input                      b_w_i

  , output logic [width_p-1:0] a_data_o
  , output logic [width_p-1:0] b_data_o
  );

   wire                   unused = reset_i;

   if (width_p == 0)
    begin: z
      wire unused0 = &{clk_i, a_data_i, a_addr_i, a_v_i, a_w_i};
      wire unused1 = &{clk_i, b_data_i, b_addr_i, b_v_i, b_w_i};
      assign a_data_o = '0;
      assign b_data_o = '0;
    end
   else
    begin: nz

   logic [width_p-1:0]    mem [els_p-1:0];

   // this treats the ram as an array of registers for which the
   // read addr is latched on the clock, the write
   // is done on the clock edge, and actually multiplexing
   // of the registers for reading is done after the clock edge.

   // logically, this means that reads happen in time after
   // the writes, and "simultaneous" reads and writes to the
   // register file are allowed -- IF read_write_same_addr is set.

   // note that this behavior is generally incompatible with
   // hardened 1r1w rams, so it's better not to take advantage
   // of it if not necessary

   // we explicitly 'X out the read address if valid is not set
   // to avoid accidental use of data when the valid signal was not
   // asserted. without this, the output of the register file would
   // "auto-update" based on new writes to the ram, a spooky behavior
   // that would never correspond to that of a hardened ram.

   logic [addr_width_lp-1:0] a_addr_r, b_addr_r;

   always_ff @(posedge clk_i)
     begin
        if (a_v_i)
            a_addr_r <= a_addr_i;
        else
            a_addr_r <= 'X;
          
        if (b_v_i)
            b_addr_r <= b_addr_i;
        else
            b_addr_r <= 'X;

`ifndef BSG_HIDE_FROM_SYNTHESIS
        // if addresses match and this is forbidden, then nuke the read address

        if (a_addr_i == b_addr_i && a_v_i && b_v_i && (a_w_i || b_w_i) && !read_write_same_addr_p)
          begin
             if (!disable_collision_warning_p)
               begin
                 $error("X'ing matched read address %x (%m)",a_addr_i);
               end
             a_addr_r <= 'X;
             b_addr_r <= 'X;
          end
`endif

     end

   assign a_data_o = mem[a_addr_r];
   assign b_data_o = mem[b_addr_r];

	always_ff @(posedge clk_i)
    begin
	  if (a_v_i & a_w_i)
            mem[a_addr_i] <= a_data_i;
	  if (b_v_i & b_w_i)
            mem[b_addr_i] <= b_data_i;
    end
  end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_2rw_sync_synth)

// MBT 7/7/2016
// DWP 11/27/2019
//
// 3 read-port, 1 write-port ram
//
// reads are synchronous
//
// although we could merge this with normal bsg_mem_1r1w
// and select with a parameter, we do not do this because
// it's typically a very big change to the instantiating code
// to move to/from sync/async, and we want to reflect this.
//
// NOTE: Users of BaseJump STL should not instantiate this module directly
// they should use bsg_mem_3r1w_sync.

//`include "bsg_defines.sv"

module bsg_mem_3r1w_sync_synth #(parameter `BSG_INV_PARAM(width_p)
				 , parameter `BSG_INV_PARAM(els_p)
				 , parameter read_write_same_addr_p=0
				 , parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
				 )
   (input   clk_i
    , input reset_i

    , input                     w_v_i
    , input [addr_width_lp-1:0] w_addr_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0]       w_data_i

    // currently unused
    , input                      r0_v_i
    , input [addr_width_lp-1:0]  r0_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r0_data_o

    , input                      r1_v_i
    , input [addr_width_lp-1:0]  r1_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r1_data_o

    , input                      r2_v_i
    , input [addr_width_lp-1:0]  r2_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r2_data_o
    );

   wire                   unused = reset_i;

   if (width_p == 0)
    begin: z
      wire unused0 = &{clk_i, w_v_i, w_addr_i, w_data_i, r0_v_i, r0_addr_i, r1_v_i, r1_addr_i, r2_v_i, r2_addr_i};
      assign r0_data_o = '0;
      assign r1_data_o = '0;
      assign r2_data_o = '0;
    end
   else
    begin: nz

   logic [width_p-1:0]    mem [els_p-1:0];

   // keep consistent with bsg_ip_cores/bsg_mem/bsg_mem_3r1w_sync.sv
   // keep consistent with bsg_ip_cores/hard/bsg_mem/bsg_mem_3r1w_sync.sv

   // this treats the ram as an array of registers for which the
   // read addr is latched on the clock, the write
   // is done on the clock edge, and actually multiplexing
   // of the registers for reading is done after the clock edge.

   // logically, this means that reads happen in time after
   // the writes, and "simultaneous" reads and writes to the
   // register file are allowed -- IF read_write_same_addr is set.

   // note that this behavior is generally incompatible with
   // hardened 1r1w rams, so it's better not to take advantage
   // of it if not necessary

   // we explicitly 'X out the read address if valid is not set
   // to avoid accidental use of data when the valid signal was not
   // asserted. without this, the output of the register file would
   // "auto-update" based on new writes to the ram, a spooky behavior
   // that would never correspond to that of a hardened ram.

   //the read logic, register the input
   logic [addr_width_lp-1:0]  r0_addr_r, r1_addr_r, r2_addr_r;

   always_ff @(posedge clk_i)
     if (r0_v_i)
       r0_addr_r <= r0_addr_i;
     else
       r0_addr_r <= 'X;

   always_ff @(posedge clk_i)
     if (r1_v_i)
       r1_addr_r <= r1_addr_i;
     else
       r1_addr_r <= 'X;

   always_ff @(posedge clk_i)
     if (r2_v_i)
       r2_addr_r <= r2_addr_i;
     else
       r2_addr_r <= 'X;

   assign r0_data_o = mem[ r0_addr_r ];
   assign r1_data_o = mem[ r1_addr_r ];
   assign r2_data_o = mem[ r2_addr_r ];

   //the write logic, the memory is treated as dff array
   always_ff @(posedge clk_i)
     if (w_v_i)
       mem[w_addr_i] <= w_data_i;

    end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_3r1w_sync_synth)
// MBT 4/1/2014
// DWP 11/27/2019
//
// 3 read-port, 1 write-port ram
//
// reads are asynchronous
//
// this file should not be directly instantiated by end programmers
// use bsg_mem_3r1w instead
//

//`include "bsg_defines.sv"

module bsg_mem_3r1w_synth #(parameter `BSG_INV_PARAM(width_p)
			    , parameter `BSG_INV_PARAM(els_p)
			    , parameter read_write_same_addr_p=0
			    , parameter addr_width_lp=`BSG_SAFE_CLOG2(els_p)
			    )
   (input   w_clk_i
    , input w_reset_i

    , input                     w_v_i
    , input [addr_width_lp-1:0] w_addr_i
    , input [`BSG_SAFE_MINUS(width_p, 1):0]       w_data_i

    , input                      r0_v_i
    , input [addr_width_lp-1:0]  r0_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r0_data_o

    , input                      r1_v_i
    , input [addr_width_lp-1:0]  r1_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r1_data_o

    , input                      r2_v_i
    , input [addr_width_lp-1:0]  r2_addr_i
    , output logic [`BSG_SAFE_MINUS(width_p, 1):0] r2_data_o
    );

   wire                   unused = w_reset_i;

   if (width_p == 0)
    begin: z
      wire unused0 = &{w_clk_i, w_v_i, w_addr_i, w_data_i, r0_v_i, r0_addr_i, r1_v_i, r1_addr_i, r2_v_i, r2_addr_i};
      assign r0_data_o = '0;
      assign r1_data_o = '0;
      assign r2_data_o = '0;
    end
   else
    begin: nz

   logic [width_p-1:0]    mem [els_p-1:0];

   // this implementation ignores the r_v_i
   assign r2_data_o = mem[r2_addr_i];
   assign r1_data_o = mem[r1_addr_i];
   assign r0_data_o = mem[r0_addr_i];

   wire                   unused = w_reset_i;

   always_ff @(posedge w_clk_i)
     if (w_v_i)
       begin
          mem[w_addr_i] <= w_data_i;
       end
    end
endmodule

//`BSG_ABSTRACT_MODULE(bsg_mem_3r1w_synth)


module bp_be_dcache_decoder_00_00000ffe
(
  pkt_i,
  decode_o
);

  input [22:0] pkt_i;
  output [32:0] decode_o;
  wire [32:0] decode_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,decode_o_4_,decode_o_3_,
  decode_o_2_,decode_o_1_,decode_o_0_,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,
  N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,
  N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
  N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,
  N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,
  N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,
  N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,
  N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,
  N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,
  N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,
  N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,
  N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,
  N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,
  N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,
  N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,
  N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,
  N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,
  N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,
  N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,
  N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,
  N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,
  N362,N363,N364,N365,N366,N367,N368,N369,N371,N372,N373,N374,N375,N376,N377,N378,
  N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,
  N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,
  N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,
  N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,
  N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458;
  assign decode_o[17] = 1'b0;
  assign decode_o_4_ = pkt_i[22];
  assign decode_o[4] = decode_o_4_;
  assign decode_o_3_ = pkt_i[21];
  assign decode_o[3] = decode_o_3_;
  assign decode_o_2_ = pkt_i[20];
  assign decode_o[2] = decode_o_2_;
  assign decode_o_1_ = pkt_i[19];
  assign decode_o[1] = decode_o_1_;
  assign decode_o_0_ = pkt_i[18];
  assign decode_o[0] = decode_o_0_;
  assign N14 = N26 | N342;
  assign N15 = N105 | N14;
  assign N16 = ~N15;
  assign N17 = N105 | N23;
  assign N18 = ~N17;
  assign decode_o[16] = N16 | N18;
  assign N19 = ~pkt_i[14];
  assign N20 = pkt_i[16] | pkt_i[17];
  assign N21 = N255 | N20;
  assign N22 = N19 | N21;
  assign N23 = pkt_i[13] | N22;
  assign N24 = pkt_i[12] | N23;
  assign N25 = ~N24;
  assign N26 = ~pkt_i[13];
  assign N27 = N26 | N22;
  assign N28 = pkt_i[12] | N27;
  assign N29 = ~N28;
  assign decode_o[15] = N25 | N29;
  assign N30 = pkt_i[17] | pkt_i[16];
  assign N31 = N26 | N105;
  assign N32 = N30 | N278;
  assign N33 = N32 | N31;
  assign N34 = N30 | N261;
  assign N35 = N34 | N262;
  assign N37 = N34 | N273;
  assign N38 = N34 | N265;
  assign N40 = pkt_i[17] | N99;
  assign N41 = N40 | N272;
  assign N42 = N41 | N273;
  assign N43 = N255 | pkt_i[14];
  assign N44 = N40 | N43;
  assign N45 = N44 | N262;
  assign N47 = N41 | N262;
  assign N48 = N44 | N265;
  assign N50 = N41 | N265;
  assign N51 = N44 | N31;
  assign N53 = N41 | N31;
  assign N54 = N40 | N261;
  assign N55 = N54 | N273;
  assign N57 = N40 | N278;
  assign N58 = N57 | N273;
  assign N59 = N54 | N262;
  assign N61 = N57 | N262;
  assign N62 = N54 | N265;
  assign N64 = N57 | N265;
  assign N65 = N54 | N31;
  assign N67 = N57 | N31;
  assign N68 = N98 | pkt_i[16];
  assign N69 = N68 | N272;
  assign N70 = N69 | N273;
  assign N72 = N44 | N273;
  assign N73 = N69 | N262;
  assign N75 = N305 & N268;
  assign N76 = N99 & N255;
  assign N77 = N76 & N314;
  assign N78 = pkt_i[17] & pkt_i[13];
  assign N79 = pkt_i[13] & N105;
  assign N80 = N76 & N79;
  assign N81 = N329 & pkt_i[13];
  assign N82 = pkt_i[17] & pkt_i[14];
  assign N83 = pkt_i[14] & N105;
  assign N84 = N76 & N83;
  assign N85 = N305 & N19;
  assign N86 = N98 & N99;
  assign N87 = N86 & N19;
  assign N89 = N26 | N102;
  assign N90 = pkt_i[12] | N89;
  assign N91 = ~N90;
  assign decode_o[10] = N91 | N97;
  assign N92 = N105 | N103;
  assign N93 = ~N92;
  assign N94 = N19 | N101;
  assign N95 = pkt_i[13] | N94;
  assign N96 = pkt_i[12] | N95;
  assign N97 = ~N96;
  assign decode_o[11] = N93 | N97;
  assign N98 = ~pkt_i[17];
  assign N99 = ~pkt_i[16];
  assign N100 = N99 | N98;
  assign N101 = pkt_i[15] | N100;
  assign N102 = pkt_i[14] | N101;
  assign N103 = pkt_i[13] | N102;
  assign N104 = pkt_i[12] | N103;
  assign decode_o[9] = ~N104;
  assign N105 = ~pkt_i[12];
  assign N106 = pkt_i[13] | N109;
  assign N107 = N105 | N106;
  assign N108 = ~N107;
  assign decode_o[12] = N108 | N117;
  assign N109 = N19 | N256;
  assign N110 = N26 | N109;
  assign N111 = pkt_i[12] | N110;
  assign N112 = ~N111;
  assign N113 = pkt_i[16] & pkt_i[17];
  assign N114 = pkt_i[15] & N113;
  assign N115 = pkt_i[14] & N114;
  assign N116 = pkt_i[13] & N115;
  assign N117 = pkt_i[12] & N116;
  assign decode_o[13] = N112 | N117;
  assign N118 = N105 | N121;
  assign N119 = ~N118;
  assign N120 = N253 | N119;
  assign N121 = N26 | N128;
  assign N122 = pkt_i[12] | N121;
  assign N123 = ~N122;
  assign N124 = N120 | N123;
  assign N125 = N105 | N129;
  assign N126 = ~N125;
  assign N127 = N124 | N126;
  assign N128 = pkt_i[14] | N341;
  assign N129 = pkt_i[13] | N128;
  assign N130 = pkt_i[12] | N129;
  assign N131 = ~N130;
  assign N132 = N127 | N131;
  assign N133 = N132 | N337;
  assign N134 = N133 | N339;
  assign N135 = N134 | N345;
  assign N136 = ~N259;
  assign N137 = N135 | N136;
  assign N138 = N26 | N147;
  assign N139 = N105 | N138;
  assign N140 = ~N139;
  assign N141 = pkt_i[12] | N138;
  assign N142 = ~N141;
  assign N143 = N140 | N142;
  assign N144 = N105 | N148;
  assign N145 = ~N144;
  assign N146 = N143 | N145;
  assign N147 = pkt_i[14] | N21;
  assign N148 = pkt_i[13] | N147;
  assign N149 = pkt_i[12] | N148;
  assign N150 = ~N149;
  assign N151 = N146 | N150;
  assign N152 = pkt_i[12] | N158;
  assign N153 = ~N152;
  assign N154 = N151 | N153;
  assign N155 = pkt_i[16] | N98;
  assign N156 = pkt_i[15] | N155;
  assign N157 = N19 | N156;
  assign N158 = pkt_i[13] | N157;
  assign N159 = N105 | N158;
  assign N160 = ~N159;
  assign N161 = N154 | N160;
  assign N162 = ~N104;
  assign N163 = N161 | N162;
  assign N164 = N131 | N126;
  assign N165 = N164 | N123;
  assign N166 = N165 | N119;
  assign N167 = N166 | N345;
  assign N168 = N167 | N339;
  assign N169 = N168 | N337;
  assign N170 = N169 | N150;
  assign N171 = N170 | N145;
  assign N172 = N171 | N142;
  assign N173 = N172 | N140;
  assign N174 = N173 | N16;
  assign N175 = N174 | N25;
  assign N176 = N175 | N18;
  assign N177 = N176 | N29;
  assign N178 = pkt_i[12] | N181;
  assign N179 = ~N178;
  assign N180 = N177 | N179;
  assign N181 = pkt_i[13] | N188;
  assign N182 = N105 | N181;
  assign N183 = ~N182;
  assign N184 = N180 | N183;
  assign N185 = pkt_i[12] | N189;
  assign N186 = ~N185;
  assign N187 = N184 | N186;
  assign N188 = pkt_i[14] | N203;
  assign N189 = N26 | N188;
  assign N190 = N105 | N189;
  assign N191 = ~N190;
  assign N192 = N187 | N191;
  assign N193 = pkt_i[12] | N196;
  assign N194 = ~N193;
  assign N195 = N192 | N194;
  assign N196 = pkt_i[13] | N204;
  assign N197 = N105 | N196;
  assign N198 = ~N197;
  assign N199 = N195 | N198;
  assign N200 = pkt_i[12] | N205;
  assign N201 = ~N200;
  assign N202 = N199 | N201;
  assign N203 = pkt_i[15] | N234;
  assign N204 = N19 | N203;
  assign N205 = N26 | N204;
  assign N206 = N105 | N205;
  assign N207 = ~N206;
  assign N208 = N202 | N207;
  assign N209 = pkt_i[12] | N212;
  assign N210 = ~N209;
  assign N211 = N208 | N210;
  assign N212 = pkt_i[13] | N219;
  assign N213 = N105 | N212;
  assign N214 = ~N213;
  assign N215 = N211 | N214;
  assign N216 = pkt_i[12] | N220;
  assign N217 = ~N216;
  assign N218 = N215 | N217;
  assign N219 = pkt_i[14] | N235;
  assign N220 = N26 | N219;
  assign N221 = N105 | N220;
  assign N222 = ~N221;
  assign N223 = N218 | N222;
  assign N224 = pkt_i[12] | N227;
  assign N225 = ~N224;
  assign N226 = N223 | N225;
  assign N227 = pkt_i[13] | N236;
  assign N228 = N105 | N227;
  assign N229 = ~N228;
  assign N230 = N226 | N229;
  assign N231 = pkt_i[12] | N237;
  assign N232 = ~N231;
  assign N233 = N230 | N232;
  assign N234 = N99 | pkt_i[17];
  assign N235 = N255 | N234;
  assign N236 = N19 | N235;
  assign N237 = N26 | N236;
  assign N238 = N105 | N237;
  assign N239 = ~N238;
  assign N240 = N233 | N239;
  assign N241 = pkt_i[12] | N244;
  assign N242 = ~N241;
  assign N243 = N240 | N242;
  assign N244 = pkt_i[13] | N247;
  assign N245 = N105 | N244;
  assign N246 = ~N245;
  assign decode_o[25] = N243 | N246;
  assign N247 = pkt_i[14] | N156;
  assign N248 = N26 | N247;
  assign N249 = pkt_i[12] | N248;
  assign N250 = ~N249;
  assign N251 = N105 | N248;
  assign N252 = ~N251;
  assign N253 = N250 | N252;
  assign N254 = N253 | N153;
  assign decode_o[26] = N254 | N160;
  assign N255 = ~pkt_i[15];
  assign N256 = N255 | N100;
  assign N257 = pkt_i[14] | N256;
  assign N258 = pkt_i[13] | N257;
  assign N259 = pkt_i[12] | N258;
  assign decode_o[24] = ~N259;
  assign N260 = N98 | N99;
  assign N261 = N255 | N19;
  assign N262 = pkt_i[13] | N105;
  assign N263 = N260 | N261;
  assign N264 = N263 | N262;
  assign N265 = N26 | pkt_i[12];
  assign N266 = N263 | N265;
  assign N267 = pkt_i[17] & pkt_i[16];
  assign N268 = pkt_i[13] & pkt_i[12];
  assign N269 = N267 & N310;
  assign N270 = N269 & N268;
  assign N272 = pkt_i[15] | pkt_i[14];
  assign N273 = pkt_i[13] | pkt_i[12];
  assign N274 = N260 | N272;
  assign N275 = N274 | N273;
  assign N276 = N274 | N265;
  assign N277 = N274 | N262;
  assign N278 = pkt_i[15] | N19;
  assign N279 = N260 | N278;
  assign N280 = N279 | N273;
  assign N282 = N255 & N19;
  assign N283 = N26 & N105;
  assign N284 = N86 & N282;
  assign N285 = N284 & N283;
  assign N286 = N32 | N273;
  assign N287 = N296 | N273;
  assign N289 = N293 | N262;
  assign N290 = N32 | N262;
  assign N291 = N296 | N262;
  assign N293 = N30 | N272;
  assign N294 = N293 | N265;
  assign N295 = N32 | N265;
  assign N296 = N30 | N43;
  assign N297 = N296 | N265;
  assign N298 = N69 | N265;
  assign N299 = N68 | N278;
  assign N300 = N299 | N273;
  assign N302 = N98 & pkt_i[15];
  assign N303 = pkt_i[14] & pkt_i[12];
  assign N304 = N302 & N303;
  assign N305 = N99 & pkt_i[15];
  assign N306 = N305 & N303;
  assign N307 = pkt_i[17] & N255;
  assign N308 = N307 & N303;
  assign N309 = N98 & pkt_i[16];
  assign N310 = pkt_i[15] & pkt_i[14];
  assign N311 = N309 & N310;
  assign N312 = pkt_i[14] & pkt_i[13];
  assign N313 = N307 & N312;
  assign N314 = pkt_i[14] & N26;
  assign N315 = N322 & N314;
  assign N316 = N315 & N105;
  assign N317 = N320 & N312;
  assign N318 = N317 & N105;
  assign N319 = N305 & N312;
  assign N320 = pkt_i[17] & N99;
  assign N321 = N320 & pkt_i[15];
  assign N322 = pkt_i[16] & pkt_i[15];
  assign N323 = N19 & pkt_i[12];
  assign N324 = N322 & N323;
  assign N325 = pkt_i[17] & N19;
  assign N326 = N325 & N268;
  assign N327 = N19 & pkt_i[13];
  assign N328 = N322 & N327;
  assign N329 = N99 & N19;
  assign N330 = N329 & N268;
  assign N331 = pkt_i[17] & pkt_i[15];
  assign N332 = N331 & N19;
  assign N333 = N19 & N26;
  assign N334 = N320 & N333;
  assign N336 = pkt_i[12] | N14;
  assign N337 = ~N336;
  assign N338 = N105 | N343;
  assign N339 = ~N338;
  assign N340 = N337 | N339;
  assign N341 = pkt_i[15] | N20;
  assign N342 = N19 | N341;
  assign N343 = pkt_i[13] | N342;
  assign N344 = pkt_i[12] | N343;
  assign N345 = ~N344;
  assign N346 = N340 | N345;
  assign N364 = decode_o_3_ | decode_o_4_;
  assign N365 = decode_o_2_ | N364;
  assign N366 = decode_o_1_ | N365;
  assign N367 = decode_o_0_ | N366;
  assign N368 = decode_o[7] | decode_o[8];
  assign N369 = decode_o[6] | N368;
  assign decode_o[14] = decode_o[5] | N369;
  assign decode_o[8:5] = (N0)? { 1'b0, 1'b0, 1'b0, 1'b1 } : 
                         (N1)? { 1'b0, 1'b0, 1'b1, 1'b0 } : 
                         (N2)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                         (N3)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                         (N4)? { 1'b0, 1'b1, 1'b0, 1'b1 } : 
                         (N5)? { 1'b0, 1'b1, 1'b1, 1'b0 } : 
                         (N6)? { 1'b0, 1'b1, 1'b1, 1'b1 } : 
                         (N7)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                         (N8)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                         (N9)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                         (N10)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                         (N11)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N36;
  assign N1 = N39;
  assign N2 = N46;
  assign N3 = N49;
  assign N4 = N52;
  assign N5 = N56;
  assign N6 = N60;
  assign N7 = N63;
  assign N8 = N66;
  assign N9 = N71;
  assign N10 = N74;
  assign N11 = N88;
  assign decode_o[31] = (N12)? 1'b1 : 
                        (N357)? 1'b0 : 
                        (N360)? 1'b1 : 
                        (N363)? 1'b1 : 
                        (N354)? 1'b0 : 1'b0;
  assign N12 = N347;
  assign decode_o[32] = (N12)? 1'b1 : 
                        (N357)? 1'b1 : 
                        (N355)? 1'b0 : 
                        (N13)? 1'b0 : 
                        (N13)? 1'b0 : 1'b0;
  assign N13 = 1'b0;
  assign N36 = N371 | N372;
  assign N371 = ~N33;
  assign N372 = ~N35;
  assign N39 = N373 | N374;
  assign N373 = ~N37;
  assign N374 = ~N38;
  assign N46 = N375 | N376;
  assign N375 = ~N42;
  assign N376 = ~N45;
  assign N49 = N377 | N378;
  assign N377 = ~N47;
  assign N378 = ~N48;
  assign N52 = N379 | N380;
  assign N379 = ~N50;
  assign N380 = ~N51;
  assign N56 = N381 | N382;
  assign N381 = ~N53;
  assign N382 = ~N55;
  assign N60 = N383 | N384;
  assign N383 = ~N58;
  assign N384 = ~N59;
  assign N63 = N385 | N386;
  assign N385 = ~N61;
  assign N386 = ~N62;
  assign N66 = N387 | N388;
  assign N387 = ~N64;
  assign N388 = ~N65;
  assign N71 = N389 | N390;
  assign N389 = ~N67;
  assign N390 = ~N70;
  assign N74 = N391 | N392;
  assign N391 = ~N72;
  assign N392 = ~N73;
  assign N88 = N75 | N401;
  assign N401 = N77 | N400;
  assign N400 = N78 | N399;
  assign N399 = N80 | N398;
  assign N398 = N81 | N397;
  assign N397 = N82 | N396;
  assign N396 = N84 | N395;
  assign N395 = N331 | N394;
  assign N394 = N85 | N393;
  assign N393 = N267 | N87;
  assign decode_o[30] = N402 | N137;
  assign N402 = decode_o[14] | decode_o[16];
  assign decode_o[28] = N404 | N163;
  assign N404 = decode_o[14] & N403;
  assign N403 = ~decode_o[16];
  assign N271 = N407 | N270;
  assign N407 = N405 | N406;
  assign N405 = ~N264;
  assign N406 = ~N266;
  assign N281 = N412 | N413;
  assign N412 = N410 | N411;
  assign N410 = N408 | N409;
  assign N408 = ~N275;
  assign N409 = ~N276;
  assign N411 = ~N277;
  assign N413 = ~N280;
  assign N288 = N415 | N416;
  assign N415 = N285 | N414;
  assign N414 = ~N286;
  assign N416 = ~N287;
  assign N292 = N419 | N420;
  assign N419 = N417 | N418;
  assign N417 = ~N289;
  assign N418 = ~N290;
  assign N420 = ~N291;
  assign N301 = N439 | N373;
  assign N439 = N438 | N371;
  assign N438 = N436 | N437;
  assign N436 = N434 | N435;
  assign N434 = N432 | N433;
  assign N432 = N430 | N431;
  assign N430 = N428 | N429;
  assign N428 = N427 | N391;
  assign N427 = N426 | N389;
  assign N426 = N425 | N387;
  assign N425 = N424 | N385;
  assign N424 = N423 | N383;
  assign N423 = N422 | N381;
  assign N422 = N421 | N379;
  assign N421 = N375 | N377;
  assign N429 = ~N294;
  assign N431 = ~N295;
  assign N433 = ~N297;
  assign N435 = ~N298;
  assign N437 = ~N300;
  assign N335 = N304 | N452;
  assign N452 = N306 | N451;
  assign N451 = N308 | N450;
  assign N450 = N311 | N449;
  assign N449 = N313 | N448;
  assign N448 = N316 | N447;
  assign N447 = N318 | N446;
  assign N446 = N319 | N445;
  assign N445 = N321 | N444;
  assign N444 = N324 | N443;
  assign N443 = N326 | N442;
  assign N442 = N328 | N441;
  assign N441 = N330 | N440;
  assign N440 = N332 | N334;
  assign decode_o[23] = N271;
  assign decode_o[22] = N281;
  assign decode_o[18] = N288;
  assign decode_o[19] = N292;
  assign decode_o[20] = N301;
  assign decode_o[21] = N335;
  assign decode_o[27] = N454 & N455;
  assign N454 = N453 | decode_o[20];
  assign N453 = decode_o[18] | decode_o[19];
  assign N455 = ~N346;
  assign N347 = decode_o[25] & decode_o[18];
  assign N348 = decode_o[25] & decode_o[19];
  assign N349 = decode_o[25] & decode_o[20];
  assign N350 = decode_o[26] & decode_o[20];
  assign N351 = N348 | N347;
  assign N352 = N349 | N351;
  assign N353 = N350 | N352;
  assign N354 = ~N353;
  assign N355 = ~N351;
  assign decode_o[29] = decode_o[30] & N458;
  assign N458 = N456 | N457;
  assign N456 = decode_o[24] | decode_o[26];
  assign N457 = decode_o[25] & N367;
  assign N356 = ~N347;
  assign N357 = N348 & N356;
  assign N358 = ~N348;
  assign N359 = N356 & N358;
  assign N360 = N349 & N359;
  assign N361 = ~N349;
  assign N362 = N359 & N361;
  assign N363 = N350 & N362;

endmodule



module bsg_mem_1rw_sync_mask_write_bit_000000b8_00000040_1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [183:0] data_i;
  input [5:0] addr_i;
  input [183:0] w_mask_i;
  output [183:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [183:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  addr_i,
  data_i,
  write_mask_i,
  data_o
);

  input [8:0] addr_i;
  input [63:0] data_i;
  input [7:0] write_mask_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [63:0] data_o;

  bsg_mem_1rw_sync_mask_write_byte_synth
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .w_i(w_i),
    .addr_i(addr_i),
    .data_i(data_i),
    .write_mask_i(write_mask_i),
    .data_o(data_o)
  );


endmodule



module bsg_dff_reset_width_p1
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  wire [0:0] data_o;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_width_p45
(
  clk_i,
  data_i,
  data_o
);

  input [44:0] data_i;
  output [44:0] data_o;
  input clk_i;
  wire [44:0] data_o;
  reg data_o_44_sv2v_reg,data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,
  data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,
  data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,
  data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,
  data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,
  data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,
  data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,
  data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_decode_00000008
(
  i,
  o
);

  input [2:0] i;
  output [7:0] o;
  wire [7:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_mux_000002aa_2
(
  data_i,
  sel_i,
  data_o
);

  input [1363:0] data_i;
  input [0:0] sel_i;
  output [681:0] data_o;
  wire [681:0] data_o;
  wire N0,N1;
  assign data_o[681] = (N1)? data_i[681] : 
                       (N0)? data_i[1363] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[680] = (N1)? data_i[680] : 
                       (N0)? data_i[1362] : 1'b0;
  assign data_o[679] = (N1)? data_i[679] : 
                       (N0)? data_i[1361] : 1'b0;
  assign data_o[678] = (N1)? data_i[678] : 
                       (N0)? data_i[1360] : 1'b0;
  assign data_o[677] = (N1)? data_i[677] : 
                       (N0)? data_i[1359] : 1'b0;
  assign data_o[676] = (N1)? data_i[676] : 
                       (N0)? data_i[1358] : 1'b0;
  assign data_o[675] = (N1)? data_i[675] : 
                       (N0)? data_i[1357] : 1'b0;
  assign data_o[674] = (N1)? data_i[674] : 
                       (N0)? data_i[1356] : 1'b0;
  assign data_o[673] = (N1)? data_i[673] : 
                       (N0)? data_i[1355] : 1'b0;
  assign data_o[672] = (N1)? data_i[672] : 
                       (N0)? data_i[1354] : 1'b0;
  assign data_o[671] = (N1)? data_i[671] : 
                       (N0)? data_i[1353] : 1'b0;
  assign data_o[670] = (N1)? data_i[670] : 
                       (N0)? data_i[1352] : 1'b0;
  assign data_o[669] = (N1)? data_i[669] : 
                       (N0)? data_i[1351] : 1'b0;
  assign data_o[668] = (N1)? data_i[668] : 
                       (N0)? data_i[1350] : 1'b0;
  assign data_o[667] = (N1)? data_i[667] : 
                       (N0)? data_i[1349] : 1'b0;
  assign data_o[666] = (N1)? data_i[666] : 
                       (N0)? data_i[1348] : 1'b0;
  assign data_o[665] = (N1)? data_i[665] : 
                       (N0)? data_i[1347] : 1'b0;
  assign data_o[664] = (N1)? data_i[664] : 
                       (N0)? data_i[1346] : 1'b0;
  assign data_o[663] = (N1)? data_i[663] : 
                       (N0)? data_i[1345] : 1'b0;
  assign data_o[662] = (N1)? data_i[662] : 
                       (N0)? data_i[1344] : 1'b0;
  assign data_o[661] = (N1)? data_i[661] : 
                       (N0)? data_i[1343] : 1'b0;
  assign data_o[660] = (N1)? data_i[660] : 
                       (N0)? data_i[1342] : 1'b0;
  assign data_o[659] = (N1)? data_i[659] : 
                       (N0)? data_i[1341] : 1'b0;
  assign data_o[658] = (N1)? data_i[658] : 
                       (N0)? data_i[1340] : 1'b0;
  assign data_o[657] = (N1)? data_i[657] : 
                       (N0)? data_i[1339] : 1'b0;
  assign data_o[656] = (N1)? data_i[656] : 
                       (N0)? data_i[1338] : 1'b0;
  assign data_o[655] = (N1)? data_i[655] : 
                       (N0)? data_i[1337] : 1'b0;
  assign data_o[654] = (N1)? data_i[654] : 
                       (N0)? data_i[1336] : 1'b0;
  assign data_o[653] = (N1)? data_i[653] : 
                       (N0)? data_i[1335] : 1'b0;
  assign data_o[652] = (N1)? data_i[652] : 
                       (N0)? data_i[1334] : 1'b0;
  assign data_o[651] = (N1)? data_i[651] : 
                       (N0)? data_i[1333] : 1'b0;
  assign data_o[650] = (N1)? data_i[650] : 
                       (N0)? data_i[1332] : 1'b0;
  assign data_o[649] = (N1)? data_i[649] : 
                       (N0)? data_i[1331] : 1'b0;
  assign data_o[648] = (N1)? data_i[648] : 
                       (N0)? data_i[1330] : 1'b0;
  assign data_o[647] = (N1)? data_i[647] : 
                       (N0)? data_i[1329] : 1'b0;
  assign data_o[646] = (N1)? data_i[646] : 
                       (N0)? data_i[1328] : 1'b0;
  assign data_o[645] = (N1)? data_i[645] : 
                       (N0)? data_i[1327] : 1'b0;
  assign data_o[644] = (N1)? data_i[644] : 
                       (N0)? data_i[1326] : 1'b0;
  assign data_o[643] = (N1)? data_i[643] : 
                       (N0)? data_i[1325] : 1'b0;
  assign data_o[642] = (N1)? data_i[642] : 
                       (N0)? data_i[1324] : 1'b0;
  assign data_o[641] = (N1)? data_i[641] : 
                       (N0)? data_i[1323] : 1'b0;
  assign data_o[640] = (N1)? data_i[640] : 
                       (N0)? data_i[1322] : 1'b0;
  assign data_o[639] = (N1)? data_i[639] : 
                       (N0)? data_i[1321] : 1'b0;
  assign data_o[638] = (N1)? data_i[638] : 
                       (N0)? data_i[1320] : 1'b0;
  assign data_o[637] = (N1)? data_i[637] : 
                       (N0)? data_i[1319] : 1'b0;
  assign data_o[636] = (N1)? data_i[636] : 
                       (N0)? data_i[1318] : 1'b0;
  assign data_o[635] = (N1)? data_i[635] : 
                       (N0)? data_i[1317] : 1'b0;
  assign data_o[634] = (N1)? data_i[634] : 
                       (N0)? data_i[1316] : 1'b0;
  assign data_o[633] = (N1)? data_i[633] : 
                       (N0)? data_i[1315] : 1'b0;
  assign data_o[632] = (N1)? data_i[632] : 
                       (N0)? data_i[1314] : 1'b0;
  assign data_o[631] = (N1)? data_i[631] : 
                       (N0)? data_i[1313] : 1'b0;
  assign data_o[630] = (N1)? data_i[630] : 
                       (N0)? data_i[1312] : 1'b0;
  assign data_o[629] = (N1)? data_i[629] : 
                       (N0)? data_i[1311] : 1'b0;
  assign data_o[628] = (N1)? data_i[628] : 
                       (N0)? data_i[1310] : 1'b0;
  assign data_o[627] = (N1)? data_i[627] : 
                       (N0)? data_i[1309] : 1'b0;
  assign data_o[626] = (N1)? data_i[626] : 
                       (N0)? data_i[1308] : 1'b0;
  assign data_o[625] = (N1)? data_i[625] : 
                       (N0)? data_i[1307] : 1'b0;
  assign data_o[624] = (N1)? data_i[624] : 
                       (N0)? data_i[1306] : 1'b0;
  assign data_o[623] = (N1)? data_i[623] : 
                       (N0)? data_i[1305] : 1'b0;
  assign data_o[622] = (N1)? data_i[622] : 
                       (N0)? data_i[1304] : 1'b0;
  assign data_o[621] = (N1)? data_i[621] : 
                       (N0)? data_i[1303] : 1'b0;
  assign data_o[620] = (N1)? data_i[620] : 
                       (N0)? data_i[1302] : 1'b0;
  assign data_o[619] = (N1)? data_i[619] : 
                       (N0)? data_i[1301] : 1'b0;
  assign data_o[618] = (N1)? data_i[618] : 
                       (N0)? data_i[1300] : 1'b0;
  assign data_o[617] = (N1)? data_i[617] : 
                       (N0)? data_i[1299] : 1'b0;
  assign data_o[616] = (N1)? data_i[616] : 
                       (N0)? data_i[1298] : 1'b0;
  assign data_o[615] = (N1)? data_i[615] : 
                       (N0)? data_i[1297] : 1'b0;
  assign data_o[614] = (N1)? data_i[614] : 
                       (N0)? data_i[1296] : 1'b0;
  assign data_o[613] = (N1)? data_i[613] : 
                       (N0)? data_i[1295] : 1'b0;
  assign data_o[612] = (N1)? data_i[612] : 
                       (N0)? data_i[1294] : 1'b0;
  assign data_o[611] = (N1)? data_i[611] : 
                       (N0)? data_i[1293] : 1'b0;
  assign data_o[610] = (N1)? data_i[610] : 
                       (N0)? data_i[1292] : 1'b0;
  assign data_o[609] = (N1)? data_i[609] : 
                       (N0)? data_i[1291] : 1'b0;
  assign data_o[608] = (N1)? data_i[608] : 
                       (N0)? data_i[1290] : 1'b0;
  assign data_o[607] = (N1)? data_i[607] : 
                       (N0)? data_i[1289] : 1'b0;
  assign data_o[606] = (N1)? data_i[606] : 
                       (N0)? data_i[1288] : 1'b0;
  assign data_o[605] = (N1)? data_i[605] : 
                       (N0)? data_i[1287] : 1'b0;
  assign data_o[604] = (N1)? data_i[604] : 
                       (N0)? data_i[1286] : 1'b0;
  assign data_o[603] = (N1)? data_i[603] : 
                       (N0)? data_i[1285] : 1'b0;
  assign data_o[602] = (N1)? data_i[602] : 
                       (N0)? data_i[1284] : 1'b0;
  assign data_o[601] = (N1)? data_i[601] : 
                       (N0)? data_i[1283] : 1'b0;
  assign data_o[600] = (N1)? data_i[600] : 
                       (N0)? data_i[1282] : 1'b0;
  assign data_o[599] = (N1)? data_i[599] : 
                       (N0)? data_i[1281] : 1'b0;
  assign data_o[598] = (N1)? data_i[598] : 
                       (N0)? data_i[1280] : 1'b0;
  assign data_o[597] = (N1)? data_i[597] : 
                       (N0)? data_i[1279] : 1'b0;
  assign data_o[596] = (N1)? data_i[596] : 
                       (N0)? data_i[1278] : 1'b0;
  assign data_o[595] = (N1)? data_i[595] : 
                       (N0)? data_i[1277] : 1'b0;
  assign data_o[594] = (N1)? data_i[594] : 
                       (N0)? data_i[1276] : 1'b0;
  assign data_o[593] = (N1)? data_i[593] : 
                       (N0)? data_i[1275] : 1'b0;
  assign data_o[592] = (N1)? data_i[592] : 
                       (N0)? data_i[1274] : 1'b0;
  assign data_o[591] = (N1)? data_i[591] : 
                       (N0)? data_i[1273] : 1'b0;
  assign data_o[590] = (N1)? data_i[590] : 
                       (N0)? data_i[1272] : 1'b0;
  assign data_o[589] = (N1)? data_i[589] : 
                       (N0)? data_i[1271] : 1'b0;
  assign data_o[588] = (N1)? data_i[588] : 
                       (N0)? data_i[1270] : 1'b0;
  assign data_o[587] = (N1)? data_i[587] : 
                       (N0)? data_i[1269] : 1'b0;
  assign data_o[586] = (N1)? data_i[586] : 
                       (N0)? data_i[1268] : 1'b0;
  assign data_o[585] = (N1)? data_i[585] : 
                       (N0)? data_i[1267] : 1'b0;
  assign data_o[584] = (N1)? data_i[584] : 
                       (N0)? data_i[1266] : 1'b0;
  assign data_o[583] = (N1)? data_i[583] : 
                       (N0)? data_i[1265] : 1'b0;
  assign data_o[582] = (N1)? data_i[582] : 
                       (N0)? data_i[1264] : 1'b0;
  assign data_o[581] = (N1)? data_i[581] : 
                       (N0)? data_i[1263] : 1'b0;
  assign data_o[580] = (N1)? data_i[580] : 
                       (N0)? data_i[1262] : 1'b0;
  assign data_o[579] = (N1)? data_i[579] : 
                       (N0)? data_i[1261] : 1'b0;
  assign data_o[578] = (N1)? data_i[578] : 
                       (N0)? data_i[1260] : 1'b0;
  assign data_o[577] = (N1)? data_i[577] : 
                       (N0)? data_i[1259] : 1'b0;
  assign data_o[576] = (N1)? data_i[576] : 
                       (N0)? data_i[1258] : 1'b0;
  assign data_o[575] = (N1)? data_i[575] : 
                       (N0)? data_i[1257] : 1'b0;
  assign data_o[574] = (N1)? data_i[574] : 
                       (N0)? data_i[1256] : 1'b0;
  assign data_o[573] = (N1)? data_i[573] : 
                       (N0)? data_i[1255] : 1'b0;
  assign data_o[572] = (N1)? data_i[572] : 
                       (N0)? data_i[1254] : 1'b0;
  assign data_o[571] = (N1)? data_i[571] : 
                       (N0)? data_i[1253] : 1'b0;
  assign data_o[570] = (N1)? data_i[570] : 
                       (N0)? data_i[1252] : 1'b0;
  assign data_o[569] = (N1)? data_i[569] : 
                       (N0)? data_i[1251] : 1'b0;
  assign data_o[568] = (N1)? data_i[568] : 
                       (N0)? data_i[1250] : 1'b0;
  assign data_o[567] = (N1)? data_i[567] : 
                       (N0)? data_i[1249] : 1'b0;
  assign data_o[566] = (N1)? data_i[566] : 
                       (N0)? data_i[1248] : 1'b0;
  assign data_o[565] = (N1)? data_i[565] : 
                       (N0)? data_i[1247] : 1'b0;
  assign data_o[564] = (N1)? data_i[564] : 
                       (N0)? data_i[1246] : 1'b0;
  assign data_o[563] = (N1)? data_i[563] : 
                       (N0)? data_i[1245] : 1'b0;
  assign data_o[562] = (N1)? data_i[562] : 
                       (N0)? data_i[1244] : 1'b0;
  assign data_o[561] = (N1)? data_i[561] : 
                       (N0)? data_i[1243] : 1'b0;
  assign data_o[560] = (N1)? data_i[560] : 
                       (N0)? data_i[1242] : 1'b0;
  assign data_o[559] = (N1)? data_i[559] : 
                       (N0)? data_i[1241] : 1'b0;
  assign data_o[558] = (N1)? data_i[558] : 
                       (N0)? data_i[1240] : 1'b0;
  assign data_o[557] = (N1)? data_i[557] : 
                       (N0)? data_i[1239] : 1'b0;
  assign data_o[556] = (N1)? data_i[556] : 
                       (N0)? data_i[1238] : 1'b0;
  assign data_o[555] = (N1)? data_i[555] : 
                       (N0)? data_i[1237] : 1'b0;
  assign data_o[554] = (N1)? data_i[554] : 
                       (N0)? data_i[1236] : 1'b0;
  assign data_o[553] = (N1)? data_i[553] : 
                       (N0)? data_i[1235] : 1'b0;
  assign data_o[552] = (N1)? data_i[552] : 
                       (N0)? data_i[1234] : 1'b0;
  assign data_o[551] = (N1)? data_i[551] : 
                       (N0)? data_i[1233] : 1'b0;
  assign data_o[550] = (N1)? data_i[550] : 
                       (N0)? data_i[1232] : 1'b0;
  assign data_o[549] = (N1)? data_i[549] : 
                       (N0)? data_i[1231] : 1'b0;
  assign data_o[548] = (N1)? data_i[548] : 
                       (N0)? data_i[1230] : 1'b0;
  assign data_o[547] = (N1)? data_i[547] : 
                       (N0)? data_i[1229] : 1'b0;
  assign data_o[546] = (N1)? data_i[546] : 
                       (N0)? data_i[1228] : 1'b0;
  assign data_o[545] = (N1)? data_i[545] : 
                       (N0)? data_i[1227] : 1'b0;
  assign data_o[544] = (N1)? data_i[544] : 
                       (N0)? data_i[1226] : 1'b0;
  assign data_o[543] = (N1)? data_i[543] : 
                       (N0)? data_i[1225] : 1'b0;
  assign data_o[542] = (N1)? data_i[542] : 
                       (N0)? data_i[1224] : 1'b0;
  assign data_o[541] = (N1)? data_i[541] : 
                       (N0)? data_i[1223] : 1'b0;
  assign data_o[540] = (N1)? data_i[540] : 
                       (N0)? data_i[1222] : 1'b0;
  assign data_o[539] = (N1)? data_i[539] : 
                       (N0)? data_i[1221] : 1'b0;
  assign data_o[538] = (N1)? data_i[538] : 
                       (N0)? data_i[1220] : 1'b0;
  assign data_o[537] = (N1)? data_i[537] : 
                       (N0)? data_i[1219] : 1'b0;
  assign data_o[536] = (N1)? data_i[536] : 
                       (N0)? data_i[1218] : 1'b0;
  assign data_o[535] = (N1)? data_i[535] : 
                       (N0)? data_i[1217] : 1'b0;
  assign data_o[534] = (N1)? data_i[534] : 
                       (N0)? data_i[1216] : 1'b0;
  assign data_o[533] = (N1)? data_i[533] : 
                       (N0)? data_i[1215] : 1'b0;
  assign data_o[532] = (N1)? data_i[532] : 
                       (N0)? data_i[1214] : 1'b0;
  assign data_o[531] = (N1)? data_i[531] : 
                       (N0)? data_i[1213] : 1'b0;
  assign data_o[530] = (N1)? data_i[530] : 
                       (N0)? data_i[1212] : 1'b0;
  assign data_o[529] = (N1)? data_i[529] : 
                       (N0)? data_i[1211] : 1'b0;
  assign data_o[528] = (N1)? data_i[528] : 
                       (N0)? data_i[1210] : 1'b0;
  assign data_o[527] = (N1)? data_i[527] : 
                       (N0)? data_i[1209] : 1'b0;
  assign data_o[526] = (N1)? data_i[526] : 
                       (N0)? data_i[1208] : 1'b0;
  assign data_o[525] = (N1)? data_i[525] : 
                       (N0)? data_i[1207] : 1'b0;
  assign data_o[524] = (N1)? data_i[524] : 
                       (N0)? data_i[1206] : 1'b0;
  assign data_o[523] = (N1)? data_i[523] : 
                       (N0)? data_i[1205] : 1'b0;
  assign data_o[522] = (N1)? data_i[522] : 
                       (N0)? data_i[1204] : 1'b0;
  assign data_o[521] = (N1)? data_i[521] : 
                       (N0)? data_i[1203] : 1'b0;
  assign data_o[520] = (N1)? data_i[520] : 
                       (N0)? data_i[1202] : 1'b0;
  assign data_o[519] = (N1)? data_i[519] : 
                       (N0)? data_i[1201] : 1'b0;
  assign data_o[518] = (N1)? data_i[518] : 
                       (N0)? data_i[1200] : 1'b0;
  assign data_o[517] = (N1)? data_i[517] : 
                       (N0)? data_i[1199] : 1'b0;
  assign data_o[516] = (N1)? data_i[516] : 
                       (N0)? data_i[1198] : 1'b0;
  assign data_o[515] = (N1)? data_i[515] : 
                       (N0)? data_i[1197] : 1'b0;
  assign data_o[514] = (N1)? data_i[514] : 
                       (N0)? data_i[1196] : 1'b0;
  assign data_o[513] = (N1)? data_i[513] : 
                       (N0)? data_i[1195] : 1'b0;
  assign data_o[512] = (N1)? data_i[512] : 
                       (N0)? data_i[1194] : 1'b0;
  assign data_o[511] = (N1)? data_i[511] : 
                       (N0)? data_i[1193] : 1'b0;
  assign data_o[510] = (N1)? data_i[510] : 
                       (N0)? data_i[1192] : 1'b0;
  assign data_o[509] = (N1)? data_i[509] : 
                       (N0)? data_i[1191] : 1'b0;
  assign data_o[508] = (N1)? data_i[508] : 
                       (N0)? data_i[1190] : 1'b0;
  assign data_o[507] = (N1)? data_i[507] : 
                       (N0)? data_i[1189] : 1'b0;
  assign data_o[506] = (N1)? data_i[506] : 
                       (N0)? data_i[1188] : 1'b0;
  assign data_o[505] = (N1)? data_i[505] : 
                       (N0)? data_i[1187] : 1'b0;
  assign data_o[504] = (N1)? data_i[504] : 
                       (N0)? data_i[1186] : 1'b0;
  assign data_o[503] = (N1)? data_i[503] : 
                       (N0)? data_i[1185] : 1'b0;
  assign data_o[502] = (N1)? data_i[502] : 
                       (N0)? data_i[1184] : 1'b0;
  assign data_o[501] = (N1)? data_i[501] : 
                       (N0)? data_i[1183] : 1'b0;
  assign data_o[500] = (N1)? data_i[500] : 
                       (N0)? data_i[1182] : 1'b0;
  assign data_o[499] = (N1)? data_i[499] : 
                       (N0)? data_i[1181] : 1'b0;
  assign data_o[498] = (N1)? data_i[498] : 
                       (N0)? data_i[1180] : 1'b0;
  assign data_o[497] = (N1)? data_i[497] : 
                       (N0)? data_i[1179] : 1'b0;
  assign data_o[496] = (N1)? data_i[496] : 
                       (N0)? data_i[1178] : 1'b0;
  assign data_o[495] = (N1)? data_i[495] : 
                       (N0)? data_i[1177] : 1'b0;
  assign data_o[494] = (N1)? data_i[494] : 
                       (N0)? data_i[1176] : 1'b0;
  assign data_o[493] = (N1)? data_i[493] : 
                       (N0)? data_i[1175] : 1'b0;
  assign data_o[492] = (N1)? data_i[492] : 
                       (N0)? data_i[1174] : 1'b0;
  assign data_o[491] = (N1)? data_i[491] : 
                       (N0)? data_i[1173] : 1'b0;
  assign data_o[490] = (N1)? data_i[490] : 
                       (N0)? data_i[1172] : 1'b0;
  assign data_o[489] = (N1)? data_i[489] : 
                       (N0)? data_i[1171] : 1'b0;
  assign data_o[488] = (N1)? data_i[488] : 
                       (N0)? data_i[1170] : 1'b0;
  assign data_o[487] = (N1)? data_i[487] : 
                       (N0)? data_i[1169] : 1'b0;
  assign data_o[486] = (N1)? data_i[486] : 
                       (N0)? data_i[1168] : 1'b0;
  assign data_o[485] = (N1)? data_i[485] : 
                       (N0)? data_i[1167] : 1'b0;
  assign data_o[484] = (N1)? data_i[484] : 
                       (N0)? data_i[1166] : 1'b0;
  assign data_o[483] = (N1)? data_i[483] : 
                       (N0)? data_i[1165] : 1'b0;
  assign data_o[482] = (N1)? data_i[482] : 
                       (N0)? data_i[1164] : 1'b0;
  assign data_o[481] = (N1)? data_i[481] : 
                       (N0)? data_i[1163] : 1'b0;
  assign data_o[480] = (N1)? data_i[480] : 
                       (N0)? data_i[1162] : 1'b0;
  assign data_o[479] = (N1)? data_i[479] : 
                       (N0)? data_i[1161] : 1'b0;
  assign data_o[478] = (N1)? data_i[478] : 
                       (N0)? data_i[1160] : 1'b0;
  assign data_o[477] = (N1)? data_i[477] : 
                       (N0)? data_i[1159] : 1'b0;
  assign data_o[476] = (N1)? data_i[476] : 
                       (N0)? data_i[1158] : 1'b0;
  assign data_o[475] = (N1)? data_i[475] : 
                       (N0)? data_i[1157] : 1'b0;
  assign data_o[474] = (N1)? data_i[474] : 
                       (N0)? data_i[1156] : 1'b0;
  assign data_o[473] = (N1)? data_i[473] : 
                       (N0)? data_i[1155] : 1'b0;
  assign data_o[472] = (N1)? data_i[472] : 
                       (N0)? data_i[1154] : 1'b0;
  assign data_o[471] = (N1)? data_i[471] : 
                       (N0)? data_i[1153] : 1'b0;
  assign data_o[470] = (N1)? data_i[470] : 
                       (N0)? data_i[1152] : 1'b0;
  assign data_o[469] = (N1)? data_i[469] : 
                       (N0)? data_i[1151] : 1'b0;
  assign data_o[468] = (N1)? data_i[468] : 
                       (N0)? data_i[1150] : 1'b0;
  assign data_o[467] = (N1)? data_i[467] : 
                       (N0)? data_i[1149] : 1'b0;
  assign data_o[466] = (N1)? data_i[466] : 
                       (N0)? data_i[1148] : 1'b0;
  assign data_o[465] = (N1)? data_i[465] : 
                       (N0)? data_i[1147] : 1'b0;
  assign data_o[464] = (N1)? data_i[464] : 
                       (N0)? data_i[1146] : 1'b0;
  assign data_o[463] = (N1)? data_i[463] : 
                       (N0)? data_i[1145] : 1'b0;
  assign data_o[462] = (N1)? data_i[462] : 
                       (N0)? data_i[1144] : 1'b0;
  assign data_o[461] = (N1)? data_i[461] : 
                       (N0)? data_i[1143] : 1'b0;
  assign data_o[460] = (N1)? data_i[460] : 
                       (N0)? data_i[1142] : 1'b0;
  assign data_o[459] = (N1)? data_i[459] : 
                       (N0)? data_i[1141] : 1'b0;
  assign data_o[458] = (N1)? data_i[458] : 
                       (N0)? data_i[1140] : 1'b0;
  assign data_o[457] = (N1)? data_i[457] : 
                       (N0)? data_i[1139] : 1'b0;
  assign data_o[456] = (N1)? data_i[456] : 
                       (N0)? data_i[1138] : 1'b0;
  assign data_o[455] = (N1)? data_i[455] : 
                       (N0)? data_i[1137] : 1'b0;
  assign data_o[454] = (N1)? data_i[454] : 
                       (N0)? data_i[1136] : 1'b0;
  assign data_o[453] = (N1)? data_i[453] : 
                       (N0)? data_i[1135] : 1'b0;
  assign data_o[452] = (N1)? data_i[452] : 
                       (N0)? data_i[1134] : 1'b0;
  assign data_o[451] = (N1)? data_i[451] : 
                       (N0)? data_i[1133] : 1'b0;
  assign data_o[450] = (N1)? data_i[450] : 
                       (N0)? data_i[1132] : 1'b0;
  assign data_o[449] = (N1)? data_i[449] : 
                       (N0)? data_i[1131] : 1'b0;
  assign data_o[448] = (N1)? data_i[448] : 
                       (N0)? data_i[1130] : 1'b0;
  assign data_o[447] = (N1)? data_i[447] : 
                       (N0)? data_i[1129] : 1'b0;
  assign data_o[446] = (N1)? data_i[446] : 
                       (N0)? data_i[1128] : 1'b0;
  assign data_o[445] = (N1)? data_i[445] : 
                       (N0)? data_i[1127] : 1'b0;
  assign data_o[444] = (N1)? data_i[444] : 
                       (N0)? data_i[1126] : 1'b0;
  assign data_o[443] = (N1)? data_i[443] : 
                       (N0)? data_i[1125] : 1'b0;
  assign data_o[442] = (N1)? data_i[442] : 
                       (N0)? data_i[1124] : 1'b0;
  assign data_o[441] = (N1)? data_i[441] : 
                       (N0)? data_i[1123] : 1'b0;
  assign data_o[440] = (N1)? data_i[440] : 
                       (N0)? data_i[1122] : 1'b0;
  assign data_o[439] = (N1)? data_i[439] : 
                       (N0)? data_i[1121] : 1'b0;
  assign data_o[438] = (N1)? data_i[438] : 
                       (N0)? data_i[1120] : 1'b0;
  assign data_o[437] = (N1)? data_i[437] : 
                       (N0)? data_i[1119] : 1'b0;
  assign data_o[436] = (N1)? data_i[436] : 
                       (N0)? data_i[1118] : 1'b0;
  assign data_o[435] = (N1)? data_i[435] : 
                       (N0)? data_i[1117] : 1'b0;
  assign data_o[434] = (N1)? data_i[434] : 
                       (N0)? data_i[1116] : 1'b0;
  assign data_o[433] = (N1)? data_i[433] : 
                       (N0)? data_i[1115] : 1'b0;
  assign data_o[432] = (N1)? data_i[432] : 
                       (N0)? data_i[1114] : 1'b0;
  assign data_o[431] = (N1)? data_i[431] : 
                       (N0)? data_i[1113] : 1'b0;
  assign data_o[430] = (N1)? data_i[430] : 
                       (N0)? data_i[1112] : 1'b0;
  assign data_o[429] = (N1)? data_i[429] : 
                       (N0)? data_i[1111] : 1'b0;
  assign data_o[428] = (N1)? data_i[428] : 
                       (N0)? data_i[1110] : 1'b0;
  assign data_o[427] = (N1)? data_i[427] : 
                       (N0)? data_i[1109] : 1'b0;
  assign data_o[426] = (N1)? data_i[426] : 
                       (N0)? data_i[1108] : 1'b0;
  assign data_o[425] = (N1)? data_i[425] : 
                       (N0)? data_i[1107] : 1'b0;
  assign data_o[424] = (N1)? data_i[424] : 
                       (N0)? data_i[1106] : 1'b0;
  assign data_o[423] = (N1)? data_i[423] : 
                       (N0)? data_i[1105] : 1'b0;
  assign data_o[422] = (N1)? data_i[422] : 
                       (N0)? data_i[1104] : 1'b0;
  assign data_o[421] = (N1)? data_i[421] : 
                       (N0)? data_i[1103] : 1'b0;
  assign data_o[420] = (N1)? data_i[420] : 
                       (N0)? data_i[1102] : 1'b0;
  assign data_o[419] = (N1)? data_i[419] : 
                       (N0)? data_i[1101] : 1'b0;
  assign data_o[418] = (N1)? data_i[418] : 
                       (N0)? data_i[1100] : 1'b0;
  assign data_o[417] = (N1)? data_i[417] : 
                       (N0)? data_i[1099] : 1'b0;
  assign data_o[416] = (N1)? data_i[416] : 
                       (N0)? data_i[1098] : 1'b0;
  assign data_o[415] = (N1)? data_i[415] : 
                       (N0)? data_i[1097] : 1'b0;
  assign data_o[414] = (N1)? data_i[414] : 
                       (N0)? data_i[1096] : 1'b0;
  assign data_o[413] = (N1)? data_i[413] : 
                       (N0)? data_i[1095] : 1'b0;
  assign data_o[412] = (N1)? data_i[412] : 
                       (N0)? data_i[1094] : 1'b0;
  assign data_o[411] = (N1)? data_i[411] : 
                       (N0)? data_i[1093] : 1'b0;
  assign data_o[410] = (N1)? data_i[410] : 
                       (N0)? data_i[1092] : 1'b0;
  assign data_o[409] = (N1)? data_i[409] : 
                       (N0)? data_i[1091] : 1'b0;
  assign data_o[408] = (N1)? data_i[408] : 
                       (N0)? data_i[1090] : 1'b0;
  assign data_o[407] = (N1)? data_i[407] : 
                       (N0)? data_i[1089] : 1'b0;
  assign data_o[406] = (N1)? data_i[406] : 
                       (N0)? data_i[1088] : 1'b0;
  assign data_o[405] = (N1)? data_i[405] : 
                       (N0)? data_i[1087] : 1'b0;
  assign data_o[404] = (N1)? data_i[404] : 
                       (N0)? data_i[1086] : 1'b0;
  assign data_o[403] = (N1)? data_i[403] : 
                       (N0)? data_i[1085] : 1'b0;
  assign data_o[402] = (N1)? data_i[402] : 
                       (N0)? data_i[1084] : 1'b0;
  assign data_o[401] = (N1)? data_i[401] : 
                       (N0)? data_i[1083] : 1'b0;
  assign data_o[400] = (N1)? data_i[400] : 
                       (N0)? data_i[1082] : 1'b0;
  assign data_o[399] = (N1)? data_i[399] : 
                       (N0)? data_i[1081] : 1'b0;
  assign data_o[398] = (N1)? data_i[398] : 
                       (N0)? data_i[1080] : 1'b0;
  assign data_o[397] = (N1)? data_i[397] : 
                       (N0)? data_i[1079] : 1'b0;
  assign data_o[396] = (N1)? data_i[396] : 
                       (N0)? data_i[1078] : 1'b0;
  assign data_o[395] = (N1)? data_i[395] : 
                       (N0)? data_i[1077] : 1'b0;
  assign data_o[394] = (N1)? data_i[394] : 
                       (N0)? data_i[1076] : 1'b0;
  assign data_o[393] = (N1)? data_i[393] : 
                       (N0)? data_i[1075] : 1'b0;
  assign data_o[392] = (N1)? data_i[392] : 
                       (N0)? data_i[1074] : 1'b0;
  assign data_o[391] = (N1)? data_i[391] : 
                       (N0)? data_i[1073] : 1'b0;
  assign data_o[390] = (N1)? data_i[390] : 
                       (N0)? data_i[1072] : 1'b0;
  assign data_o[389] = (N1)? data_i[389] : 
                       (N0)? data_i[1071] : 1'b0;
  assign data_o[388] = (N1)? data_i[388] : 
                       (N0)? data_i[1070] : 1'b0;
  assign data_o[387] = (N1)? data_i[387] : 
                       (N0)? data_i[1069] : 1'b0;
  assign data_o[386] = (N1)? data_i[386] : 
                       (N0)? data_i[1068] : 1'b0;
  assign data_o[385] = (N1)? data_i[385] : 
                       (N0)? data_i[1067] : 1'b0;
  assign data_o[384] = (N1)? data_i[384] : 
                       (N0)? data_i[1066] : 1'b0;
  assign data_o[383] = (N1)? data_i[383] : 
                       (N0)? data_i[1065] : 1'b0;
  assign data_o[382] = (N1)? data_i[382] : 
                       (N0)? data_i[1064] : 1'b0;
  assign data_o[381] = (N1)? data_i[381] : 
                       (N0)? data_i[1063] : 1'b0;
  assign data_o[380] = (N1)? data_i[380] : 
                       (N0)? data_i[1062] : 1'b0;
  assign data_o[379] = (N1)? data_i[379] : 
                       (N0)? data_i[1061] : 1'b0;
  assign data_o[378] = (N1)? data_i[378] : 
                       (N0)? data_i[1060] : 1'b0;
  assign data_o[377] = (N1)? data_i[377] : 
                       (N0)? data_i[1059] : 1'b0;
  assign data_o[376] = (N1)? data_i[376] : 
                       (N0)? data_i[1058] : 1'b0;
  assign data_o[375] = (N1)? data_i[375] : 
                       (N0)? data_i[1057] : 1'b0;
  assign data_o[374] = (N1)? data_i[374] : 
                       (N0)? data_i[1056] : 1'b0;
  assign data_o[373] = (N1)? data_i[373] : 
                       (N0)? data_i[1055] : 1'b0;
  assign data_o[372] = (N1)? data_i[372] : 
                       (N0)? data_i[1054] : 1'b0;
  assign data_o[371] = (N1)? data_i[371] : 
                       (N0)? data_i[1053] : 1'b0;
  assign data_o[370] = (N1)? data_i[370] : 
                       (N0)? data_i[1052] : 1'b0;
  assign data_o[369] = (N1)? data_i[369] : 
                       (N0)? data_i[1051] : 1'b0;
  assign data_o[368] = (N1)? data_i[368] : 
                       (N0)? data_i[1050] : 1'b0;
  assign data_o[367] = (N1)? data_i[367] : 
                       (N0)? data_i[1049] : 1'b0;
  assign data_o[366] = (N1)? data_i[366] : 
                       (N0)? data_i[1048] : 1'b0;
  assign data_o[365] = (N1)? data_i[365] : 
                       (N0)? data_i[1047] : 1'b0;
  assign data_o[364] = (N1)? data_i[364] : 
                       (N0)? data_i[1046] : 1'b0;
  assign data_o[363] = (N1)? data_i[363] : 
                       (N0)? data_i[1045] : 1'b0;
  assign data_o[362] = (N1)? data_i[362] : 
                       (N0)? data_i[1044] : 1'b0;
  assign data_o[361] = (N1)? data_i[361] : 
                       (N0)? data_i[1043] : 1'b0;
  assign data_o[360] = (N1)? data_i[360] : 
                       (N0)? data_i[1042] : 1'b0;
  assign data_o[359] = (N1)? data_i[359] : 
                       (N0)? data_i[1041] : 1'b0;
  assign data_o[358] = (N1)? data_i[358] : 
                       (N0)? data_i[1040] : 1'b0;
  assign data_o[357] = (N1)? data_i[357] : 
                       (N0)? data_i[1039] : 1'b0;
  assign data_o[356] = (N1)? data_i[356] : 
                       (N0)? data_i[1038] : 1'b0;
  assign data_o[355] = (N1)? data_i[355] : 
                       (N0)? data_i[1037] : 1'b0;
  assign data_o[354] = (N1)? data_i[354] : 
                       (N0)? data_i[1036] : 1'b0;
  assign data_o[353] = (N1)? data_i[353] : 
                       (N0)? data_i[1035] : 1'b0;
  assign data_o[352] = (N1)? data_i[352] : 
                       (N0)? data_i[1034] : 1'b0;
  assign data_o[351] = (N1)? data_i[351] : 
                       (N0)? data_i[1033] : 1'b0;
  assign data_o[350] = (N1)? data_i[350] : 
                       (N0)? data_i[1032] : 1'b0;
  assign data_o[349] = (N1)? data_i[349] : 
                       (N0)? data_i[1031] : 1'b0;
  assign data_o[348] = (N1)? data_i[348] : 
                       (N0)? data_i[1030] : 1'b0;
  assign data_o[347] = (N1)? data_i[347] : 
                       (N0)? data_i[1029] : 1'b0;
  assign data_o[346] = (N1)? data_i[346] : 
                       (N0)? data_i[1028] : 1'b0;
  assign data_o[345] = (N1)? data_i[345] : 
                       (N0)? data_i[1027] : 1'b0;
  assign data_o[344] = (N1)? data_i[344] : 
                       (N0)? data_i[1026] : 1'b0;
  assign data_o[343] = (N1)? data_i[343] : 
                       (N0)? data_i[1025] : 1'b0;
  assign data_o[342] = (N1)? data_i[342] : 
                       (N0)? data_i[1024] : 1'b0;
  assign data_o[341] = (N1)? data_i[341] : 
                       (N0)? data_i[1023] : 1'b0;
  assign data_o[340] = (N1)? data_i[340] : 
                       (N0)? data_i[1022] : 1'b0;
  assign data_o[339] = (N1)? data_i[339] : 
                       (N0)? data_i[1021] : 1'b0;
  assign data_o[338] = (N1)? data_i[338] : 
                       (N0)? data_i[1020] : 1'b0;
  assign data_o[337] = (N1)? data_i[337] : 
                       (N0)? data_i[1019] : 1'b0;
  assign data_o[336] = (N1)? data_i[336] : 
                       (N0)? data_i[1018] : 1'b0;
  assign data_o[335] = (N1)? data_i[335] : 
                       (N0)? data_i[1017] : 1'b0;
  assign data_o[334] = (N1)? data_i[334] : 
                       (N0)? data_i[1016] : 1'b0;
  assign data_o[333] = (N1)? data_i[333] : 
                       (N0)? data_i[1015] : 1'b0;
  assign data_o[332] = (N1)? data_i[332] : 
                       (N0)? data_i[1014] : 1'b0;
  assign data_o[331] = (N1)? data_i[331] : 
                       (N0)? data_i[1013] : 1'b0;
  assign data_o[330] = (N1)? data_i[330] : 
                       (N0)? data_i[1012] : 1'b0;
  assign data_o[329] = (N1)? data_i[329] : 
                       (N0)? data_i[1011] : 1'b0;
  assign data_o[328] = (N1)? data_i[328] : 
                       (N0)? data_i[1010] : 1'b0;
  assign data_o[327] = (N1)? data_i[327] : 
                       (N0)? data_i[1009] : 1'b0;
  assign data_o[326] = (N1)? data_i[326] : 
                       (N0)? data_i[1008] : 1'b0;
  assign data_o[325] = (N1)? data_i[325] : 
                       (N0)? data_i[1007] : 1'b0;
  assign data_o[324] = (N1)? data_i[324] : 
                       (N0)? data_i[1006] : 1'b0;
  assign data_o[323] = (N1)? data_i[323] : 
                       (N0)? data_i[1005] : 1'b0;
  assign data_o[322] = (N1)? data_i[322] : 
                       (N0)? data_i[1004] : 1'b0;
  assign data_o[321] = (N1)? data_i[321] : 
                       (N0)? data_i[1003] : 1'b0;
  assign data_o[320] = (N1)? data_i[320] : 
                       (N0)? data_i[1002] : 1'b0;
  assign data_o[319] = (N1)? data_i[319] : 
                       (N0)? data_i[1001] : 1'b0;
  assign data_o[318] = (N1)? data_i[318] : 
                       (N0)? data_i[1000] : 1'b0;
  assign data_o[317] = (N1)? data_i[317] : 
                       (N0)? data_i[999] : 1'b0;
  assign data_o[316] = (N1)? data_i[316] : 
                       (N0)? data_i[998] : 1'b0;
  assign data_o[315] = (N1)? data_i[315] : 
                       (N0)? data_i[997] : 1'b0;
  assign data_o[314] = (N1)? data_i[314] : 
                       (N0)? data_i[996] : 1'b0;
  assign data_o[313] = (N1)? data_i[313] : 
                       (N0)? data_i[995] : 1'b0;
  assign data_o[312] = (N1)? data_i[312] : 
                       (N0)? data_i[994] : 1'b0;
  assign data_o[311] = (N1)? data_i[311] : 
                       (N0)? data_i[993] : 1'b0;
  assign data_o[310] = (N1)? data_i[310] : 
                       (N0)? data_i[992] : 1'b0;
  assign data_o[309] = (N1)? data_i[309] : 
                       (N0)? data_i[991] : 1'b0;
  assign data_o[308] = (N1)? data_i[308] : 
                       (N0)? data_i[990] : 1'b0;
  assign data_o[307] = (N1)? data_i[307] : 
                       (N0)? data_i[989] : 1'b0;
  assign data_o[306] = (N1)? data_i[306] : 
                       (N0)? data_i[988] : 1'b0;
  assign data_o[305] = (N1)? data_i[305] : 
                       (N0)? data_i[987] : 1'b0;
  assign data_o[304] = (N1)? data_i[304] : 
                       (N0)? data_i[986] : 1'b0;
  assign data_o[303] = (N1)? data_i[303] : 
                       (N0)? data_i[985] : 1'b0;
  assign data_o[302] = (N1)? data_i[302] : 
                       (N0)? data_i[984] : 1'b0;
  assign data_o[301] = (N1)? data_i[301] : 
                       (N0)? data_i[983] : 1'b0;
  assign data_o[300] = (N1)? data_i[300] : 
                       (N0)? data_i[982] : 1'b0;
  assign data_o[299] = (N1)? data_i[299] : 
                       (N0)? data_i[981] : 1'b0;
  assign data_o[298] = (N1)? data_i[298] : 
                       (N0)? data_i[980] : 1'b0;
  assign data_o[297] = (N1)? data_i[297] : 
                       (N0)? data_i[979] : 1'b0;
  assign data_o[296] = (N1)? data_i[296] : 
                       (N0)? data_i[978] : 1'b0;
  assign data_o[295] = (N1)? data_i[295] : 
                       (N0)? data_i[977] : 1'b0;
  assign data_o[294] = (N1)? data_i[294] : 
                       (N0)? data_i[976] : 1'b0;
  assign data_o[293] = (N1)? data_i[293] : 
                       (N0)? data_i[975] : 1'b0;
  assign data_o[292] = (N1)? data_i[292] : 
                       (N0)? data_i[974] : 1'b0;
  assign data_o[291] = (N1)? data_i[291] : 
                       (N0)? data_i[973] : 1'b0;
  assign data_o[290] = (N1)? data_i[290] : 
                       (N0)? data_i[972] : 1'b0;
  assign data_o[289] = (N1)? data_i[289] : 
                       (N0)? data_i[971] : 1'b0;
  assign data_o[288] = (N1)? data_i[288] : 
                       (N0)? data_i[970] : 1'b0;
  assign data_o[287] = (N1)? data_i[287] : 
                       (N0)? data_i[969] : 1'b0;
  assign data_o[286] = (N1)? data_i[286] : 
                       (N0)? data_i[968] : 1'b0;
  assign data_o[285] = (N1)? data_i[285] : 
                       (N0)? data_i[967] : 1'b0;
  assign data_o[284] = (N1)? data_i[284] : 
                       (N0)? data_i[966] : 1'b0;
  assign data_o[283] = (N1)? data_i[283] : 
                       (N0)? data_i[965] : 1'b0;
  assign data_o[282] = (N1)? data_i[282] : 
                       (N0)? data_i[964] : 1'b0;
  assign data_o[281] = (N1)? data_i[281] : 
                       (N0)? data_i[963] : 1'b0;
  assign data_o[280] = (N1)? data_i[280] : 
                       (N0)? data_i[962] : 1'b0;
  assign data_o[279] = (N1)? data_i[279] : 
                       (N0)? data_i[961] : 1'b0;
  assign data_o[278] = (N1)? data_i[278] : 
                       (N0)? data_i[960] : 1'b0;
  assign data_o[277] = (N1)? data_i[277] : 
                       (N0)? data_i[959] : 1'b0;
  assign data_o[276] = (N1)? data_i[276] : 
                       (N0)? data_i[958] : 1'b0;
  assign data_o[275] = (N1)? data_i[275] : 
                       (N0)? data_i[957] : 1'b0;
  assign data_o[274] = (N1)? data_i[274] : 
                       (N0)? data_i[956] : 1'b0;
  assign data_o[273] = (N1)? data_i[273] : 
                       (N0)? data_i[955] : 1'b0;
  assign data_o[272] = (N1)? data_i[272] : 
                       (N0)? data_i[954] : 1'b0;
  assign data_o[271] = (N1)? data_i[271] : 
                       (N0)? data_i[953] : 1'b0;
  assign data_o[270] = (N1)? data_i[270] : 
                       (N0)? data_i[952] : 1'b0;
  assign data_o[269] = (N1)? data_i[269] : 
                       (N0)? data_i[951] : 1'b0;
  assign data_o[268] = (N1)? data_i[268] : 
                       (N0)? data_i[950] : 1'b0;
  assign data_o[267] = (N1)? data_i[267] : 
                       (N0)? data_i[949] : 1'b0;
  assign data_o[266] = (N1)? data_i[266] : 
                       (N0)? data_i[948] : 1'b0;
  assign data_o[265] = (N1)? data_i[265] : 
                       (N0)? data_i[947] : 1'b0;
  assign data_o[264] = (N1)? data_i[264] : 
                       (N0)? data_i[946] : 1'b0;
  assign data_o[263] = (N1)? data_i[263] : 
                       (N0)? data_i[945] : 1'b0;
  assign data_o[262] = (N1)? data_i[262] : 
                       (N0)? data_i[944] : 1'b0;
  assign data_o[261] = (N1)? data_i[261] : 
                       (N0)? data_i[943] : 1'b0;
  assign data_o[260] = (N1)? data_i[260] : 
                       (N0)? data_i[942] : 1'b0;
  assign data_o[259] = (N1)? data_i[259] : 
                       (N0)? data_i[941] : 1'b0;
  assign data_o[258] = (N1)? data_i[258] : 
                       (N0)? data_i[940] : 1'b0;
  assign data_o[257] = (N1)? data_i[257] : 
                       (N0)? data_i[939] : 1'b0;
  assign data_o[256] = (N1)? data_i[256] : 
                       (N0)? data_i[938] : 1'b0;
  assign data_o[255] = (N1)? data_i[255] : 
                       (N0)? data_i[937] : 1'b0;
  assign data_o[254] = (N1)? data_i[254] : 
                       (N0)? data_i[936] : 1'b0;
  assign data_o[253] = (N1)? data_i[253] : 
                       (N0)? data_i[935] : 1'b0;
  assign data_o[252] = (N1)? data_i[252] : 
                       (N0)? data_i[934] : 1'b0;
  assign data_o[251] = (N1)? data_i[251] : 
                       (N0)? data_i[933] : 1'b0;
  assign data_o[250] = (N1)? data_i[250] : 
                       (N0)? data_i[932] : 1'b0;
  assign data_o[249] = (N1)? data_i[249] : 
                       (N0)? data_i[931] : 1'b0;
  assign data_o[248] = (N1)? data_i[248] : 
                       (N0)? data_i[930] : 1'b0;
  assign data_o[247] = (N1)? data_i[247] : 
                       (N0)? data_i[929] : 1'b0;
  assign data_o[246] = (N1)? data_i[246] : 
                       (N0)? data_i[928] : 1'b0;
  assign data_o[245] = (N1)? data_i[245] : 
                       (N0)? data_i[927] : 1'b0;
  assign data_o[244] = (N1)? data_i[244] : 
                       (N0)? data_i[926] : 1'b0;
  assign data_o[243] = (N1)? data_i[243] : 
                       (N0)? data_i[925] : 1'b0;
  assign data_o[242] = (N1)? data_i[242] : 
                       (N0)? data_i[924] : 1'b0;
  assign data_o[241] = (N1)? data_i[241] : 
                       (N0)? data_i[923] : 1'b0;
  assign data_o[240] = (N1)? data_i[240] : 
                       (N0)? data_i[922] : 1'b0;
  assign data_o[239] = (N1)? data_i[239] : 
                       (N0)? data_i[921] : 1'b0;
  assign data_o[238] = (N1)? data_i[238] : 
                       (N0)? data_i[920] : 1'b0;
  assign data_o[237] = (N1)? data_i[237] : 
                       (N0)? data_i[919] : 1'b0;
  assign data_o[236] = (N1)? data_i[236] : 
                       (N0)? data_i[918] : 1'b0;
  assign data_o[235] = (N1)? data_i[235] : 
                       (N0)? data_i[917] : 1'b0;
  assign data_o[234] = (N1)? data_i[234] : 
                       (N0)? data_i[916] : 1'b0;
  assign data_o[233] = (N1)? data_i[233] : 
                       (N0)? data_i[915] : 1'b0;
  assign data_o[232] = (N1)? data_i[232] : 
                       (N0)? data_i[914] : 1'b0;
  assign data_o[231] = (N1)? data_i[231] : 
                       (N0)? data_i[913] : 1'b0;
  assign data_o[230] = (N1)? data_i[230] : 
                       (N0)? data_i[912] : 1'b0;
  assign data_o[229] = (N1)? data_i[229] : 
                       (N0)? data_i[911] : 1'b0;
  assign data_o[228] = (N1)? data_i[228] : 
                       (N0)? data_i[910] : 1'b0;
  assign data_o[227] = (N1)? data_i[227] : 
                       (N0)? data_i[909] : 1'b0;
  assign data_o[226] = (N1)? data_i[226] : 
                       (N0)? data_i[908] : 1'b0;
  assign data_o[225] = (N1)? data_i[225] : 
                       (N0)? data_i[907] : 1'b0;
  assign data_o[224] = (N1)? data_i[224] : 
                       (N0)? data_i[906] : 1'b0;
  assign data_o[223] = (N1)? data_i[223] : 
                       (N0)? data_i[905] : 1'b0;
  assign data_o[222] = (N1)? data_i[222] : 
                       (N0)? data_i[904] : 1'b0;
  assign data_o[221] = (N1)? data_i[221] : 
                       (N0)? data_i[903] : 1'b0;
  assign data_o[220] = (N1)? data_i[220] : 
                       (N0)? data_i[902] : 1'b0;
  assign data_o[219] = (N1)? data_i[219] : 
                       (N0)? data_i[901] : 1'b0;
  assign data_o[218] = (N1)? data_i[218] : 
                       (N0)? data_i[900] : 1'b0;
  assign data_o[217] = (N1)? data_i[217] : 
                       (N0)? data_i[899] : 1'b0;
  assign data_o[216] = (N1)? data_i[216] : 
                       (N0)? data_i[898] : 1'b0;
  assign data_o[215] = (N1)? data_i[215] : 
                       (N0)? data_i[897] : 1'b0;
  assign data_o[214] = (N1)? data_i[214] : 
                       (N0)? data_i[896] : 1'b0;
  assign data_o[213] = (N1)? data_i[213] : 
                       (N0)? data_i[895] : 1'b0;
  assign data_o[212] = (N1)? data_i[212] : 
                       (N0)? data_i[894] : 1'b0;
  assign data_o[211] = (N1)? data_i[211] : 
                       (N0)? data_i[893] : 1'b0;
  assign data_o[210] = (N1)? data_i[210] : 
                       (N0)? data_i[892] : 1'b0;
  assign data_o[209] = (N1)? data_i[209] : 
                       (N0)? data_i[891] : 1'b0;
  assign data_o[208] = (N1)? data_i[208] : 
                       (N0)? data_i[890] : 1'b0;
  assign data_o[207] = (N1)? data_i[207] : 
                       (N0)? data_i[889] : 1'b0;
  assign data_o[206] = (N1)? data_i[206] : 
                       (N0)? data_i[888] : 1'b0;
  assign data_o[205] = (N1)? data_i[205] : 
                       (N0)? data_i[887] : 1'b0;
  assign data_o[204] = (N1)? data_i[204] : 
                       (N0)? data_i[886] : 1'b0;
  assign data_o[203] = (N1)? data_i[203] : 
                       (N0)? data_i[885] : 1'b0;
  assign data_o[202] = (N1)? data_i[202] : 
                       (N0)? data_i[884] : 1'b0;
  assign data_o[201] = (N1)? data_i[201] : 
                       (N0)? data_i[883] : 1'b0;
  assign data_o[200] = (N1)? data_i[200] : 
                       (N0)? data_i[882] : 1'b0;
  assign data_o[199] = (N1)? data_i[199] : 
                       (N0)? data_i[881] : 1'b0;
  assign data_o[198] = (N1)? data_i[198] : 
                       (N0)? data_i[880] : 1'b0;
  assign data_o[197] = (N1)? data_i[197] : 
                       (N0)? data_i[879] : 1'b0;
  assign data_o[196] = (N1)? data_i[196] : 
                       (N0)? data_i[878] : 1'b0;
  assign data_o[195] = (N1)? data_i[195] : 
                       (N0)? data_i[877] : 1'b0;
  assign data_o[194] = (N1)? data_i[194] : 
                       (N0)? data_i[876] : 1'b0;
  assign data_o[193] = (N1)? data_i[193] : 
                       (N0)? data_i[875] : 1'b0;
  assign data_o[192] = (N1)? data_i[192] : 
                       (N0)? data_i[874] : 1'b0;
  assign data_o[191] = (N1)? data_i[191] : 
                       (N0)? data_i[873] : 1'b0;
  assign data_o[190] = (N1)? data_i[190] : 
                       (N0)? data_i[872] : 1'b0;
  assign data_o[189] = (N1)? data_i[189] : 
                       (N0)? data_i[871] : 1'b0;
  assign data_o[188] = (N1)? data_i[188] : 
                       (N0)? data_i[870] : 1'b0;
  assign data_o[187] = (N1)? data_i[187] : 
                       (N0)? data_i[869] : 1'b0;
  assign data_o[186] = (N1)? data_i[186] : 
                       (N0)? data_i[868] : 1'b0;
  assign data_o[185] = (N1)? data_i[185] : 
                       (N0)? data_i[867] : 1'b0;
  assign data_o[184] = (N1)? data_i[184] : 
                       (N0)? data_i[866] : 1'b0;
  assign data_o[183] = (N1)? data_i[183] : 
                       (N0)? data_i[865] : 1'b0;
  assign data_o[182] = (N1)? data_i[182] : 
                       (N0)? data_i[864] : 1'b0;
  assign data_o[181] = (N1)? data_i[181] : 
                       (N0)? data_i[863] : 1'b0;
  assign data_o[180] = (N1)? data_i[180] : 
                       (N0)? data_i[862] : 1'b0;
  assign data_o[179] = (N1)? data_i[179] : 
                       (N0)? data_i[861] : 1'b0;
  assign data_o[178] = (N1)? data_i[178] : 
                       (N0)? data_i[860] : 1'b0;
  assign data_o[177] = (N1)? data_i[177] : 
                       (N0)? data_i[859] : 1'b0;
  assign data_o[176] = (N1)? data_i[176] : 
                       (N0)? data_i[858] : 1'b0;
  assign data_o[175] = (N1)? data_i[175] : 
                       (N0)? data_i[857] : 1'b0;
  assign data_o[174] = (N1)? data_i[174] : 
                       (N0)? data_i[856] : 1'b0;
  assign data_o[173] = (N1)? data_i[173] : 
                       (N0)? data_i[855] : 1'b0;
  assign data_o[172] = (N1)? data_i[172] : 
                       (N0)? data_i[854] : 1'b0;
  assign data_o[171] = (N1)? data_i[171] : 
                       (N0)? data_i[853] : 1'b0;
  assign data_o[170] = (N1)? data_i[170] : 
                       (N0)? data_i[852] : 1'b0;
  assign data_o[169] = (N1)? data_i[169] : 
                       (N0)? data_i[851] : 1'b0;
  assign data_o[168] = (N1)? data_i[168] : 
                       (N0)? data_i[850] : 1'b0;
  assign data_o[167] = (N1)? data_i[167] : 
                       (N0)? data_i[849] : 1'b0;
  assign data_o[166] = (N1)? data_i[166] : 
                       (N0)? data_i[848] : 1'b0;
  assign data_o[165] = (N1)? data_i[165] : 
                       (N0)? data_i[847] : 1'b0;
  assign data_o[164] = (N1)? data_i[164] : 
                       (N0)? data_i[846] : 1'b0;
  assign data_o[163] = (N1)? data_i[163] : 
                       (N0)? data_i[845] : 1'b0;
  assign data_o[162] = (N1)? data_i[162] : 
                       (N0)? data_i[844] : 1'b0;
  assign data_o[161] = (N1)? data_i[161] : 
                       (N0)? data_i[843] : 1'b0;
  assign data_o[160] = (N1)? data_i[160] : 
                       (N0)? data_i[842] : 1'b0;
  assign data_o[159] = (N1)? data_i[159] : 
                       (N0)? data_i[841] : 1'b0;
  assign data_o[158] = (N1)? data_i[158] : 
                       (N0)? data_i[840] : 1'b0;
  assign data_o[157] = (N1)? data_i[157] : 
                       (N0)? data_i[839] : 1'b0;
  assign data_o[156] = (N1)? data_i[156] : 
                       (N0)? data_i[838] : 1'b0;
  assign data_o[155] = (N1)? data_i[155] : 
                       (N0)? data_i[837] : 1'b0;
  assign data_o[154] = (N1)? data_i[154] : 
                       (N0)? data_i[836] : 1'b0;
  assign data_o[153] = (N1)? data_i[153] : 
                       (N0)? data_i[835] : 1'b0;
  assign data_o[152] = (N1)? data_i[152] : 
                       (N0)? data_i[834] : 1'b0;
  assign data_o[151] = (N1)? data_i[151] : 
                       (N0)? data_i[833] : 1'b0;
  assign data_o[150] = (N1)? data_i[150] : 
                       (N0)? data_i[832] : 1'b0;
  assign data_o[149] = (N1)? data_i[149] : 
                       (N0)? data_i[831] : 1'b0;
  assign data_o[148] = (N1)? data_i[148] : 
                       (N0)? data_i[830] : 1'b0;
  assign data_o[147] = (N1)? data_i[147] : 
                       (N0)? data_i[829] : 1'b0;
  assign data_o[146] = (N1)? data_i[146] : 
                       (N0)? data_i[828] : 1'b0;
  assign data_o[145] = (N1)? data_i[145] : 
                       (N0)? data_i[827] : 1'b0;
  assign data_o[144] = (N1)? data_i[144] : 
                       (N0)? data_i[826] : 1'b0;
  assign data_o[143] = (N1)? data_i[143] : 
                       (N0)? data_i[825] : 1'b0;
  assign data_o[142] = (N1)? data_i[142] : 
                       (N0)? data_i[824] : 1'b0;
  assign data_o[141] = (N1)? data_i[141] : 
                       (N0)? data_i[823] : 1'b0;
  assign data_o[140] = (N1)? data_i[140] : 
                       (N0)? data_i[822] : 1'b0;
  assign data_o[139] = (N1)? data_i[139] : 
                       (N0)? data_i[821] : 1'b0;
  assign data_o[138] = (N1)? data_i[138] : 
                       (N0)? data_i[820] : 1'b0;
  assign data_o[137] = (N1)? data_i[137] : 
                       (N0)? data_i[819] : 1'b0;
  assign data_o[136] = (N1)? data_i[136] : 
                       (N0)? data_i[818] : 1'b0;
  assign data_o[135] = (N1)? data_i[135] : 
                       (N0)? data_i[817] : 1'b0;
  assign data_o[134] = (N1)? data_i[134] : 
                       (N0)? data_i[816] : 1'b0;
  assign data_o[133] = (N1)? data_i[133] : 
                       (N0)? data_i[815] : 1'b0;
  assign data_o[132] = (N1)? data_i[132] : 
                       (N0)? data_i[814] : 1'b0;
  assign data_o[131] = (N1)? data_i[131] : 
                       (N0)? data_i[813] : 1'b0;
  assign data_o[130] = (N1)? data_i[130] : 
                       (N0)? data_i[812] : 1'b0;
  assign data_o[129] = (N1)? data_i[129] : 
                       (N0)? data_i[811] : 1'b0;
  assign data_o[128] = (N1)? data_i[128] : 
                       (N0)? data_i[810] : 1'b0;
  assign data_o[127] = (N1)? data_i[127] : 
                       (N0)? data_i[809] : 1'b0;
  assign data_o[126] = (N1)? data_i[126] : 
                       (N0)? data_i[808] : 1'b0;
  assign data_o[125] = (N1)? data_i[125] : 
                       (N0)? data_i[807] : 1'b0;
  assign data_o[124] = (N1)? data_i[124] : 
                       (N0)? data_i[806] : 1'b0;
  assign data_o[123] = (N1)? data_i[123] : 
                       (N0)? data_i[805] : 1'b0;
  assign data_o[122] = (N1)? data_i[122] : 
                       (N0)? data_i[804] : 1'b0;
  assign data_o[121] = (N1)? data_i[121] : 
                       (N0)? data_i[803] : 1'b0;
  assign data_o[120] = (N1)? data_i[120] : 
                       (N0)? data_i[802] : 1'b0;
  assign data_o[119] = (N1)? data_i[119] : 
                       (N0)? data_i[801] : 1'b0;
  assign data_o[118] = (N1)? data_i[118] : 
                       (N0)? data_i[800] : 1'b0;
  assign data_o[117] = (N1)? data_i[117] : 
                       (N0)? data_i[799] : 1'b0;
  assign data_o[116] = (N1)? data_i[116] : 
                       (N0)? data_i[798] : 1'b0;
  assign data_o[115] = (N1)? data_i[115] : 
                       (N0)? data_i[797] : 1'b0;
  assign data_o[114] = (N1)? data_i[114] : 
                       (N0)? data_i[796] : 1'b0;
  assign data_o[113] = (N1)? data_i[113] : 
                       (N0)? data_i[795] : 1'b0;
  assign data_o[112] = (N1)? data_i[112] : 
                       (N0)? data_i[794] : 1'b0;
  assign data_o[111] = (N1)? data_i[111] : 
                       (N0)? data_i[793] : 1'b0;
  assign data_o[110] = (N1)? data_i[110] : 
                       (N0)? data_i[792] : 1'b0;
  assign data_o[109] = (N1)? data_i[109] : 
                       (N0)? data_i[791] : 1'b0;
  assign data_o[108] = (N1)? data_i[108] : 
                       (N0)? data_i[790] : 1'b0;
  assign data_o[107] = (N1)? data_i[107] : 
                       (N0)? data_i[789] : 1'b0;
  assign data_o[106] = (N1)? data_i[106] : 
                       (N0)? data_i[788] : 1'b0;
  assign data_o[105] = (N1)? data_i[105] : 
                       (N0)? data_i[787] : 1'b0;
  assign data_o[104] = (N1)? data_i[104] : 
                       (N0)? data_i[786] : 1'b0;
  assign data_o[103] = (N1)? data_i[103] : 
                       (N0)? data_i[785] : 1'b0;
  assign data_o[102] = (N1)? data_i[102] : 
                       (N0)? data_i[784] : 1'b0;
  assign data_o[101] = (N1)? data_i[101] : 
                       (N0)? data_i[783] : 1'b0;
  assign data_o[100] = (N1)? data_i[100] : 
                       (N0)? data_i[782] : 1'b0;
  assign data_o[99] = (N1)? data_i[99] : 
                      (N0)? data_i[781] : 1'b0;
  assign data_o[98] = (N1)? data_i[98] : 
                      (N0)? data_i[780] : 1'b0;
  assign data_o[97] = (N1)? data_i[97] : 
                      (N0)? data_i[779] : 1'b0;
  assign data_o[96] = (N1)? data_i[96] : 
                      (N0)? data_i[778] : 1'b0;
  assign data_o[95] = (N1)? data_i[95] : 
                      (N0)? data_i[777] : 1'b0;
  assign data_o[94] = (N1)? data_i[94] : 
                      (N0)? data_i[776] : 1'b0;
  assign data_o[93] = (N1)? data_i[93] : 
                      (N0)? data_i[775] : 1'b0;
  assign data_o[92] = (N1)? data_i[92] : 
                      (N0)? data_i[774] : 1'b0;
  assign data_o[91] = (N1)? data_i[91] : 
                      (N0)? data_i[773] : 1'b0;
  assign data_o[90] = (N1)? data_i[90] : 
                      (N0)? data_i[772] : 1'b0;
  assign data_o[89] = (N1)? data_i[89] : 
                      (N0)? data_i[771] : 1'b0;
  assign data_o[88] = (N1)? data_i[88] : 
                      (N0)? data_i[770] : 1'b0;
  assign data_o[87] = (N1)? data_i[87] : 
                      (N0)? data_i[769] : 1'b0;
  assign data_o[86] = (N1)? data_i[86] : 
                      (N0)? data_i[768] : 1'b0;
  assign data_o[85] = (N1)? data_i[85] : 
                      (N0)? data_i[767] : 1'b0;
  assign data_o[84] = (N1)? data_i[84] : 
                      (N0)? data_i[766] : 1'b0;
  assign data_o[83] = (N1)? data_i[83] : 
                      (N0)? data_i[765] : 1'b0;
  assign data_o[82] = (N1)? data_i[82] : 
                      (N0)? data_i[764] : 1'b0;
  assign data_o[81] = (N1)? data_i[81] : 
                      (N0)? data_i[763] : 1'b0;
  assign data_o[80] = (N1)? data_i[80] : 
                      (N0)? data_i[762] : 1'b0;
  assign data_o[79] = (N1)? data_i[79] : 
                      (N0)? data_i[761] : 1'b0;
  assign data_o[78] = (N1)? data_i[78] : 
                      (N0)? data_i[760] : 1'b0;
  assign data_o[77] = (N1)? data_i[77] : 
                      (N0)? data_i[759] : 1'b0;
  assign data_o[76] = (N1)? data_i[76] : 
                      (N0)? data_i[758] : 1'b0;
  assign data_o[75] = (N1)? data_i[75] : 
                      (N0)? data_i[757] : 1'b0;
  assign data_o[74] = (N1)? data_i[74] : 
                      (N0)? data_i[756] : 1'b0;
  assign data_o[73] = (N1)? data_i[73] : 
                      (N0)? data_i[755] : 1'b0;
  assign data_o[72] = (N1)? data_i[72] : 
                      (N0)? data_i[754] : 1'b0;
  assign data_o[71] = (N1)? data_i[71] : 
                      (N0)? data_i[753] : 1'b0;
  assign data_o[70] = (N1)? data_i[70] : 
                      (N0)? data_i[752] : 1'b0;
  assign data_o[69] = (N1)? data_i[69] : 
                      (N0)? data_i[751] : 1'b0;
  assign data_o[68] = (N1)? data_i[68] : 
                      (N0)? data_i[750] : 1'b0;
  assign data_o[67] = (N1)? data_i[67] : 
                      (N0)? data_i[749] : 1'b0;
  assign data_o[66] = (N1)? data_i[66] : 
                      (N0)? data_i[748] : 1'b0;
  assign data_o[65] = (N1)? data_i[65] : 
                      (N0)? data_i[747] : 1'b0;
  assign data_o[64] = (N1)? data_i[64] : 
                      (N0)? data_i[746] : 1'b0;
  assign data_o[63] = (N1)? data_i[63] : 
                      (N0)? data_i[745] : 1'b0;
  assign data_o[62] = (N1)? data_i[62] : 
                      (N0)? data_i[744] : 1'b0;
  assign data_o[61] = (N1)? data_i[61] : 
                      (N0)? data_i[743] : 1'b0;
  assign data_o[60] = (N1)? data_i[60] : 
                      (N0)? data_i[742] : 1'b0;
  assign data_o[59] = (N1)? data_i[59] : 
                      (N0)? data_i[741] : 1'b0;
  assign data_o[58] = (N1)? data_i[58] : 
                      (N0)? data_i[740] : 1'b0;
  assign data_o[57] = (N1)? data_i[57] : 
                      (N0)? data_i[739] : 1'b0;
  assign data_o[56] = (N1)? data_i[56] : 
                      (N0)? data_i[738] : 1'b0;
  assign data_o[55] = (N1)? data_i[55] : 
                      (N0)? data_i[737] : 1'b0;
  assign data_o[54] = (N1)? data_i[54] : 
                      (N0)? data_i[736] : 1'b0;
  assign data_o[53] = (N1)? data_i[53] : 
                      (N0)? data_i[735] : 1'b0;
  assign data_o[52] = (N1)? data_i[52] : 
                      (N0)? data_i[734] : 1'b0;
  assign data_o[51] = (N1)? data_i[51] : 
                      (N0)? data_i[733] : 1'b0;
  assign data_o[50] = (N1)? data_i[50] : 
                      (N0)? data_i[732] : 1'b0;
  assign data_o[49] = (N1)? data_i[49] : 
                      (N0)? data_i[731] : 1'b0;
  assign data_o[48] = (N1)? data_i[48] : 
                      (N0)? data_i[730] : 1'b0;
  assign data_o[47] = (N1)? data_i[47] : 
                      (N0)? data_i[729] : 1'b0;
  assign data_o[46] = (N1)? data_i[46] : 
                      (N0)? data_i[728] : 1'b0;
  assign data_o[45] = (N1)? data_i[45] : 
                      (N0)? data_i[727] : 1'b0;
  assign data_o[44] = (N1)? data_i[44] : 
                      (N0)? data_i[726] : 1'b0;
  assign data_o[43] = (N1)? data_i[43] : 
                      (N0)? data_i[725] : 1'b0;
  assign data_o[42] = (N1)? data_i[42] : 
                      (N0)? data_i[724] : 1'b0;
  assign data_o[41] = (N1)? data_i[41] : 
                      (N0)? data_i[723] : 1'b0;
  assign data_o[40] = (N1)? data_i[40] : 
                      (N0)? data_i[722] : 1'b0;
  assign data_o[39] = (N1)? data_i[39] : 
                      (N0)? data_i[721] : 1'b0;
  assign data_o[38] = (N1)? data_i[38] : 
                      (N0)? data_i[720] : 1'b0;
  assign data_o[37] = (N1)? data_i[37] : 
                      (N0)? data_i[719] : 1'b0;
  assign data_o[36] = (N1)? data_i[36] : 
                      (N0)? data_i[718] : 1'b0;
  assign data_o[35] = (N1)? data_i[35] : 
                      (N0)? data_i[717] : 1'b0;
  assign data_o[34] = (N1)? data_i[34] : 
                      (N0)? data_i[716] : 1'b0;
  assign data_o[33] = (N1)? data_i[33] : 
                      (N0)? data_i[715] : 1'b0;
  assign data_o[32] = (N1)? data_i[32] : 
                      (N0)? data_i[714] : 1'b0;
  assign data_o[31] = (N1)? data_i[31] : 
                      (N0)? data_i[713] : 1'b0;
  assign data_o[30] = (N1)? data_i[30] : 
                      (N0)? data_i[712] : 1'b0;
  assign data_o[29] = (N1)? data_i[29] : 
                      (N0)? data_i[711] : 1'b0;
  assign data_o[28] = (N1)? data_i[28] : 
                      (N0)? data_i[710] : 1'b0;
  assign data_o[27] = (N1)? data_i[27] : 
                      (N0)? data_i[709] : 1'b0;
  assign data_o[26] = (N1)? data_i[26] : 
                      (N0)? data_i[708] : 1'b0;
  assign data_o[25] = (N1)? data_i[25] : 
                      (N0)? data_i[707] : 1'b0;
  assign data_o[24] = (N1)? data_i[24] : 
                      (N0)? data_i[706] : 1'b0;
  assign data_o[23] = (N1)? data_i[23] : 
                      (N0)? data_i[705] : 1'b0;
  assign data_o[22] = (N1)? data_i[22] : 
                      (N0)? data_i[704] : 1'b0;
  assign data_o[21] = (N1)? data_i[21] : 
                      (N0)? data_i[703] : 1'b0;
  assign data_o[20] = (N1)? data_i[20] : 
                      (N0)? data_i[702] : 1'b0;
  assign data_o[19] = (N1)? data_i[19] : 
                      (N0)? data_i[701] : 1'b0;
  assign data_o[18] = (N1)? data_i[18] : 
                      (N0)? data_i[700] : 1'b0;
  assign data_o[17] = (N1)? data_i[17] : 
                      (N0)? data_i[699] : 1'b0;
  assign data_o[16] = (N1)? data_i[16] : 
                      (N0)? data_i[698] : 1'b0;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[697] : 1'b0;
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[696] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[695] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[694] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[693] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[692] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[691] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[690] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[689] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[688] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[687] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[686] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[685] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[684] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[683] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[682] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_dff_000002ab
(
  clk_i,
  data_i,
  data_o
);

  input [682:0] data_i;
  output [682:0] data_o;
  input clk_i;
  wire [682:0] data_o;
  reg data_o_682_sv2v_reg,data_o_681_sv2v_reg,data_o_680_sv2v_reg,data_o_679_sv2v_reg,
  data_o_678_sv2v_reg,data_o_677_sv2v_reg,data_o_676_sv2v_reg,data_o_675_sv2v_reg,
  data_o_674_sv2v_reg,data_o_673_sv2v_reg,data_o_672_sv2v_reg,data_o_671_sv2v_reg,
  data_o_670_sv2v_reg,data_o_669_sv2v_reg,data_o_668_sv2v_reg,data_o_667_sv2v_reg,
  data_o_666_sv2v_reg,data_o_665_sv2v_reg,data_o_664_sv2v_reg,data_o_663_sv2v_reg,
  data_o_662_sv2v_reg,data_o_661_sv2v_reg,data_o_660_sv2v_reg,data_o_659_sv2v_reg,
  data_o_658_sv2v_reg,data_o_657_sv2v_reg,data_o_656_sv2v_reg,data_o_655_sv2v_reg,
  data_o_654_sv2v_reg,data_o_653_sv2v_reg,data_o_652_sv2v_reg,data_o_651_sv2v_reg,
  data_o_650_sv2v_reg,data_o_649_sv2v_reg,data_o_648_sv2v_reg,data_o_647_sv2v_reg,
  data_o_646_sv2v_reg,data_o_645_sv2v_reg,data_o_644_sv2v_reg,data_o_643_sv2v_reg,
  data_o_642_sv2v_reg,data_o_641_sv2v_reg,data_o_640_sv2v_reg,data_o_639_sv2v_reg,
  data_o_638_sv2v_reg,data_o_637_sv2v_reg,data_o_636_sv2v_reg,data_o_635_sv2v_reg,
  data_o_634_sv2v_reg,data_o_633_sv2v_reg,data_o_632_sv2v_reg,data_o_631_sv2v_reg,
  data_o_630_sv2v_reg,data_o_629_sv2v_reg,data_o_628_sv2v_reg,data_o_627_sv2v_reg,
  data_o_626_sv2v_reg,data_o_625_sv2v_reg,data_o_624_sv2v_reg,data_o_623_sv2v_reg,
  data_o_622_sv2v_reg,data_o_621_sv2v_reg,data_o_620_sv2v_reg,data_o_619_sv2v_reg,
  data_o_618_sv2v_reg,data_o_617_sv2v_reg,data_o_616_sv2v_reg,data_o_615_sv2v_reg,
  data_o_614_sv2v_reg,data_o_613_sv2v_reg,data_o_612_sv2v_reg,data_o_611_sv2v_reg,
  data_o_610_sv2v_reg,data_o_609_sv2v_reg,data_o_608_sv2v_reg,data_o_607_sv2v_reg,
  data_o_606_sv2v_reg,data_o_605_sv2v_reg,data_o_604_sv2v_reg,data_o_603_sv2v_reg,
  data_o_602_sv2v_reg,data_o_601_sv2v_reg,data_o_600_sv2v_reg,data_o_599_sv2v_reg,
  data_o_598_sv2v_reg,data_o_597_sv2v_reg,data_o_596_sv2v_reg,data_o_595_sv2v_reg,
  data_o_594_sv2v_reg,data_o_593_sv2v_reg,data_o_592_sv2v_reg,data_o_591_sv2v_reg,
  data_o_590_sv2v_reg,data_o_589_sv2v_reg,data_o_588_sv2v_reg,data_o_587_sv2v_reg,
  data_o_586_sv2v_reg,data_o_585_sv2v_reg,data_o_584_sv2v_reg,data_o_583_sv2v_reg,
  data_o_582_sv2v_reg,data_o_581_sv2v_reg,data_o_580_sv2v_reg,data_o_579_sv2v_reg,
  data_o_578_sv2v_reg,data_o_577_sv2v_reg,data_o_576_sv2v_reg,data_o_575_sv2v_reg,
  data_o_574_sv2v_reg,data_o_573_sv2v_reg,data_o_572_sv2v_reg,data_o_571_sv2v_reg,
  data_o_570_sv2v_reg,data_o_569_sv2v_reg,data_o_568_sv2v_reg,data_o_567_sv2v_reg,
  data_o_566_sv2v_reg,data_o_565_sv2v_reg,data_o_564_sv2v_reg,data_o_563_sv2v_reg,
  data_o_562_sv2v_reg,data_o_561_sv2v_reg,data_o_560_sv2v_reg,data_o_559_sv2v_reg,
  data_o_558_sv2v_reg,data_o_557_sv2v_reg,data_o_556_sv2v_reg,data_o_555_sv2v_reg,
  data_o_554_sv2v_reg,data_o_553_sv2v_reg,data_o_552_sv2v_reg,data_o_551_sv2v_reg,
  data_o_550_sv2v_reg,data_o_549_sv2v_reg,data_o_548_sv2v_reg,data_o_547_sv2v_reg,
  data_o_546_sv2v_reg,data_o_545_sv2v_reg,data_o_544_sv2v_reg,data_o_543_sv2v_reg,
  data_o_542_sv2v_reg,data_o_541_sv2v_reg,data_o_540_sv2v_reg,data_o_539_sv2v_reg,
  data_o_538_sv2v_reg,data_o_537_sv2v_reg,data_o_536_sv2v_reg,data_o_535_sv2v_reg,
  data_o_534_sv2v_reg,data_o_533_sv2v_reg,data_o_532_sv2v_reg,data_o_531_sv2v_reg,
  data_o_530_sv2v_reg,data_o_529_sv2v_reg,data_o_528_sv2v_reg,data_o_527_sv2v_reg,
  data_o_526_sv2v_reg,data_o_525_sv2v_reg,data_o_524_sv2v_reg,data_o_523_sv2v_reg,
  data_o_522_sv2v_reg,data_o_521_sv2v_reg,data_o_520_sv2v_reg,data_o_519_sv2v_reg,
  data_o_518_sv2v_reg,data_o_517_sv2v_reg,data_o_516_sv2v_reg,data_o_515_sv2v_reg,
  data_o_514_sv2v_reg,data_o_513_sv2v_reg,data_o_512_sv2v_reg,data_o_511_sv2v_reg,
  data_o_510_sv2v_reg,data_o_509_sv2v_reg,data_o_508_sv2v_reg,data_o_507_sv2v_reg,
  data_o_506_sv2v_reg,data_o_505_sv2v_reg,data_o_504_sv2v_reg,data_o_503_sv2v_reg,
  data_o_502_sv2v_reg,data_o_501_sv2v_reg,data_o_500_sv2v_reg,data_o_499_sv2v_reg,
  data_o_498_sv2v_reg,data_o_497_sv2v_reg,data_o_496_sv2v_reg,data_o_495_sv2v_reg,
  data_o_494_sv2v_reg,data_o_493_sv2v_reg,data_o_492_sv2v_reg,data_o_491_sv2v_reg,
  data_o_490_sv2v_reg,data_o_489_sv2v_reg,data_o_488_sv2v_reg,data_o_487_sv2v_reg,
  data_o_486_sv2v_reg,data_o_485_sv2v_reg,data_o_484_sv2v_reg,data_o_483_sv2v_reg,
  data_o_482_sv2v_reg,data_o_481_sv2v_reg,data_o_480_sv2v_reg,data_o_479_sv2v_reg,
  data_o_478_sv2v_reg,data_o_477_sv2v_reg,data_o_476_sv2v_reg,data_o_475_sv2v_reg,
  data_o_474_sv2v_reg,data_o_473_sv2v_reg,data_o_472_sv2v_reg,data_o_471_sv2v_reg,
  data_o_470_sv2v_reg,data_o_469_sv2v_reg,data_o_468_sv2v_reg,data_o_467_sv2v_reg,
  data_o_466_sv2v_reg,data_o_465_sv2v_reg,data_o_464_sv2v_reg,data_o_463_sv2v_reg,
  data_o_462_sv2v_reg,data_o_461_sv2v_reg,data_o_460_sv2v_reg,data_o_459_sv2v_reg,
  data_o_458_sv2v_reg,data_o_457_sv2v_reg,data_o_456_sv2v_reg,data_o_455_sv2v_reg,
  data_o_454_sv2v_reg,data_o_453_sv2v_reg,data_o_452_sv2v_reg,data_o_451_sv2v_reg,
  data_o_450_sv2v_reg,data_o_449_sv2v_reg,data_o_448_sv2v_reg,data_o_447_sv2v_reg,
  data_o_446_sv2v_reg,data_o_445_sv2v_reg,data_o_444_sv2v_reg,data_o_443_sv2v_reg,
  data_o_442_sv2v_reg,data_o_441_sv2v_reg,data_o_440_sv2v_reg,data_o_439_sv2v_reg,
  data_o_438_sv2v_reg,data_o_437_sv2v_reg,data_o_436_sv2v_reg,data_o_435_sv2v_reg,
  data_o_434_sv2v_reg,data_o_433_sv2v_reg,data_o_432_sv2v_reg,data_o_431_sv2v_reg,
  data_o_430_sv2v_reg,data_o_429_sv2v_reg,data_o_428_sv2v_reg,data_o_427_sv2v_reg,
  data_o_426_sv2v_reg,data_o_425_sv2v_reg,data_o_424_sv2v_reg,data_o_423_sv2v_reg,
  data_o_422_sv2v_reg,data_o_421_sv2v_reg,data_o_420_sv2v_reg,data_o_419_sv2v_reg,
  data_o_418_sv2v_reg,data_o_417_sv2v_reg,data_o_416_sv2v_reg,data_o_415_sv2v_reg,
  data_o_414_sv2v_reg,data_o_413_sv2v_reg,data_o_412_sv2v_reg,data_o_411_sv2v_reg,
  data_o_410_sv2v_reg,data_o_409_sv2v_reg,data_o_408_sv2v_reg,data_o_407_sv2v_reg,
  data_o_406_sv2v_reg,data_o_405_sv2v_reg,data_o_404_sv2v_reg,data_o_403_sv2v_reg,
  data_o_402_sv2v_reg,data_o_401_sv2v_reg,data_o_400_sv2v_reg,data_o_399_sv2v_reg,
  data_o_398_sv2v_reg,data_o_397_sv2v_reg,data_o_396_sv2v_reg,data_o_395_sv2v_reg,
  data_o_394_sv2v_reg,data_o_393_sv2v_reg,data_o_392_sv2v_reg,data_o_391_sv2v_reg,
  data_o_390_sv2v_reg,data_o_389_sv2v_reg,data_o_388_sv2v_reg,data_o_387_sv2v_reg,
  data_o_386_sv2v_reg,data_o_385_sv2v_reg,data_o_384_sv2v_reg,data_o_383_sv2v_reg,
  data_o_382_sv2v_reg,data_o_381_sv2v_reg,data_o_380_sv2v_reg,data_o_379_sv2v_reg,
  data_o_378_sv2v_reg,data_o_377_sv2v_reg,data_o_376_sv2v_reg,data_o_375_sv2v_reg,
  data_o_374_sv2v_reg,data_o_373_sv2v_reg,data_o_372_sv2v_reg,data_o_371_sv2v_reg,
  data_o_370_sv2v_reg,data_o_369_sv2v_reg,data_o_368_sv2v_reg,data_o_367_sv2v_reg,
  data_o_366_sv2v_reg,data_o_365_sv2v_reg,data_o_364_sv2v_reg,data_o_363_sv2v_reg,
  data_o_362_sv2v_reg,data_o_361_sv2v_reg,data_o_360_sv2v_reg,data_o_359_sv2v_reg,
  data_o_358_sv2v_reg,data_o_357_sv2v_reg,data_o_356_sv2v_reg,data_o_355_sv2v_reg,
  data_o_354_sv2v_reg,data_o_353_sv2v_reg,data_o_352_sv2v_reg,data_o_351_sv2v_reg,
  data_o_350_sv2v_reg,data_o_349_sv2v_reg,data_o_348_sv2v_reg,data_o_347_sv2v_reg,
  data_o_346_sv2v_reg,data_o_345_sv2v_reg,data_o_344_sv2v_reg,data_o_343_sv2v_reg,
  data_o_342_sv2v_reg,data_o_341_sv2v_reg,data_o_340_sv2v_reg,data_o_339_sv2v_reg,
  data_o_338_sv2v_reg,data_o_337_sv2v_reg,data_o_336_sv2v_reg,data_o_335_sv2v_reg,
  data_o_334_sv2v_reg,data_o_333_sv2v_reg,data_o_332_sv2v_reg,data_o_331_sv2v_reg,
  data_o_330_sv2v_reg,data_o_329_sv2v_reg,data_o_328_sv2v_reg,data_o_327_sv2v_reg,
  data_o_326_sv2v_reg,data_o_325_sv2v_reg,data_o_324_sv2v_reg,data_o_323_sv2v_reg,
  data_o_322_sv2v_reg,data_o_321_sv2v_reg,data_o_320_sv2v_reg,data_o_319_sv2v_reg,
  data_o_318_sv2v_reg,data_o_317_sv2v_reg,data_o_316_sv2v_reg,data_o_315_sv2v_reg,
  data_o_314_sv2v_reg,data_o_313_sv2v_reg,data_o_312_sv2v_reg,data_o_311_sv2v_reg,
  data_o_310_sv2v_reg,data_o_309_sv2v_reg,data_o_308_sv2v_reg,data_o_307_sv2v_reg,
  data_o_306_sv2v_reg,data_o_305_sv2v_reg,data_o_304_sv2v_reg,data_o_303_sv2v_reg,
  data_o_302_sv2v_reg,data_o_301_sv2v_reg,data_o_300_sv2v_reg,data_o_299_sv2v_reg,
  data_o_298_sv2v_reg,data_o_297_sv2v_reg,data_o_296_sv2v_reg,data_o_295_sv2v_reg,
  data_o_294_sv2v_reg,data_o_293_sv2v_reg,data_o_292_sv2v_reg,data_o_291_sv2v_reg,
  data_o_290_sv2v_reg,data_o_289_sv2v_reg,data_o_288_sv2v_reg,data_o_287_sv2v_reg,
  data_o_286_sv2v_reg,data_o_285_sv2v_reg,data_o_284_sv2v_reg,data_o_283_sv2v_reg,
  data_o_282_sv2v_reg,data_o_281_sv2v_reg,data_o_280_sv2v_reg,data_o_279_sv2v_reg,
  data_o_278_sv2v_reg,data_o_277_sv2v_reg,data_o_276_sv2v_reg,data_o_275_sv2v_reg,
  data_o_274_sv2v_reg,data_o_273_sv2v_reg,data_o_272_sv2v_reg,data_o_271_sv2v_reg,
  data_o_270_sv2v_reg,data_o_269_sv2v_reg,data_o_268_sv2v_reg,data_o_267_sv2v_reg,
  data_o_266_sv2v_reg,data_o_265_sv2v_reg,data_o_264_sv2v_reg,data_o_263_sv2v_reg,
  data_o_262_sv2v_reg,data_o_261_sv2v_reg,data_o_260_sv2v_reg,data_o_259_sv2v_reg,
  data_o_258_sv2v_reg,data_o_257_sv2v_reg,data_o_256_sv2v_reg,data_o_255_sv2v_reg,
  data_o_254_sv2v_reg,data_o_253_sv2v_reg,data_o_252_sv2v_reg,data_o_251_sv2v_reg,
  data_o_250_sv2v_reg,data_o_249_sv2v_reg,data_o_248_sv2v_reg,data_o_247_sv2v_reg,
  data_o_246_sv2v_reg,data_o_245_sv2v_reg,data_o_244_sv2v_reg,data_o_243_sv2v_reg,
  data_o_242_sv2v_reg,data_o_241_sv2v_reg,data_o_240_sv2v_reg,data_o_239_sv2v_reg,
  data_o_238_sv2v_reg,data_o_237_sv2v_reg,data_o_236_sv2v_reg,data_o_235_sv2v_reg,
  data_o_234_sv2v_reg,data_o_233_sv2v_reg,data_o_232_sv2v_reg,data_o_231_sv2v_reg,
  data_o_230_sv2v_reg,data_o_229_sv2v_reg,data_o_228_sv2v_reg,data_o_227_sv2v_reg,
  data_o_226_sv2v_reg,data_o_225_sv2v_reg,data_o_224_sv2v_reg,data_o_223_sv2v_reg,
  data_o_222_sv2v_reg,data_o_221_sv2v_reg,data_o_220_sv2v_reg,data_o_219_sv2v_reg,
  data_o_218_sv2v_reg,data_o_217_sv2v_reg,data_o_216_sv2v_reg,data_o_215_sv2v_reg,
  data_o_214_sv2v_reg,data_o_213_sv2v_reg,data_o_212_sv2v_reg,data_o_211_sv2v_reg,
  data_o_210_sv2v_reg,data_o_209_sv2v_reg,data_o_208_sv2v_reg,data_o_207_sv2v_reg,
  data_o_206_sv2v_reg,data_o_205_sv2v_reg,data_o_204_sv2v_reg,data_o_203_sv2v_reg,
  data_o_202_sv2v_reg,data_o_201_sv2v_reg,data_o_200_sv2v_reg,data_o_199_sv2v_reg,
  data_o_198_sv2v_reg,data_o_197_sv2v_reg,data_o_196_sv2v_reg,data_o_195_sv2v_reg,
  data_o_194_sv2v_reg,data_o_193_sv2v_reg,data_o_192_sv2v_reg,data_o_191_sv2v_reg,
  data_o_190_sv2v_reg,data_o_189_sv2v_reg,data_o_188_sv2v_reg,data_o_187_sv2v_reg,
  data_o_186_sv2v_reg,data_o_185_sv2v_reg,data_o_184_sv2v_reg,data_o_183_sv2v_reg,
  data_o_182_sv2v_reg,data_o_181_sv2v_reg,data_o_180_sv2v_reg,data_o_179_sv2v_reg,
  data_o_178_sv2v_reg,data_o_177_sv2v_reg,data_o_176_sv2v_reg,data_o_175_sv2v_reg,
  data_o_174_sv2v_reg,data_o_173_sv2v_reg,data_o_172_sv2v_reg,data_o_171_sv2v_reg,
  data_o_170_sv2v_reg,data_o_169_sv2v_reg,data_o_168_sv2v_reg,data_o_167_sv2v_reg,
  data_o_166_sv2v_reg,data_o_165_sv2v_reg,data_o_164_sv2v_reg,data_o_163_sv2v_reg,
  data_o_162_sv2v_reg,data_o_161_sv2v_reg,data_o_160_sv2v_reg,data_o_159_sv2v_reg,
  data_o_158_sv2v_reg,data_o_157_sv2v_reg,data_o_156_sv2v_reg,data_o_155_sv2v_reg,
  data_o_154_sv2v_reg,data_o_153_sv2v_reg,data_o_152_sv2v_reg,data_o_151_sv2v_reg,
  data_o_150_sv2v_reg,data_o_149_sv2v_reg,data_o_148_sv2v_reg,data_o_147_sv2v_reg,
  data_o_146_sv2v_reg,data_o_145_sv2v_reg,data_o_144_sv2v_reg,data_o_143_sv2v_reg,
  data_o_142_sv2v_reg,data_o_141_sv2v_reg,data_o_140_sv2v_reg,data_o_139_sv2v_reg,
  data_o_138_sv2v_reg,data_o_137_sv2v_reg,data_o_136_sv2v_reg,data_o_135_sv2v_reg,
  data_o_134_sv2v_reg,data_o_133_sv2v_reg,data_o_132_sv2v_reg,data_o_131_sv2v_reg,
  data_o_130_sv2v_reg,data_o_129_sv2v_reg,data_o_128_sv2v_reg,data_o_127_sv2v_reg,
  data_o_126_sv2v_reg,data_o_125_sv2v_reg,data_o_124_sv2v_reg,data_o_123_sv2v_reg,
  data_o_122_sv2v_reg,data_o_121_sv2v_reg,data_o_120_sv2v_reg,data_o_119_sv2v_reg,
  data_o_118_sv2v_reg,data_o_117_sv2v_reg,data_o_116_sv2v_reg,data_o_115_sv2v_reg,
  data_o_114_sv2v_reg,data_o_113_sv2v_reg,data_o_112_sv2v_reg,data_o_111_sv2v_reg,
  data_o_110_sv2v_reg,data_o_109_sv2v_reg,data_o_108_sv2v_reg,data_o_107_sv2v_reg,
  data_o_106_sv2v_reg,data_o_105_sv2v_reg,data_o_104_sv2v_reg,data_o_103_sv2v_reg,
  data_o_102_sv2v_reg,data_o_101_sv2v_reg,data_o_100_sv2v_reg,data_o_99_sv2v_reg,
  data_o_98_sv2v_reg,data_o_97_sv2v_reg,data_o_96_sv2v_reg,data_o_95_sv2v_reg,
  data_o_94_sv2v_reg,data_o_93_sv2v_reg,data_o_92_sv2v_reg,data_o_91_sv2v_reg,
  data_o_90_sv2v_reg,data_o_89_sv2v_reg,data_o_88_sv2v_reg,data_o_87_sv2v_reg,
  data_o_86_sv2v_reg,data_o_85_sv2v_reg,data_o_84_sv2v_reg,data_o_83_sv2v_reg,
  data_o_82_sv2v_reg,data_o_81_sv2v_reg,data_o_80_sv2v_reg,data_o_79_sv2v_reg,data_o_78_sv2v_reg,
  data_o_77_sv2v_reg,data_o_76_sv2v_reg,data_o_75_sv2v_reg,data_o_74_sv2v_reg,
  data_o_73_sv2v_reg,data_o_72_sv2v_reg,data_o_71_sv2v_reg,data_o_70_sv2v_reg,
  data_o_69_sv2v_reg,data_o_68_sv2v_reg,data_o_67_sv2v_reg,data_o_66_sv2v_reg,
  data_o_65_sv2v_reg,data_o_64_sv2v_reg,data_o_63_sv2v_reg,data_o_62_sv2v_reg,
  data_o_61_sv2v_reg,data_o_60_sv2v_reg,data_o_59_sv2v_reg,data_o_58_sv2v_reg,data_o_57_sv2v_reg,
  data_o_56_sv2v_reg,data_o_55_sv2v_reg,data_o_54_sv2v_reg,data_o_53_sv2v_reg,
  data_o_52_sv2v_reg,data_o_51_sv2v_reg,data_o_50_sv2v_reg,data_o_49_sv2v_reg,
  data_o_48_sv2v_reg,data_o_47_sv2v_reg,data_o_46_sv2v_reg,data_o_45_sv2v_reg,
  data_o_44_sv2v_reg,data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,
  data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,
  data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,
  data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,
  data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,
  data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[682] = data_o_682_sv2v_reg;
  assign data_o[681] = data_o_681_sv2v_reg;
  assign data_o[680] = data_o_680_sv2v_reg;
  assign data_o[679] = data_o_679_sv2v_reg;
  assign data_o[678] = data_o_678_sv2v_reg;
  assign data_o[677] = data_o_677_sv2v_reg;
  assign data_o[676] = data_o_676_sv2v_reg;
  assign data_o[675] = data_o_675_sv2v_reg;
  assign data_o[674] = data_o_674_sv2v_reg;
  assign data_o[673] = data_o_673_sv2v_reg;
  assign data_o[672] = data_o_672_sv2v_reg;
  assign data_o[671] = data_o_671_sv2v_reg;
  assign data_o[670] = data_o_670_sv2v_reg;
  assign data_o[669] = data_o_669_sv2v_reg;
  assign data_o[668] = data_o_668_sv2v_reg;
  assign data_o[667] = data_o_667_sv2v_reg;
  assign data_o[666] = data_o_666_sv2v_reg;
  assign data_o[665] = data_o_665_sv2v_reg;
  assign data_o[664] = data_o_664_sv2v_reg;
  assign data_o[663] = data_o_663_sv2v_reg;
  assign data_o[662] = data_o_662_sv2v_reg;
  assign data_o[661] = data_o_661_sv2v_reg;
  assign data_o[660] = data_o_660_sv2v_reg;
  assign data_o[659] = data_o_659_sv2v_reg;
  assign data_o[658] = data_o_658_sv2v_reg;
  assign data_o[657] = data_o_657_sv2v_reg;
  assign data_o[656] = data_o_656_sv2v_reg;
  assign data_o[655] = data_o_655_sv2v_reg;
  assign data_o[654] = data_o_654_sv2v_reg;
  assign data_o[653] = data_o_653_sv2v_reg;
  assign data_o[652] = data_o_652_sv2v_reg;
  assign data_o[651] = data_o_651_sv2v_reg;
  assign data_o[650] = data_o_650_sv2v_reg;
  assign data_o[649] = data_o_649_sv2v_reg;
  assign data_o[648] = data_o_648_sv2v_reg;
  assign data_o[647] = data_o_647_sv2v_reg;
  assign data_o[646] = data_o_646_sv2v_reg;
  assign data_o[645] = data_o_645_sv2v_reg;
  assign data_o[644] = data_o_644_sv2v_reg;
  assign data_o[643] = data_o_643_sv2v_reg;
  assign data_o[642] = data_o_642_sv2v_reg;
  assign data_o[641] = data_o_641_sv2v_reg;
  assign data_o[640] = data_o_640_sv2v_reg;
  assign data_o[639] = data_o_639_sv2v_reg;
  assign data_o[638] = data_o_638_sv2v_reg;
  assign data_o[637] = data_o_637_sv2v_reg;
  assign data_o[636] = data_o_636_sv2v_reg;
  assign data_o[635] = data_o_635_sv2v_reg;
  assign data_o[634] = data_o_634_sv2v_reg;
  assign data_o[633] = data_o_633_sv2v_reg;
  assign data_o[632] = data_o_632_sv2v_reg;
  assign data_o[631] = data_o_631_sv2v_reg;
  assign data_o[630] = data_o_630_sv2v_reg;
  assign data_o[629] = data_o_629_sv2v_reg;
  assign data_o[628] = data_o_628_sv2v_reg;
  assign data_o[627] = data_o_627_sv2v_reg;
  assign data_o[626] = data_o_626_sv2v_reg;
  assign data_o[625] = data_o_625_sv2v_reg;
  assign data_o[624] = data_o_624_sv2v_reg;
  assign data_o[623] = data_o_623_sv2v_reg;
  assign data_o[622] = data_o_622_sv2v_reg;
  assign data_o[621] = data_o_621_sv2v_reg;
  assign data_o[620] = data_o_620_sv2v_reg;
  assign data_o[619] = data_o_619_sv2v_reg;
  assign data_o[618] = data_o_618_sv2v_reg;
  assign data_o[617] = data_o_617_sv2v_reg;
  assign data_o[616] = data_o_616_sv2v_reg;
  assign data_o[615] = data_o_615_sv2v_reg;
  assign data_o[614] = data_o_614_sv2v_reg;
  assign data_o[613] = data_o_613_sv2v_reg;
  assign data_o[612] = data_o_612_sv2v_reg;
  assign data_o[611] = data_o_611_sv2v_reg;
  assign data_o[610] = data_o_610_sv2v_reg;
  assign data_o[609] = data_o_609_sv2v_reg;
  assign data_o[608] = data_o_608_sv2v_reg;
  assign data_o[607] = data_o_607_sv2v_reg;
  assign data_o[606] = data_o_606_sv2v_reg;
  assign data_o[605] = data_o_605_sv2v_reg;
  assign data_o[604] = data_o_604_sv2v_reg;
  assign data_o[603] = data_o_603_sv2v_reg;
  assign data_o[602] = data_o_602_sv2v_reg;
  assign data_o[601] = data_o_601_sv2v_reg;
  assign data_o[600] = data_o_600_sv2v_reg;
  assign data_o[599] = data_o_599_sv2v_reg;
  assign data_o[598] = data_o_598_sv2v_reg;
  assign data_o[597] = data_o_597_sv2v_reg;
  assign data_o[596] = data_o_596_sv2v_reg;
  assign data_o[595] = data_o_595_sv2v_reg;
  assign data_o[594] = data_o_594_sv2v_reg;
  assign data_o[593] = data_o_593_sv2v_reg;
  assign data_o[592] = data_o_592_sv2v_reg;
  assign data_o[591] = data_o_591_sv2v_reg;
  assign data_o[590] = data_o_590_sv2v_reg;
  assign data_o[589] = data_o_589_sv2v_reg;
  assign data_o[588] = data_o_588_sv2v_reg;
  assign data_o[587] = data_o_587_sv2v_reg;
  assign data_o[586] = data_o_586_sv2v_reg;
  assign data_o[585] = data_o_585_sv2v_reg;
  assign data_o[584] = data_o_584_sv2v_reg;
  assign data_o[583] = data_o_583_sv2v_reg;
  assign data_o[582] = data_o_582_sv2v_reg;
  assign data_o[581] = data_o_581_sv2v_reg;
  assign data_o[580] = data_o_580_sv2v_reg;
  assign data_o[579] = data_o_579_sv2v_reg;
  assign data_o[578] = data_o_578_sv2v_reg;
  assign data_o[577] = data_o_577_sv2v_reg;
  assign data_o[576] = data_o_576_sv2v_reg;
  assign data_o[575] = data_o_575_sv2v_reg;
  assign data_o[574] = data_o_574_sv2v_reg;
  assign data_o[573] = data_o_573_sv2v_reg;
  assign data_o[572] = data_o_572_sv2v_reg;
  assign data_o[571] = data_o_571_sv2v_reg;
  assign data_o[570] = data_o_570_sv2v_reg;
  assign data_o[569] = data_o_569_sv2v_reg;
  assign data_o[568] = data_o_568_sv2v_reg;
  assign data_o[567] = data_o_567_sv2v_reg;
  assign data_o[566] = data_o_566_sv2v_reg;
  assign data_o[565] = data_o_565_sv2v_reg;
  assign data_o[564] = data_o_564_sv2v_reg;
  assign data_o[563] = data_o_563_sv2v_reg;
  assign data_o[562] = data_o_562_sv2v_reg;
  assign data_o[561] = data_o_561_sv2v_reg;
  assign data_o[560] = data_o_560_sv2v_reg;
  assign data_o[559] = data_o_559_sv2v_reg;
  assign data_o[558] = data_o_558_sv2v_reg;
  assign data_o[557] = data_o_557_sv2v_reg;
  assign data_o[556] = data_o_556_sv2v_reg;
  assign data_o[555] = data_o_555_sv2v_reg;
  assign data_o[554] = data_o_554_sv2v_reg;
  assign data_o[553] = data_o_553_sv2v_reg;
  assign data_o[552] = data_o_552_sv2v_reg;
  assign data_o[551] = data_o_551_sv2v_reg;
  assign data_o[550] = data_o_550_sv2v_reg;
  assign data_o[549] = data_o_549_sv2v_reg;
  assign data_o[548] = data_o_548_sv2v_reg;
  assign data_o[547] = data_o_547_sv2v_reg;
  assign data_o[546] = data_o_546_sv2v_reg;
  assign data_o[545] = data_o_545_sv2v_reg;
  assign data_o[544] = data_o_544_sv2v_reg;
  assign data_o[543] = data_o_543_sv2v_reg;
  assign data_o[542] = data_o_542_sv2v_reg;
  assign data_o[541] = data_o_541_sv2v_reg;
  assign data_o[540] = data_o_540_sv2v_reg;
  assign data_o[539] = data_o_539_sv2v_reg;
  assign data_o[538] = data_o_538_sv2v_reg;
  assign data_o[537] = data_o_537_sv2v_reg;
  assign data_o[536] = data_o_536_sv2v_reg;
  assign data_o[535] = data_o_535_sv2v_reg;
  assign data_o[534] = data_o_534_sv2v_reg;
  assign data_o[533] = data_o_533_sv2v_reg;
  assign data_o[532] = data_o_532_sv2v_reg;
  assign data_o[531] = data_o_531_sv2v_reg;
  assign data_o[530] = data_o_530_sv2v_reg;
  assign data_o[529] = data_o_529_sv2v_reg;
  assign data_o[528] = data_o_528_sv2v_reg;
  assign data_o[527] = data_o_527_sv2v_reg;
  assign data_o[526] = data_o_526_sv2v_reg;
  assign data_o[525] = data_o_525_sv2v_reg;
  assign data_o[524] = data_o_524_sv2v_reg;
  assign data_o[523] = data_o_523_sv2v_reg;
  assign data_o[522] = data_o_522_sv2v_reg;
  assign data_o[521] = data_o_521_sv2v_reg;
  assign data_o[520] = data_o_520_sv2v_reg;
  assign data_o[519] = data_o_519_sv2v_reg;
  assign data_o[518] = data_o_518_sv2v_reg;
  assign data_o[517] = data_o_517_sv2v_reg;
  assign data_o[516] = data_o_516_sv2v_reg;
  assign data_o[515] = data_o_515_sv2v_reg;
  assign data_o[514] = data_o_514_sv2v_reg;
  assign data_o[513] = data_o_513_sv2v_reg;
  assign data_o[512] = data_o_512_sv2v_reg;
  assign data_o[511] = data_o_511_sv2v_reg;
  assign data_o[510] = data_o_510_sv2v_reg;
  assign data_o[509] = data_o_509_sv2v_reg;
  assign data_o[508] = data_o_508_sv2v_reg;
  assign data_o[507] = data_o_507_sv2v_reg;
  assign data_o[506] = data_o_506_sv2v_reg;
  assign data_o[505] = data_o_505_sv2v_reg;
  assign data_o[504] = data_o_504_sv2v_reg;
  assign data_o[503] = data_o_503_sv2v_reg;
  assign data_o[502] = data_o_502_sv2v_reg;
  assign data_o[501] = data_o_501_sv2v_reg;
  assign data_o[500] = data_o_500_sv2v_reg;
  assign data_o[499] = data_o_499_sv2v_reg;
  assign data_o[498] = data_o_498_sv2v_reg;
  assign data_o[497] = data_o_497_sv2v_reg;
  assign data_o[496] = data_o_496_sv2v_reg;
  assign data_o[495] = data_o_495_sv2v_reg;
  assign data_o[494] = data_o_494_sv2v_reg;
  assign data_o[493] = data_o_493_sv2v_reg;
  assign data_o[492] = data_o_492_sv2v_reg;
  assign data_o[491] = data_o_491_sv2v_reg;
  assign data_o[490] = data_o_490_sv2v_reg;
  assign data_o[489] = data_o_489_sv2v_reg;
  assign data_o[488] = data_o_488_sv2v_reg;
  assign data_o[487] = data_o_487_sv2v_reg;
  assign data_o[486] = data_o_486_sv2v_reg;
  assign data_o[485] = data_o_485_sv2v_reg;
  assign data_o[484] = data_o_484_sv2v_reg;
  assign data_o[483] = data_o_483_sv2v_reg;
  assign data_o[482] = data_o_482_sv2v_reg;
  assign data_o[481] = data_o_481_sv2v_reg;
  assign data_o[480] = data_o_480_sv2v_reg;
  assign data_o[479] = data_o_479_sv2v_reg;
  assign data_o[478] = data_o_478_sv2v_reg;
  assign data_o[477] = data_o_477_sv2v_reg;
  assign data_o[476] = data_o_476_sv2v_reg;
  assign data_o[475] = data_o_475_sv2v_reg;
  assign data_o[474] = data_o_474_sv2v_reg;
  assign data_o[473] = data_o_473_sv2v_reg;
  assign data_o[472] = data_o_472_sv2v_reg;
  assign data_o[471] = data_o_471_sv2v_reg;
  assign data_o[470] = data_o_470_sv2v_reg;
  assign data_o[469] = data_o_469_sv2v_reg;
  assign data_o[468] = data_o_468_sv2v_reg;
  assign data_o[467] = data_o_467_sv2v_reg;
  assign data_o[466] = data_o_466_sv2v_reg;
  assign data_o[465] = data_o_465_sv2v_reg;
  assign data_o[464] = data_o_464_sv2v_reg;
  assign data_o[463] = data_o_463_sv2v_reg;
  assign data_o[462] = data_o_462_sv2v_reg;
  assign data_o[461] = data_o_461_sv2v_reg;
  assign data_o[460] = data_o_460_sv2v_reg;
  assign data_o[459] = data_o_459_sv2v_reg;
  assign data_o[458] = data_o_458_sv2v_reg;
  assign data_o[457] = data_o_457_sv2v_reg;
  assign data_o[456] = data_o_456_sv2v_reg;
  assign data_o[455] = data_o_455_sv2v_reg;
  assign data_o[454] = data_o_454_sv2v_reg;
  assign data_o[453] = data_o_453_sv2v_reg;
  assign data_o[452] = data_o_452_sv2v_reg;
  assign data_o[451] = data_o_451_sv2v_reg;
  assign data_o[450] = data_o_450_sv2v_reg;
  assign data_o[449] = data_o_449_sv2v_reg;
  assign data_o[448] = data_o_448_sv2v_reg;
  assign data_o[447] = data_o_447_sv2v_reg;
  assign data_o[446] = data_o_446_sv2v_reg;
  assign data_o[445] = data_o_445_sv2v_reg;
  assign data_o[444] = data_o_444_sv2v_reg;
  assign data_o[443] = data_o_443_sv2v_reg;
  assign data_o[442] = data_o_442_sv2v_reg;
  assign data_o[441] = data_o_441_sv2v_reg;
  assign data_o[440] = data_o_440_sv2v_reg;
  assign data_o[439] = data_o_439_sv2v_reg;
  assign data_o[438] = data_o_438_sv2v_reg;
  assign data_o[437] = data_o_437_sv2v_reg;
  assign data_o[436] = data_o_436_sv2v_reg;
  assign data_o[435] = data_o_435_sv2v_reg;
  assign data_o[434] = data_o_434_sv2v_reg;
  assign data_o[433] = data_o_433_sv2v_reg;
  assign data_o[432] = data_o_432_sv2v_reg;
  assign data_o[431] = data_o_431_sv2v_reg;
  assign data_o[430] = data_o_430_sv2v_reg;
  assign data_o[429] = data_o_429_sv2v_reg;
  assign data_o[428] = data_o_428_sv2v_reg;
  assign data_o[427] = data_o_427_sv2v_reg;
  assign data_o[426] = data_o_426_sv2v_reg;
  assign data_o[425] = data_o_425_sv2v_reg;
  assign data_o[424] = data_o_424_sv2v_reg;
  assign data_o[423] = data_o_423_sv2v_reg;
  assign data_o[422] = data_o_422_sv2v_reg;
  assign data_o[421] = data_o_421_sv2v_reg;
  assign data_o[420] = data_o_420_sv2v_reg;
  assign data_o[419] = data_o_419_sv2v_reg;
  assign data_o[418] = data_o_418_sv2v_reg;
  assign data_o[417] = data_o_417_sv2v_reg;
  assign data_o[416] = data_o_416_sv2v_reg;
  assign data_o[415] = data_o_415_sv2v_reg;
  assign data_o[414] = data_o_414_sv2v_reg;
  assign data_o[413] = data_o_413_sv2v_reg;
  assign data_o[412] = data_o_412_sv2v_reg;
  assign data_o[411] = data_o_411_sv2v_reg;
  assign data_o[410] = data_o_410_sv2v_reg;
  assign data_o[409] = data_o_409_sv2v_reg;
  assign data_o[408] = data_o_408_sv2v_reg;
  assign data_o[407] = data_o_407_sv2v_reg;
  assign data_o[406] = data_o_406_sv2v_reg;
  assign data_o[405] = data_o_405_sv2v_reg;
  assign data_o[404] = data_o_404_sv2v_reg;
  assign data_o[403] = data_o_403_sv2v_reg;
  assign data_o[402] = data_o_402_sv2v_reg;
  assign data_o[401] = data_o_401_sv2v_reg;
  assign data_o[400] = data_o_400_sv2v_reg;
  assign data_o[399] = data_o_399_sv2v_reg;
  assign data_o[398] = data_o_398_sv2v_reg;
  assign data_o[397] = data_o_397_sv2v_reg;
  assign data_o[396] = data_o_396_sv2v_reg;
  assign data_o[395] = data_o_395_sv2v_reg;
  assign data_o[394] = data_o_394_sv2v_reg;
  assign data_o[393] = data_o_393_sv2v_reg;
  assign data_o[392] = data_o_392_sv2v_reg;
  assign data_o[391] = data_o_391_sv2v_reg;
  assign data_o[390] = data_o_390_sv2v_reg;
  assign data_o[389] = data_o_389_sv2v_reg;
  assign data_o[388] = data_o_388_sv2v_reg;
  assign data_o[387] = data_o_387_sv2v_reg;
  assign data_o[386] = data_o_386_sv2v_reg;
  assign data_o[385] = data_o_385_sv2v_reg;
  assign data_o[384] = data_o_384_sv2v_reg;
  assign data_o[383] = data_o_383_sv2v_reg;
  assign data_o[382] = data_o_382_sv2v_reg;
  assign data_o[381] = data_o_381_sv2v_reg;
  assign data_o[380] = data_o_380_sv2v_reg;
  assign data_o[379] = data_o_379_sv2v_reg;
  assign data_o[378] = data_o_378_sv2v_reg;
  assign data_o[377] = data_o_377_sv2v_reg;
  assign data_o[376] = data_o_376_sv2v_reg;
  assign data_o[375] = data_o_375_sv2v_reg;
  assign data_o[374] = data_o_374_sv2v_reg;
  assign data_o[373] = data_o_373_sv2v_reg;
  assign data_o[372] = data_o_372_sv2v_reg;
  assign data_o[371] = data_o_371_sv2v_reg;
  assign data_o[370] = data_o_370_sv2v_reg;
  assign data_o[369] = data_o_369_sv2v_reg;
  assign data_o[368] = data_o_368_sv2v_reg;
  assign data_o[367] = data_o_367_sv2v_reg;
  assign data_o[366] = data_o_366_sv2v_reg;
  assign data_o[365] = data_o_365_sv2v_reg;
  assign data_o[364] = data_o_364_sv2v_reg;
  assign data_o[363] = data_o_363_sv2v_reg;
  assign data_o[362] = data_o_362_sv2v_reg;
  assign data_o[361] = data_o_361_sv2v_reg;
  assign data_o[360] = data_o_360_sv2v_reg;
  assign data_o[359] = data_o_359_sv2v_reg;
  assign data_o[358] = data_o_358_sv2v_reg;
  assign data_o[357] = data_o_357_sv2v_reg;
  assign data_o[356] = data_o_356_sv2v_reg;
  assign data_o[355] = data_o_355_sv2v_reg;
  assign data_o[354] = data_o_354_sv2v_reg;
  assign data_o[353] = data_o_353_sv2v_reg;
  assign data_o[352] = data_o_352_sv2v_reg;
  assign data_o[351] = data_o_351_sv2v_reg;
  assign data_o[350] = data_o_350_sv2v_reg;
  assign data_o[349] = data_o_349_sv2v_reg;
  assign data_o[348] = data_o_348_sv2v_reg;
  assign data_o[347] = data_o_347_sv2v_reg;
  assign data_o[346] = data_o_346_sv2v_reg;
  assign data_o[345] = data_o_345_sv2v_reg;
  assign data_o[344] = data_o_344_sv2v_reg;
  assign data_o[343] = data_o_343_sv2v_reg;
  assign data_o[342] = data_o_342_sv2v_reg;
  assign data_o[341] = data_o_341_sv2v_reg;
  assign data_o[340] = data_o_340_sv2v_reg;
  assign data_o[339] = data_o_339_sv2v_reg;
  assign data_o[338] = data_o_338_sv2v_reg;
  assign data_o[337] = data_o_337_sv2v_reg;
  assign data_o[336] = data_o_336_sv2v_reg;
  assign data_o[335] = data_o_335_sv2v_reg;
  assign data_o[334] = data_o_334_sv2v_reg;
  assign data_o[333] = data_o_333_sv2v_reg;
  assign data_o[332] = data_o_332_sv2v_reg;
  assign data_o[331] = data_o_331_sv2v_reg;
  assign data_o[330] = data_o_330_sv2v_reg;
  assign data_o[329] = data_o_329_sv2v_reg;
  assign data_o[328] = data_o_328_sv2v_reg;
  assign data_o[327] = data_o_327_sv2v_reg;
  assign data_o[326] = data_o_326_sv2v_reg;
  assign data_o[325] = data_o_325_sv2v_reg;
  assign data_o[324] = data_o_324_sv2v_reg;
  assign data_o[323] = data_o_323_sv2v_reg;
  assign data_o[322] = data_o_322_sv2v_reg;
  assign data_o[321] = data_o_321_sv2v_reg;
  assign data_o[320] = data_o_320_sv2v_reg;
  assign data_o[319] = data_o_319_sv2v_reg;
  assign data_o[318] = data_o_318_sv2v_reg;
  assign data_o[317] = data_o_317_sv2v_reg;
  assign data_o[316] = data_o_316_sv2v_reg;
  assign data_o[315] = data_o_315_sv2v_reg;
  assign data_o[314] = data_o_314_sv2v_reg;
  assign data_o[313] = data_o_313_sv2v_reg;
  assign data_o[312] = data_o_312_sv2v_reg;
  assign data_o[311] = data_o_311_sv2v_reg;
  assign data_o[310] = data_o_310_sv2v_reg;
  assign data_o[309] = data_o_309_sv2v_reg;
  assign data_o[308] = data_o_308_sv2v_reg;
  assign data_o[307] = data_o_307_sv2v_reg;
  assign data_o[306] = data_o_306_sv2v_reg;
  assign data_o[305] = data_o_305_sv2v_reg;
  assign data_o[304] = data_o_304_sv2v_reg;
  assign data_o[303] = data_o_303_sv2v_reg;
  assign data_o[302] = data_o_302_sv2v_reg;
  assign data_o[301] = data_o_301_sv2v_reg;
  assign data_o[300] = data_o_300_sv2v_reg;
  assign data_o[299] = data_o_299_sv2v_reg;
  assign data_o[298] = data_o_298_sv2v_reg;
  assign data_o[297] = data_o_297_sv2v_reg;
  assign data_o[296] = data_o_296_sv2v_reg;
  assign data_o[295] = data_o_295_sv2v_reg;
  assign data_o[294] = data_o_294_sv2v_reg;
  assign data_o[293] = data_o_293_sv2v_reg;
  assign data_o[292] = data_o_292_sv2v_reg;
  assign data_o[291] = data_o_291_sv2v_reg;
  assign data_o[290] = data_o_290_sv2v_reg;
  assign data_o[289] = data_o_289_sv2v_reg;
  assign data_o[288] = data_o_288_sv2v_reg;
  assign data_o[287] = data_o_287_sv2v_reg;
  assign data_o[286] = data_o_286_sv2v_reg;
  assign data_o[285] = data_o_285_sv2v_reg;
  assign data_o[284] = data_o_284_sv2v_reg;
  assign data_o[283] = data_o_283_sv2v_reg;
  assign data_o[282] = data_o_282_sv2v_reg;
  assign data_o[281] = data_o_281_sv2v_reg;
  assign data_o[280] = data_o_280_sv2v_reg;
  assign data_o[279] = data_o_279_sv2v_reg;
  assign data_o[278] = data_o_278_sv2v_reg;
  assign data_o[277] = data_o_277_sv2v_reg;
  assign data_o[276] = data_o_276_sv2v_reg;
  assign data_o[275] = data_o_275_sv2v_reg;
  assign data_o[274] = data_o_274_sv2v_reg;
  assign data_o[273] = data_o_273_sv2v_reg;
  assign data_o[272] = data_o_272_sv2v_reg;
  assign data_o[271] = data_o_271_sv2v_reg;
  assign data_o[270] = data_o_270_sv2v_reg;
  assign data_o[269] = data_o_269_sv2v_reg;
  assign data_o[268] = data_o_268_sv2v_reg;
  assign data_o[267] = data_o_267_sv2v_reg;
  assign data_o[266] = data_o_266_sv2v_reg;
  assign data_o[265] = data_o_265_sv2v_reg;
  assign data_o[264] = data_o_264_sv2v_reg;
  assign data_o[263] = data_o_263_sv2v_reg;
  assign data_o[262] = data_o_262_sv2v_reg;
  assign data_o[261] = data_o_261_sv2v_reg;
  assign data_o[260] = data_o_260_sv2v_reg;
  assign data_o[259] = data_o_259_sv2v_reg;
  assign data_o[258] = data_o_258_sv2v_reg;
  assign data_o[257] = data_o_257_sv2v_reg;
  assign data_o[256] = data_o_256_sv2v_reg;
  assign data_o[255] = data_o_255_sv2v_reg;
  assign data_o[254] = data_o_254_sv2v_reg;
  assign data_o[253] = data_o_253_sv2v_reg;
  assign data_o[252] = data_o_252_sv2v_reg;
  assign data_o[251] = data_o_251_sv2v_reg;
  assign data_o[250] = data_o_250_sv2v_reg;
  assign data_o[249] = data_o_249_sv2v_reg;
  assign data_o[248] = data_o_248_sv2v_reg;
  assign data_o[247] = data_o_247_sv2v_reg;
  assign data_o[246] = data_o_246_sv2v_reg;
  assign data_o[245] = data_o_245_sv2v_reg;
  assign data_o[244] = data_o_244_sv2v_reg;
  assign data_o[243] = data_o_243_sv2v_reg;
  assign data_o[242] = data_o_242_sv2v_reg;
  assign data_o[241] = data_o_241_sv2v_reg;
  assign data_o[240] = data_o_240_sv2v_reg;
  assign data_o[239] = data_o_239_sv2v_reg;
  assign data_o[238] = data_o_238_sv2v_reg;
  assign data_o[237] = data_o_237_sv2v_reg;
  assign data_o[236] = data_o_236_sv2v_reg;
  assign data_o[235] = data_o_235_sv2v_reg;
  assign data_o[234] = data_o_234_sv2v_reg;
  assign data_o[233] = data_o_233_sv2v_reg;
  assign data_o[232] = data_o_232_sv2v_reg;
  assign data_o[231] = data_o_231_sv2v_reg;
  assign data_o[230] = data_o_230_sv2v_reg;
  assign data_o[229] = data_o_229_sv2v_reg;
  assign data_o[228] = data_o_228_sv2v_reg;
  assign data_o[227] = data_o_227_sv2v_reg;
  assign data_o[226] = data_o_226_sv2v_reg;
  assign data_o[225] = data_o_225_sv2v_reg;
  assign data_o[224] = data_o_224_sv2v_reg;
  assign data_o[223] = data_o_223_sv2v_reg;
  assign data_o[222] = data_o_222_sv2v_reg;
  assign data_o[221] = data_o_221_sv2v_reg;
  assign data_o[220] = data_o_220_sv2v_reg;
  assign data_o[219] = data_o_219_sv2v_reg;
  assign data_o[218] = data_o_218_sv2v_reg;
  assign data_o[217] = data_o_217_sv2v_reg;
  assign data_o[216] = data_o_216_sv2v_reg;
  assign data_o[215] = data_o_215_sv2v_reg;
  assign data_o[214] = data_o_214_sv2v_reg;
  assign data_o[213] = data_o_213_sv2v_reg;
  assign data_o[212] = data_o_212_sv2v_reg;
  assign data_o[211] = data_o_211_sv2v_reg;
  assign data_o[210] = data_o_210_sv2v_reg;
  assign data_o[209] = data_o_209_sv2v_reg;
  assign data_o[208] = data_o_208_sv2v_reg;
  assign data_o[207] = data_o_207_sv2v_reg;
  assign data_o[206] = data_o_206_sv2v_reg;
  assign data_o[205] = data_o_205_sv2v_reg;
  assign data_o[204] = data_o_204_sv2v_reg;
  assign data_o[203] = data_o_203_sv2v_reg;
  assign data_o[202] = data_o_202_sv2v_reg;
  assign data_o[201] = data_o_201_sv2v_reg;
  assign data_o[200] = data_o_200_sv2v_reg;
  assign data_o[199] = data_o_199_sv2v_reg;
  assign data_o[198] = data_o_198_sv2v_reg;
  assign data_o[197] = data_o_197_sv2v_reg;
  assign data_o[196] = data_o_196_sv2v_reg;
  assign data_o[195] = data_o_195_sv2v_reg;
  assign data_o[194] = data_o_194_sv2v_reg;
  assign data_o[193] = data_o_193_sv2v_reg;
  assign data_o[192] = data_o_192_sv2v_reg;
  assign data_o[191] = data_o_191_sv2v_reg;
  assign data_o[190] = data_o_190_sv2v_reg;
  assign data_o[189] = data_o_189_sv2v_reg;
  assign data_o[188] = data_o_188_sv2v_reg;
  assign data_o[187] = data_o_187_sv2v_reg;
  assign data_o[186] = data_o_186_sv2v_reg;
  assign data_o[185] = data_o_185_sv2v_reg;
  assign data_o[184] = data_o_184_sv2v_reg;
  assign data_o[183] = data_o_183_sv2v_reg;
  assign data_o[182] = data_o_182_sv2v_reg;
  assign data_o[181] = data_o_181_sv2v_reg;
  assign data_o[180] = data_o_180_sv2v_reg;
  assign data_o[179] = data_o_179_sv2v_reg;
  assign data_o[178] = data_o_178_sv2v_reg;
  assign data_o[177] = data_o_177_sv2v_reg;
  assign data_o[176] = data_o_176_sv2v_reg;
  assign data_o[175] = data_o_175_sv2v_reg;
  assign data_o[174] = data_o_174_sv2v_reg;
  assign data_o[173] = data_o_173_sv2v_reg;
  assign data_o[172] = data_o_172_sv2v_reg;
  assign data_o[171] = data_o_171_sv2v_reg;
  assign data_o[170] = data_o_170_sv2v_reg;
  assign data_o[169] = data_o_169_sv2v_reg;
  assign data_o[168] = data_o_168_sv2v_reg;
  assign data_o[167] = data_o_167_sv2v_reg;
  assign data_o[166] = data_o_166_sv2v_reg;
  assign data_o[165] = data_o_165_sv2v_reg;
  assign data_o[164] = data_o_164_sv2v_reg;
  assign data_o[163] = data_o_163_sv2v_reg;
  assign data_o[162] = data_o_162_sv2v_reg;
  assign data_o[161] = data_o_161_sv2v_reg;
  assign data_o[160] = data_o_160_sv2v_reg;
  assign data_o[159] = data_o_159_sv2v_reg;
  assign data_o[158] = data_o_158_sv2v_reg;
  assign data_o[157] = data_o_157_sv2v_reg;
  assign data_o[156] = data_o_156_sv2v_reg;
  assign data_o[155] = data_o_155_sv2v_reg;
  assign data_o[154] = data_o_154_sv2v_reg;
  assign data_o[153] = data_o_153_sv2v_reg;
  assign data_o[152] = data_o_152_sv2v_reg;
  assign data_o[151] = data_o_151_sv2v_reg;
  assign data_o[150] = data_o_150_sv2v_reg;
  assign data_o[149] = data_o_149_sv2v_reg;
  assign data_o[148] = data_o_148_sv2v_reg;
  assign data_o[147] = data_o_147_sv2v_reg;
  assign data_o[146] = data_o_146_sv2v_reg;
  assign data_o[145] = data_o_145_sv2v_reg;
  assign data_o[144] = data_o_144_sv2v_reg;
  assign data_o[143] = data_o_143_sv2v_reg;
  assign data_o[142] = data_o_142_sv2v_reg;
  assign data_o[141] = data_o_141_sv2v_reg;
  assign data_o[140] = data_o_140_sv2v_reg;
  assign data_o[139] = data_o_139_sv2v_reg;
  assign data_o[138] = data_o_138_sv2v_reg;
  assign data_o[137] = data_o_137_sv2v_reg;
  assign data_o[136] = data_o_136_sv2v_reg;
  assign data_o[135] = data_o_135_sv2v_reg;
  assign data_o[134] = data_o_134_sv2v_reg;
  assign data_o[133] = data_o_133_sv2v_reg;
  assign data_o[132] = data_o_132_sv2v_reg;
  assign data_o[131] = data_o_131_sv2v_reg;
  assign data_o[130] = data_o_130_sv2v_reg;
  assign data_o[129] = data_o_129_sv2v_reg;
  assign data_o[128] = data_o_128_sv2v_reg;
  assign data_o[127] = data_o_127_sv2v_reg;
  assign data_o[126] = data_o_126_sv2v_reg;
  assign data_o[125] = data_o_125_sv2v_reg;
  assign data_o[124] = data_o_124_sv2v_reg;
  assign data_o[123] = data_o_123_sv2v_reg;
  assign data_o[122] = data_o_122_sv2v_reg;
  assign data_o[121] = data_o_121_sv2v_reg;
  assign data_o[120] = data_o_120_sv2v_reg;
  assign data_o[119] = data_o_119_sv2v_reg;
  assign data_o[118] = data_o_118_sv2v_reg;
  assign data_o[117] = data_o_117_sv2v_reg;
  assign data_o[116] = data_o_116_sv2v_reg;
  assign data_o[115] = data_o_115_sv2v_reg;
  assign data_o[114] = data_o_114_sv2v_reg;
  assign data_o[113] = data_o_113_sv2v_reg;
  assign data_o[112] = data_o_112_sv2v_reg;
  assign data_o[111] = data_o_111_sv2v_reg;
  assign data_o[110] = data_o_110_sv2v_reg;
  assign data_o[109] = data_o_109_sv2v_reg;
  assign data_o[108] = data_o_108_sv2v_reg;
  assign data_o[107] = data_o_107_sv2v_reg;
  assign data_o[106] = data_o_106_sv2v_reg;
  assign data_o[105] = data_o_105_sv2v_reg;
  assign data_o[104] = data_o_104_sv2v_reg;
  assign data_o[103] = data_o_103_sv2v_reg;
  assign data_o[102] = data_o_102_sv2v_reg;
  assign data_o[101] = data_o_101_sv2v_reg;
  assign data_o[100] = data_o_100_sv2v_reg;
  assign data_o[99] = data_o_99_sv2v_reg;
  assign data_o[98] = data_o_98_sv2v_reg;
  assign data_o[97] = data_o_97_sv2v_reg;
  assign data_o[96] = data_o_96_sv2v_reg;
  assign data_o[95] = data_o_95_sv2v_reg;
  assign data_o[94] = data_o_94_sv2v_reg;
  assign data_o[93] = data_o_93_sv2v_reg;
  assign data_o[92] = data_o_92_sv2v_reg;
  assign data_o[91] = data_o_91_sv2v_reg;
  assign data_o[90] = data_o_90_sv2v_reg;
  assign data_o[89] = data_o_89_sv2v_reg;
  assign data_o[88] = data_o_88_sv2v_reg;
  assign data_o[87] = data_o_87_sv2v_reg;
  assign data_o[86] = data_o_86_sv2v_reg;
  assign data_o[85] = data_o_85_sv2v_reg;
  assign data_o[84] = data_o_84_sv2v_reg;
  assign data_o[83] = data_o_83_sv2v_reg;
  assign data_o[82] = data_o_82_sv2v_reg;
  assign data_o[81] = data_o_81_sv2v_reg;
  assign data_o[80] = data_o_80_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_682_sv2v_reg <= data_i[682];
      data_o_681_sv2v_reg <= data_i[681];
      data_o_680_sv2v_reg <= data_i[680];
      data_o_679_sv2v_reg <= data_i[679];
      data_o_678_sv2v_reg <= data_i[678];
      data_o_677_sv2v_reg <= data_i[677];
      data_o_676_sv2v_reg <= data_i[676];
      data_o_675_sv2v_reg <= data_i[675];
      data_o_674_sv2v_reg <= data_i[674];
      data_o_673_sv2v_reg <= data_i[673];
      data_o_672_sv2v_reg <= data_i[672];
      data_o_671_sv2v_reg <= data_i[671];
      data_o_670_sv2v_reg <= data_i[670];
      data_o_669_sv2v_reg <= data_i[669];
      data_o_668_sv2v_reg <= data_i[668];
      data_o_667_sv2v_reg <= data_i[667];
      data_o_666_sv2v_reg <= data_i[666];
      data_o_665_sv2v_reg <= data_i[665];
      data_o_664_sv2v_reg <= data_i[664];
      data_o_663_sv2v_reg <= data_i[663];
      data_o_662_sv2v_reg <= data_i[662];
      data_o_661_sv2v_reg <= data_i[661];
      data_o_660_sv2v_reg <= data_i[660];
      data_o_659_sv2v_reg <= data_i[659];
      data_o_658_sv2v_reg <= data_i[658];
      data_o_657_sv2v_reg <= data_i[657];
      data_o_656_sv2v_reg <= data_i[656];
      data_o_655_sv2v_reg <= data_i[655];
      data_o_654_sv2v_reg <= data_i[654];
      data_o_653_sv2v_reg <= data_i[653];
      data_o_652_sv2v_reg <= data_i[652];
      data_o_651_sv2v_reg <= data_i[651];
      data_o_650_sv2v_reg <= data_i[650];
      data_o_649_sv2v_reg <= data_i[649];
      data_o_648_sv2v_reg <= data_i[648];
      data_o_647_sv2v_reg <= data_i[647];
      data_o_646_sv2v_reg <= data_i[646];
      data_o_645_sv2v_reg <= data_i[645];
      data_o_644_sv2v_reg <= data_i[644];
      data_o_643_sv2v_reg <= data_i[643];
      data_o_642_sv2v_reg <= data_i[642];
      data_o_641_sv2v_reg <= data_i[641];
      data_o_640_sv2v_reg <= data_i[640];
      data_o_639_sv2v_reg <= data_i[639];
      data_o_638_sv2v_reg <= data_i[638];
      data_o_637_sv2v_reg <= data_i[637];
      data_o_636_sv2v_reg <= data_i[636];
      data_o_635_sv2v_reg <= data_i[635];
      data_o_634_sv2v_reg <= data_i[634];
      data_o_633_sv2v_reg <= data_i[633];
      data_o_632_sv2v_reg <= data_i[632];
      data_o_631_sv2v_reg <= data_i[631];
      data_o_630_sv2v_reg <= data_i[630];
      data_o_629_sv2v_reg <= data_i[629];
      data_o_628_sv2v_reg <= data_i[628];
      data_o_627_sv2v_reg <= data_i[627];
      data_o_626_sv2v_reg <= data_i[626];
      data_o_625_sv2v_reg <= data_i[625];
      data_o_624_sv2v_reg <= data_i[624];
      data_o_623_sv2v_reg <= data_i[623];
      data_o_622_sv2v_reg <= data_i[622];
      data_o_621_sv2v_reg <= data_i[621];
      data_o_620_sv2v_reg <= data_i[620];
      data_o_619_sv2v_reg <= data_i[619];
      data_o_618_sv2v_reg <= data_i[618];
      data_o_617_sv2v_reg <= data_i[617];
      data_o_616_sv2v_reg <= data_i[616];
      data_o_615_sv2v_reg <= data_i[615];
      data_o_614_sv2v_reg <= data_i[614];
      data_o_613_sv2v_reg <= data_i[613];
      data_o_612_sv2v_reg <= data_i[612];
      data_o_611_sv2v_reg <= data_i[611];
      data_o_610_sv2v_reg <= data_i[610];
      data_o_609_sv2v_reg <= data_i[609];
      data_o_608_sv2v_reg <= data_i[608];
      data_o_607_sv2v_reg <= data_i[607];
      data_o_606_sv2v_reg <= data_i[606];
      data_o_605_sv2v_reg <= data_i[605];
      data_o_604_sv2v_reg <= data_i[604];
      data_o_603_sv2v_reg <= data_i[603];
      data_o_602_sv2v_reg <= data_i[602];
      data_o_601_sv2v_reg <= data_i[601];
      data_o_600_sv2v_reg <= data_i[600];
      data_o_599_sv2v_reg <= data_i[599];
      data_o_598_sv2v_reg <= data_i[598];
      data_o_597_sv2v_reg <= data_i[597];
      data_o_596_sv2v_reg <= data_i[596];
      data_o_595_sv2v_reg <= data_i[595];
      data_o_594_sv2v_reg <= data_i[594];
      data_o_593_sv2v_reg <= data_i[593];
      data_o_592_sv2v_reg <= data_i[592];
      data_o_591_sv2v_reg <= data_i[591];
      data_o_590_sv2v_reg <= data_i[590];
      data_o_589_sv2v_reg <= data_i[589];
      data_o_588_sv2v_reg <= data_i[588];
      data_o_587_sv2v_reg <= data_i[587];
      data_o_586_sv2v_reg <= data_i[586];
      data_o_585_sv2v_reg <= data_i[585];
      data_o_584_sv2v_reg <= data_i[584];
      data_o_583_sv2v_reg <= data_i[583];
      data_o_582_sv2v_reg <= data_i[582];
      data_o_581_sv2v_reg <= data_i[581];
      data_o_580_sv2v_reg <= data_i[580];
      data_o_579_sv2v_reg <= data_i[579];
      data_o_578_sv2v_reg <= data_i[578];
      data_o_577_sv2v_reg <= data_i[577];
      data_o_576_sv2v_reg <= data_i[576];
      data_o_575_sv2v_reg <= data_i[575];
      data_o_574_sv2v_reg <= data_i[574];
      data_o_573_sv2v_reg <= data_i[573];
      data_o_572_sv2v_reg <= data_i[572];
      data_o_571_sv2v_reg <= data_i[571];
      data_o_570_sv2v_reg <= data_i[570];
      data_o_569_sv2v_reg <= data_i[569];
      data_o_568_sv2v_reg <= data_i[568];
      data_o_567_sv2v_reg <= data_i[567];
      data_o_566_sv2v_reg <= data_i[566];
      data_o_565_sv2v_reg <= data_i[565];
      data_o_564_sv2v_reg <= data_i[564];
      data_o_563_sv2v_reg <= data_i[563];
      data_o_562_sv2v_reg <= data_i[562];
      data_o_561_sv2v_reg <= data_i[561];
      data_o_560_sv2v_reg <= data_i[560];
      data_o_559_sv2v_reg <= data_i[559];
      data_o_558_sv2v_reg <= data_i[558];
      data_o_557_sv2v_reg <= data_i[557];
      data_o_556_sv2v_reg <= data_i[556];
      data_o_555_sv2v_reg <= data_i[555];
      data_o_554_sv2v_reg <= data_i[554];
      data_o_553_sv2v_reg <= data_i[553];
      data_o_552_sv2v_reg <= data_i[552];
      data_o_551_sv2v_reg <= data_i[551];
      data_o_550_sv2v_reg <= data_i[550];
      data_o_549_sv2v_reg <= data_i[549];
      data_o_548_sv2v_reg <= data_i[548];
      data_o_547_sv2v_reg <= data_i[547];
      data_o_546_sv2v_reg <= data_i[546];
      data_o_545_sv2v_reg <= data_i[545];
      data_o_544_sv2v_reg <= data_i[544];
      data_o_543_sv2v_reg <= data_i[543];
      data_o_542_sv2v_reg <= data_i[542];
      data_o_541_sv2v_reg <= data_i[541];
      data_o_540_sv2v_reg <= data_i[540];
      data_o_539_sv2v_reg <= data_i[539];
      data_o_538_sv2v_reg <= data_i[538];
      data_o_537_sv2v_reg <= data_i[537];
      data_o_536_sv2v_reg <= data_i[536];
      data_o_535_sv2v_reg <= data_i[535];
      data_o_534_sv2v_reg <= data_i[534];
      data_o_533_sv2v_reg <= data_i[533];
      data_o_532_sv2v_reg <= data_i[532];
      data_o_531_sv2v_reg <= data_i[531];
      data_o_530_sv2v_reg <= data_i[530];
      data_o_529_sv2v_reg <= data_i[529];
      data_o_528_sv2v_reg <= data_i[528];
      data_o_527_sv2v_reg <= data_i[527];
      data_o_526_sv2v_reg <= data_i[526];
      data_o_525_sv2v_reg <= data_i[525];
      data_o_524_sv2v_reg <= data_i[524];
      data_o_523_sv2v_reg <= data_i[523];
      data_o_522_sv2v_reg <= data_i[522];
      data_o_521_sv2v_reg <= data_i[521];
      data_o_520_sv2v_reg <= data_i[520];
      data_o_519_sv2v_reg <= data_i[519];
      data_o_518_sv2v_reg <= data_i[518];
      data_o_517_sv2v_reg <= data_i[517];
      data_o_516_sv2v_reg <= data_i[516];
      data_o_515_sv2v_reg <= data_i[515];
      data_o_514_sv2v_reg <= data_i[514];
      data_o_513_sv2v_reg <= data_i[513];
      data_o_512_sv2v_reg <= data_i[512];
      data_o_511_sv2v_reg <= data_i[511];
      data_o_510_sv2v_reg <= data_i[510];
      data_o_509_sv2v_reg <= data_i[509];
      data_o_508_sv2v_reg <= data_i[508];
      data_o_507_sv2v_reg <= data_i[507];
      data_o_506_sv2v_reg <= data_i[506];
      data_o_505_sv2v_reg <= data_i[505];
      data_o_504_sv2v_reg <= data_i[504];
      data_o_503_sv2v_reg <= data_i[503];
      data_o_502_sv2v_reg <= data_i[502];
      data_o_501_sv2v_reg <= data_i[501];
      data_o_500_sv2v_reg <= data_i[500];
      data_o_499_sv2v_reg <= data_i[499];
      data_o_498_sv2v_reg <= data_i[498];
      data_o_497_sv2v_reg <= data_i[497];
      data_o_496_sv2v_reg <= data_i[496];
      data_o_495_sv2v_reg <= data_i[495];
      data_o_494_sv2v_reg <= data_i[494];
      data_o_493_sv2v_reg <= data_i[493];
      data_o_492_sv2v_reg <= data_i[492];
      data_o_491_sv2v_reg <= data_i[491];
      data_o_490_sv2v_reg <= data_i[490];
      data_o_489_sv2v_reg <= data_i[489];
      data_o_488_sv2v_reg <= data_i[488];
      data_o_487_sv2v_reg <= data_i[487];
      data_o_486_sv2v_reg <= data_i[486];
      data_o_485_sv2v_reg <= data_i[485];
      data_o_484_sv2v_reg <= data_i[484];
      data_o_483_sv2v_reg <= data_i[483];
      data_o_482_sv2v_reg <= data_i[482];
      data_o_481_sv2v_reg <= data_i[481];
      data_o_480_sv2v_reg <= data_i[480];
      data_o_479_sv2v_reg <= data_i[479];
      data_o_478_sv2v_reg <= data_i[478];
      data_o_477_sv2v_reg <= data_i[477];
      data_o_476_sv2v_reg <= data_i[476];
      data_o_475_sv2v_reg <= data_i[475];
      data_o_474_sv2v_reg <= data_i[474];
      data_o_473_sv2v_reg <= data_i[473];
      data_o_472_sv2v_reg <= data_i[472];
      data_o_471_sv2v_reg <= data_i[471];
      data_o_470_sv2v_reg <= data_i[470];
      data_o_469_sv2v_reg <= data_i[469];
      data_o_468_sv2v_reg <= data_i[468];
      data_o_467_sv2v_reg <= data_i[467];
      data_o_466_sv2v_reg <= data_i[466];
      data_o_465_sv2v_reg <= data_i[465];
      data_o_464_sv2v_reg <= data_i[464];
      data_o_463_sv2v_reg <= data_i[463];
      data_o_462_sv2v_reg <= data_i[462];
      data_o_461_sv2v_reg <= data_i[461];
      data_o_460_sv2v_reg <= data_i[460];
      data_o_459_sv2v_reg <= data_i[459];
      data_o_458_sv2v_reg <= data_i[458];
      data_o_457_sv2v_reg <= data_i[457];
      data_o_456_sv2v_reg <= data_i[456];
      data_o_455_sv2v_reg <= data_i[455];
      data_o_454_sv2v_reg <= data_i[454];
      data_o_453_sv2v_reg <= data_i[453];
      data_o_452_sv2v_reg <= data_i[452];
      data_o_451_sv2v_reg <= data_i[451];
      data_o_450_sv2v_reg <= data_i[450];
      data_o_449_sv2v_reg <= data_i[449];
      data_o_448_sv2v_reg <= data_i[448];
      data_o_447_sv2v_reg <= data_i[447];
      data_o_446_sv2v_reg <= data_i[446];
      data_o_445_sv2v_reg <= data_i[445];
      data_o_444_sv2v_reg <= data_i[444];
      data_o_443_sv2v_reg <= data_i[443];
      data_o_442_sv2v_reg <= data_i[442];
      data_o_441_sv2v_reg <= data_i[441];
      data_o_440_sv2v_reg <= data_i[440];
      data_o_439_sv2v_reg <= data_i[439];
      data_o_438_sv2v_reg <= data_i[438];
      data_o_437_sv2v_reg <= data_i[437];
      data_o_436_sv2v_reg <= data_i[436];
      data_o_435_sv2v_reg <= data_i[435];
      data_o_434_sv2v_reg <= data_i[434];
      data_o_433_sv2v_reg <= data_i[433];
      data_o_432_sv2v_reg <= data_i[432];
      data_o_431_sv2v_reg <= data_i[431];
      data_o_430_sv2v_reg <= data_i[430];
      data_o_429_sv2v_reg <= data_i[429];
      data_o_428_sv2v_reg <= data_i[428];
      data_o_427_sv2v_reg <= data_i[427];
      data_o_426_sv2v_reg <= data_i[426];
      data_o_425_sv2v_reg <= data_i[425];
      data_o_424_sv2v_reg <= data_i[424];
      data_o_423_sv2v_reg <= data_i[423];
      data_o_422_sv2v_reg <= data_i[422];
      data_o_421_sv2v_reg <= data_i[421];
      data_o_420_sv2v_reg <= data_i[420];
      data_o_419_sv2v_reg <= data_i[419];
      data_o_418_sv2v_reg <= data_i[418];
      data_o_417_sv2v_reg <= data_i[417];
      data_o_416_sv2v_reg <= data_i[416];
      data_o_415_sv2v_reg <= data_i[415];
      data_o_414_sv2v_reg <= data_i[414];
      data_o_413_sv2v_reg <= data_i[413];
      data_o_412_sv2v_reg <= data_i[412];
      data_o_411_sv2v_reg <= data_i[411];
      data_o_410_sv2v_reg <= data_i[410];
      data_o_409_sv2v_reg <= data_i[409];
      data_o_408_sv2v_reg <= data_i[408];
      data_o_407_sv2v_reg <= data_i[407];
      data_o_406_sv2v_reg <= data_i[406];
      data_o_405_sv2v_reg <= data_i[405];
      data_o_404_sv2v_reg <= data_i[404];
      data_o_403_sv2v_reg <= data_i[403];
      data_o_402_sv2v_reg <= data_i[402];
      data_o_401_sv2v_reg <= data_i[401];
      data_o_400_sv2v_reg <= data_i[400];
      data_o_399_sv2v_reg <= data_i[399];
      data_o_398_sv2v_reg <= data_i[398];
      data_o_397_sv2v_reg <= data_i[397];
      data_o_396_sv2v_reg <= data_i[396];
      data_o_395_sv2v_reg <= data_i[395];
      data_o_394_sv2v_reg <= data_i[394];
      data_o_393_sv2v_reg <= data_i[393];
      data_o_392_sv2v_reg <= data_i[392];
      data_o_391_sv2v_reg <= data_i[391];
      data_o_390_sv2v_reg <= data_i[390];
      data_o_389_sv2v_reg <= data_i[389];
      data_o_388_sv2v_reg <= data_i[388];
      data_o_387_sv2v_reg <= data_i[387];
      data_o_386_sv2v_reg <= data_i[386];
      data_o_385_sv2v_reg <= data_i[385];
      data_o_384_sv2v_reg <= data_i[384];
      data_o_383_sv2v_reg <= data_i[383];
      data_o_382_sv2v_reg <= data_i[382];
      data_o_381_sv2v_reg <= data_i[381];
      data_o_380_sv2v_reg <= data_i[380];
      data_o_379_sv2v_reg <= data_i[379];
      data_o_378_sv2v_reg <= data_i[378];
      data_o_377_sv2v_reg <= data_i[377];
      data_o_376_sv2v_reg <= data_i[376];
      data_o_375_sv2v_reg <= data_i[375];
      data_o_374_sv2v_reg <= data_i[374];
      data_o_373_sv2v_reg <= data_i[373];
      data_o_372_sv2v_reg <= data_i[372];
      data_o_371_sv2v_reg <= data_i[371];
      data_o_370_sv2v_reg <= data_i[370];
      data_o_369_sv2v_reg <= data_i[369];
      data_o_368_sv2v_reg <= data_i[368];
      data_o_367_sv2v_reg <= data_i[367];
      data_o_366_sv2v_reg <= data_i[366];
      data_o_365_sv2v_reg <= data_i[365];
      data_o_364_sv2v_reg <= data_i[364];
      data_o_363_sv2v_reg <= data_i[363];
      data_o_362_sv2v_reg <= data_i[362];
      data_o_361_sv2v_reg <= data_i[361];
      data_o_360_sv2v_reg <= data_i[360];
      data_o_359_sv2v_reg <= data_i[359];
      data_o_358_sv2v_reg <= data_i[358];
      data_o_357_sv2v_reg <= data_i[357];
      data_o_356_sv2v_reg <= data_i[356];
      data_o_355_sv2v_reg <= data_i[355];
      data_o_354_sv2v_reg <= data_i[354];
      data_o_353_sv2v_reg <= data_i[353];
      data_o_352_sv2v_reg <= data_i[352];
      data_o_351_sv2v_reg <= data_i[351];
      data_o_350_sv2v_reg <= data_i[350];
      data_o_349_sv2v_reg <= data_i[349];
      data_o_348_sv2v_reg <= data_i[348];
      data_o_347_sv2v_reg <= data_i[347];
      data_o_346_sv2v_reg <= data_i[346];
      data_o_345_sv2v_reg <= data_i[345];
      data_o_344_sv2v_reg <= data_i[344];
      data_o_343_sv2v_reg <= data_i[343];
      data_o_342_sv2v_reg <= data_i[342];
      data_o_341_sv2v_reg <= data_i[341];
      data_o_340_sv2v_reg <= data_i[340];
      data_o_339_sv2v_reg <= data_i[339];
      data_o_338_sv2v_reg <= data_i[338];
      data_o_337_sv2v_reg <= data_i[337];
      data_o_336_sv2v_reg <= data_i[336];
      data_o_335_sv2v_reg <= data_i[335];
      data_o_334_sv2v_reg <= data_i[334];
      data_o_333_sv2v_reg <= data_i[333];
      data_o_332_sv2v_reg <= data_i[332];
      data_o_331_sv2v_reg <= data_i[331];
      data_o_330_sv2v_reg <= data_i[330];
      data_o_329_sv2v_reg <= data_i[329];
      data_o_328_sv2v_reg <= data_i[328];
      data_o_327_sv2v_reg <= data_i[327];
      data_o_326_sv2v_reg <= data_i[326];
      data_o_325_sv2v_reg <= data_i[325];
      data_o_324_sv2v_reg <= data_i[324];
      data_o_323_sv2v_reg <= data_i[323];
      data_o_322_sv2v_reg <= data_i[322];
      data_o_321_sv2v_reg <= data_i[321];
      data_o_320_sv2v_reg <= data_i[320];
      data_o_319_sv2v_reg <= data_i[319];
      data_o_318_sv2v_reg <= data_i[318];
      data_o_317_sv2v_reg <= data_i[317];
      data_o_316_sv2v_reg <= data_i[316];
      data_o_315_sv2v_reg <= data_i[315];
      data_o_314_sv2v_reg <= data_i[314];
      data_o_313_sv2v_reg <= data_i[313];
      data_o_312_sv2v_reg <= data_i[312];
      data_o_311_sv2v_reg <= data_i[311];
      data_o_310_sv2v_reg <= data_i[310];
      data_o_309_sv2v_reg <= data_i[309];
      data_o_308_sv2v_reg <= data_i[308];
      data_o_307_sv2v_reg <= data_i[307];
      data_o_306_sv2v_reg <= data_i[306];
      data_o_305_sv2v_reg <= data_i[305];
      data_o_304_sv2v_reg <= data_i[304];
      data_o_303_sv2v_reg <= data_i[303];
      data_o_302_sv2v_reg <= data_i[302];
      data_o_301_sv2v_reg <= data_i[301];
      data_o_300_sv2v_reg <= data_i[300];
      data_o_299_sv2v_reg <= data_i[299];
      data_o_298_sv2v_reg <= data_i[298];
      data_o_297_sv2v_reg <= data_i[297];
      data_o_296_sv2v_reg <= data_i[296];
      data_o_295_sv2v_reg <= data_i[295];
      data_o_294_sv2v_reg <= data_i[294];
      data_o_293_sv2v_reg <= data_i[293];
      data_o_292_sv2v_reg <= data_i[292];
      data_o_291_sv2v_reg <= data_i[291];
      data_o_290_sv2v_reg <= data_i[290];
      data_o_289_sv2v_reg <= data_i[289];
      data_o_288_sv2v_reg <= data_i[288];
      data_o_287_sv2v_reg <= data_i[287];
      data_o_286_sv2v_reg <= data_i[286];
      data_o_285_sv2v_reg <= data_i[285];
      data_o_284_sv2v_reg <= data_i[284];
      data_o_283_sv2v_reg <= data_i[283];
      data_o_282_sv2v_reg <= data_i[282];
      data_o_281_sv2v_reg <= data_i[281];
      data_o_280_sv2v_reg <= data_i[280];
      data_o_279_sv2v_reg <= data_i[279];
      data_o_278_sv2v_reg <= data_i[278];
      data_o_277_sv2v_reg <= data_i[277];
      data_o_276_sv2v_reg <= data_i[276];
      data_o_275_sv2v_reg <= data_i[275];
      data_o_274_sv2v_reg <= data_i[274];
      data_o_273_sv2v_reg <= data_i[273];
      data_o_272_sv2v_reg <= data_i[272];
      data_o_271_sv2v_reg <= data_i[271];
      data_o_270_sv2v_reg <= data_i[270];
      data_o_269_sv2v_reg <= data_i[269];
      data_o_268_sv2v_reg <= data_i[268];
      data_o_267_sv2v_reg <= data_i[267];
      data_o_266_sv2v_reg <= data_i[266];
      data_o_265_sv2v_reg <= data_i[265];
      data_o_264_sv2v_reg <= data_i[264];
      data_o_263_sv2v_reg <= data_i[263];
      data_o_262_sv2v_reg <= data_i[262];
      data_o_261_sv2v_reg <= data_i[261];
      data_o_260_sv2v_reg <= data_i[260];
      data_o_259_sv2v_reg <= data_i[259];
      data_o_258_sv2v_reg <= data_i[258];
      data_o_257_sv2v_reg <= data_i[257];
      data_o_256_sv2v_reg <= data_i[256];
      data_o_255_sv2v_reg <= data_i[255];
      data_o_254_sv2v_reg <= data_i[254];
      data_o_253_sv2v_reg <= data_i[253];
      data_o_252_sv2v_reg <= data_i[252];
      data_o_251_sv2v_reg <= data_i[251];
      data_o_250_sv2v_reg <= data_i[250];
      data_o_249_sv2v_reg <= data_i[249];
      data_o_248_sv2v_reg <= data_i[248];
      data_o_247_sv2v_reg <= data_i[247];
      data_o_246_sv2v_reg <= data_i[246];
      data_o_245_sv2v_reg <= data_i[245];
      data_o_244_sv2v_reg <= data_i[244];
      data_o_243_sv2v_reg <= data_i[243];
      data_o_242_sv2v_reg <= data_i[242];
      data_o_241_sv2v_reg <= data_i[241];
      data_o_240_sv2v_reg <= data_i[240];
      data_o_239_sv2v_reg <= data_i[239];
      data_o_238_sv2v_reg <= data_i[238];
      data_o_237_sv2v_reg <= data_i[237];
      data_o_236_sv2v_reg <= data_i[236];
      data_o_235_sv2v_reg <= data_i[235];
      data_o_234_sv2v_reg <= data_i[234];
      data_o_233_sv2v_reg <= data_i[233];
      data_o_232_sv2v_reg <= data_i[232];
      data_o_231_sv2v_reg <= data_i[231];
      data_o_230_sv2v_reg <= data_i[230];
      data_o_229_sv2v_reg <= data_i[229];
      data_o_228_sv2v_reg <= data_i[228];
      data_o_227_sv2v_reg <= data_i[227];
      data_o_226_sv2v_reg <= data_i[226];
      data_o_225_sv2v_reg <= data_i[225];
      data_o_224_sv2v_reg <= data_i[224];
      data_o_223_sv2v_reg <= data_i[223];
      data_o_222_sv2v_reg <= data_i[222];
      data_o_221_sv2v_reg <= data_i[221];
      data_o_220_sv2v_reg <= data_i[220];
      data_o_219_sv2v_reg <= data_i[219];
      data_o_218_sv2v_reg <= data_i[218];
      data_o_217_sv2v_reg <= data_i[217];
      data_o_216_sv2v_reg <= data_i[216];
      data_o_215_sv2v_reg <= data_i[215];
      data_o_214_sv2v_reg <= data_i[214];
      data_o_213_sv2v_reg <= data_i[213];
      data_o_212_sv2v_reg <= data_i[212];
      data_o_211_sv2v_reg <= data_i[211];
      data_o_210_sv2v_reg <= data_i[210];
      data_o_209_sv2v_reg <= data_i[209];
      data_o_208_sv2v_reg <= data_i[208];
      data_o_207_sv2v_reg <= data_i[207];
      data_o_206_sv2v_reg <= data_i[206];
      data_o_205_sv2v_reg <= data_i[205];
      data_o_204_sv2v_reg <= data_i[204];
      data_o_203_sv2v_reg <= data_i[203];
      data_o_202_sv2v_reg <= data_i[202];
      data_o_201_sv2v_reg <= data_i[201];
      data_o_200_sv2v_reg <= data_i[200];
      data_o_199_sv2v_reg <= data_i[199];
      data_o_198_sv2v_reg <= data_i[198];
      data_o_197_sv2v_reg <= data_i[197];
      data_o_196_sv2v_reg <= data_i[196];
      data_o_195_sv2v_reg <= data_i[195];
      data_o_194_sv2v_reg <= data_i[194];
      data_o_193_sv2v_reg <= data_i[193];
      data_o_192_sv2v_reg <= data_i[192];
      data_o_191_sv2v_reg <= data_i[191];
      data_o_190_sv2v_reg <= data_i[190];
      data_o_189_sv2v_reg <= data_i[189];
      data_o_188_sv2v_reg <= data_i[188];
      data_o_187_sv2v_reg <= data_i[187];
      data_o_186_sv2v_reg <= data_i[186];
      data_o_185_sv2v_reg <= data_i[185];
      data_o_184_sv2v_reg <= data_i[184];
      data_o_183_sv2v_reg <= data_i[183];
      data_o_182_sv2v_reg <= data_i[182];
      data_o_181_sv2v_reg <= data_i[181];
      data_o_180_sv2v_reg <= data_i[180];
      data_o_179_sv2v_reg <= data_i[179];
      data_o_178_sv2v_reg <= data_i[178];
      data_o_177_sv2v_reg <= data_i[177];
      data_o_176_sv2v_reg <= data_i[176];
      data_o_175_sv2v_reg <= data_i[175];
      data_o_174_sv2v_reg <= data_i[174];
      data_o_173_sv2v_reg <= data_i[173];
      data_o_172_sv2v_reg <= data_i[172];
      data_o_171_sv2v_reg <= data_i[171];
      data_o_170_sv2v_reg <= data_i[170];
      data_o_169_sv2v_reg <= data_i[169];
      data_o_168_sv2v_reg <= data_i[168];
      data_o_167_sv2v_reg <= data_i[167];
      data_o_166_sv2v_reg <= data_i[166];
      data_o_165_sv2v_reg <= data_i[165];
      data_o_164_sv2v_reg <= data_i[164];
      data_o_163_sv2v_reg <= data_i[163];
      data_o_162_sv2v_reg <= data_i[162];
      data_o_161_sv2v_reg <= data_i[161];
      data_o_160_sv2v_reg <= data_i[160];
      data_o_159_sv2v_reg <= data_i[159];
      data_o_158_sv2v_reg <= data_i[158];
      data_o_157_sv2v_reg <= data_i[157];
      data_o_156_sv2v_reg <= data_i[156];
      data_o_155_sv2v_reg <= data_i[155];
      data_o_154_sv2v_reg <= data_i[154];
      data_o_153_sv2v_reg <= data_i[153];
      data_o_152_sv2v_reg <= data_i[152];
      data_o_151_sv2v_reg <= data_i[151];
      data_o_150_sv2v_reg <= data_i[150];
      data_o_149_sv2v_reg <= data_i[149];
      data_o_148_sv2v_reg <= data_i[148];
      data_o_147_sv2v_reg <= data_i[147];
      data_o_146_sv2v_reg <= data_i[146];
      data_o_145_sv2v_reg <= data_i[145];
      data_o_144_sv2v_reg <= data_i[144];
      data_o_143_sv2v_reg <= data_i[143];
      data_o_142_sv2v_reg <= data_i[142];
      data_o_141_sv2v_reg <= data_i[141];
      data_o_140_sv2v_reg <= data_i[140];
      data_o_139_sv2v_reg <= data_i[139];
      data_o_138_sv2v_reg <= data_i[138];
      data_o_137_sv2v_reg <= data_i[137];
      data_o_136_sv2v_reg <= data_i[136];
      data_o_135_sv2v_reg <= data_i[135];
      data_o_134_sv2v_reg <= data_i[134];
      data_o_133_sv2v_reg <= data_i[133];
      data_o_132_sv2v_reg <= data_i[132];
      data_o_131_sv2v_reg <= data_i[131];
      data_o_130_sv2v_reg <= data_i[130];
      data_o_129_sv2v_reg <= data_i[129];
      data_o_128_sv2v_reg <= data_i[128];
      data_o_127_sv2v_reg <= data_i[127];
      data_o_126_sv2v_reg <= data_i[126];
      data_o_125_sv2v_reg <= data_i[125];
      data_o_124_sv2v_reg <= data_i[124];
      data_o_123_sv2v_reg <= data_i[123];
      data_o_122_sv2v_reg <= data_i[122];
      data_o_121_sv2v_reg <= data_i[121];
      data_o_120_sv2v_reg <= data_i[120];
      data_o_119_sv2v_reg <= data_i[119];
      data_o_118_sv2v_reg <= data_i[118];
      data_o_117_sv2v_reg <= data_i[117];
      data_o_116_sv2v_reg <= data_i[116];
      data_o_115_sv2v_reg <= data_i[115];
      data_o_114_sv2v_reg <= data_i[114];
      data_o_113_sv2v_reg <= data_i[113];
      data_o_112_sv2v_reg <= data_i[112];
      data_o_111_sv2v_reg <= data_i[111];
      data_o_110_sv2v_reg <= data_i[110];
      data_o_109_sv2v_reg <= data_i[109];
      data_o_108_sv2v_reg <= data_i[108];
      data_o_107_sv2v_reg <= data_i[107];
      data_o_106_sv2v_reg <= data_i[106];
      data_o_105_sv2v_reg <= data_i[105];
      data_o_104_sv2v_reg <= data_i[104];
      data_o_103_sv2v_reg <= data_i[103];
      data_o_102_sv2v_reg <= data_i[102];
      data_o_101_sv2v_reg <= data_i[101];
      data_o_100_sv2v_reg <= data_i[100];
      data_o_99_sv2v_reg <= data_i[99];
      data_o_98_sv2v_reg <= data_i[98];
      data_o_97_sv2v_reg <= data_i[97];
      data_o_96_sv2v_reg <= data_i[96];
      data_o_95_sv2v_reg <= data_i[95];
      data_o_94_sv2v_reg <= data_i[94];
      data_o_93_sv2v_reg <= data_i[93];
      data_o_92_sv2v_reg <= data_i[92];
      data_o_91_sv2v_reg <= data_i[91];
      data_o_90_sv2v_reg <= data_i[90];
      data_o_89_sv2v_reg <= data_i[89];
      data_o_88_sv2v_reg <= data_i[88];
      data_o_87_sv2v_reg <= data_i[87];
      data_o_86_sv2v_reg <= data_i[86];
      data_o_85_sv2v_reg <= data_i[85];
      data_o_84_sv2v_reg <= data_i[84];
      data_o_83_sv2v_reg <= data_i[83];
      data_o_82_sv2v_reg <= data_i[82];
      data_o_81_sv2v_reg <= data_i[81];
      data_o_80_sv2v_reg <= data_i[80];
      data_o_79_sv2v_reg <= data_i[79];
      data_o_78_sv2v_reg <= data_i[78];
      data_o_77_sv2v_reg <= data_i[77];
      data_o_76_sv2v_reg <= data_i[76];
      data_o_75_sv2v_reg <= data_i[75];
      data_o_74_sv2v_reg <= data_i[74];
      data_o_73_sv2v_reg <= data_i[73];
      data_o_72_sv2v_reg <= data_i[72];
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_encode_one_hot_00000008_1
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o,v_2__0_,v_1__6_,v_1__4_,v_1__2_,v_1__0_,addr_2__4_,addr_2__0_;
  assign v_1__0_ = i[1] | i[0];
  assign v_1__2_ = i[3] | i[2];
  assign v_1__4_ = i[5] | i[4];
  assign v_1__6_ = i[7] | i[6];
  assign v_2__0_ = v_1__2_ | v_1__0_;
  assign addr_2__0_ = i[1] | i[3];
  assign addr_o[2] = v_1__6_ | v_1__4_;
  assign addr_2__4_ = i[5] | i[7];
  assign v_o = addr_o[2] | v_2__0_;
  assign addr_o[1] = v_1__2_ | v_1__6_;
  assign addr_o[0] = addr_2__0_ | addr_2__4_;

endmodule



module bsg_adder_one_hot_00000008
(
  a_i,
  b_i,
  o
);

  input [7:0] a_i;
  input [7:0] b_i;
  output [7:0] o;
  wire [7:0] o,\rof_0_.aggregate ,\rof_1_.aggregate ,\rof_2_.aggregate ,\rof_3_.aggregate ,
  \rof_4_.aggregate ,\rof_5_.aggregate ,\rof_6_.aggregate ,\rof_7_.aggregate ;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47;
  assign \rof_0_.aggregate [0] = a_i[0] & b_i[0];
  assign \rof_0_.aggregate [1] = a_i[1] & b_i[7];
  assign \rof_0_.aggregate [2] = a_i[2] & b_i[6];
  assign \rof_0_.aggregate [3] = a_i[3] & b_i[5];
  assign \rof_0_.aggregate [4] = a_i[4] & b_i[4];
  assign \rof_0_.aggregate [5] = a_i[5] & b_i[3];
  assign \rof_0_.aggregate [6] = a_i[6] & b_i[2];
  assign \rof_0_.aggregate [7] = a_i[7] & b_i[1];
  assign o[0] = N5 | \rof_0_.aggregate [0];
  assign N5 = N4 | \rof_0_.aggregate [1];
  assign N4 = N3 | \rof_0_.aggregate [2];
  assign N3 = N2 | \rof_0_.aggregate [3];
  assign N2 = N1 | \rof_0_.aggregate [4];
  assign N1 = N0 | \rof_0_.aggregate [5];
  assign N0 = \rof_0_.aggregate [7] | \rof_0_.aggregate [6];
  assign \rof_1_.aggregate [0] = a_i[0] & b_i[1];
  assign \rof_1_.aggregate [1] = a_i[1] & b_i[0];
  assign \rof_1_.aggregate [2] = a_i[2] & b_i[7];
  assign \rof_1_.aggregate [3] = a_i[3] & b_i[6];
  assign \rof_1_.aggregate [4] = a_i[4] & b_i[5];
  assign \rof_1_.aggregate [5] = a_i[5] & b_i[4];
  assign \rof_1_.aggregate [6] = a_i[6] & b_i[3];
  assign \rof_1_.aggregate [7] = a_i[7] & b_i[2];
  assign o[1] = N11 | \rof_1_.aggregate [0];
  assign N11 = N10 | \rof_1_.aggregate [1];
  assign N10 = N9 | \rof_1_.aggregate [2];
  assign N9 = N8 | \rof_1_.aggregate [3];
  assign N8 = N7 | \rof_1_.aggregate [4];
  assign N7 = N6 | \rof_1_.aggregate [5];
  assign N6 = \rof_1_.aggregate [7] | \rof_1_.aggregate [6];
  assign \rof_2_.aggregate [0] = a_i[0] & b_i[2];
  assign \rof_2_.aggregate [1] = a_i[1] & b_i[1];
  assign \rof_2_.aggregate [2] = a_i[2] & b_i[0];
  assign \rof_2_.aggregate [3] = a_i[3] & b_i[7];
  assign \rof_2_.aggregate [4] = a_i[4] & b_i[6];
  assign \rof_2_.aggregate [5] = a_i[5] & b_i[5];
  assign \rof_2_.aggregate [6] = a_i[6] & b_i[4];
  assign \rof_2_.aggregate [7] = a_i[7] & b_i[3];
  assign o[2] = N17 | \rof_2_.aggregate [0];
  assign N17 = N16 | \rof_2_.aggregate [1];
  assign N16 = N15 | \rof_2_.aggregate [2];
  assign N15 = N14 | \rof_2_.aggregate [3];
  assign N14 = N13 | \rof_2_.aggregate [4];
  assign N13 = N12 | \rof_2_.aggregate [5];
  assign N12 = \rof_2_.aggregate [7] | \rof_2_.aggregate [6];
  assign \rof_3_.aggregate [0] = a_i[0] & b_i[3];
  assign \rof_3_.aggregate [1] = a_i[1] & b_i[2];
  assign \rof_3_.aggregate [2] = a_i[2] & b_i[1];
  assign \rof_3_.aggregate [3] = a_i[3] & b_i[0];
  assign \rof_3_.aggregate [4] = a_i[4] & b_i[7];
  assign \rof_3_.aggregate [5] = a_i[5] & b_i[6];
  assign \rof_3_.aggregate [6] = a_i[6] & b_i[5];
  assign \rof_3_.aggregate [7] = a_i[7] & b_i[4];
  assign o[3] = N23 | \rof_3_.aggregate [0];
  assign N23 = N22 | \rof_3_.aggregate [1];
  assign N22 = N21 | \rof_3_.aggregate [2];
  assign N21 = N20 | \rof_3_.aggregate [3];
  assign N20 = N19 | \rof_3_.aggregate [4];
  assign N19 = N18 | \rof_3_.aggregate [5];
  assign N18 = \rof_3_.aggregate [7] | \rof_3_.aggregate [6];
  assign \rof_4_.aggregate [0] = a_i[0] & b_i[4];
  assign \rof_4_.aggregate [1] = a_i[1] & b_i[3];
  assign \rof_4_.aggregate [2] = a_i[2] & b_i[2];
  assign \rof_4_.aggregate [3] = a_i[3] & b_i[1];
  assign \rof_4_.aggregate [4] = a_i[4] & b_i[0];
  assign \rof_4_.aggregate [5] = a_i[5] & b_i[7];
  assign \rof_4_.aggregate [6] = a_i[6] & b_i[6];
  assign \rof_4_.aggregate [7] = a_i[7] & b_i[5];
  assign o[4] = N29 | \rof_4_.aggregate [0];
  assign N29 = N28 | \rof_4_.aggregate [1];
  assign N28 = N27 | \rof_4_.aggregate [2];
  assign N27 = N26 | \rof_4_.aggregate [3];
  assign N26 = N25 | \rof_4_.aggregate [4];
  assign N25 = N24 | \rof_4_.aggregate [5];
  assign N24 = \rof_4_.aggregate [7] | \rof_4_.aggregate [6];
  assign \rof_5_.aggregate [0] = a_i[0] & b_i[5];
  assign \rof_5_.aggregate [1] = a_i[1] & b_i[4];
  assign \rof_5_.aggregate [2] = a_i[2] & b_i[3];
  assign \rof_5_.aggregate [3] = a_i[3] & b_i[2];
  assign \rof_5_.aggregate [4] = a_i[4] & b_i[1];
  assign \rof_5_.aggregate [5] = a_i[5] & b_i[0];
  assign \rof_5_.aggregate [6] = a_i[6] & b_i[7];
  assign \rof_5_.aggregate [7] = a_i[7] & b_i[6];
  assign o[5] = N35 | \rof_5_.aggregate [0];
  assign N35 = N34 | \rof_5_.aggregate [1];
  assign N34 = N33 | \rof_5_.aggregate [2];
  assign N33 = N32 | \rof_5_.aggregate [3];
  assign N32 = N31 | \rof_5_.aggregate [4];
  assign N31 = N30 | \rof_5_.aggregate [5];
  assign N30 = \rof_5_.aggregate [7] | \rof_5_.aggregate [6];
  assign \rof_6_.aggregate [0] = a_i[0] & b_i[6];
  assign \rof_6_.aggregate [1] = a_i[1] & b_i[5];
  assign \rof_6_.aggregate [2] = a_i[2] & b_i[4];
  assign \rof_6_.aggregate [3] = a_i[3] & b_i[3];
  assign \rof_6_.aggregate [4] = a_i[4] & b_i[2];
  assign \rof_6_.aggregate [5] = a_i[5] & b_i[1];
  assign \rof_6_.aggregate [6] = a_i[6] & b_i[0];
  assign \rof_6_.aggregate [7] = a_i[7] & b_i[7];
  assign o[6] = N41 | \rof_6_.aggregate [0];
  assign N41 = N40 | \rof_6_.aggregate [1];
  assign N40 = N39 | \rof_6_.aggregate [2];
  assign N39 = N38 | \rof_6_.aggregate [3];
  assign N38 = N37 | \rof_6_.aggregate [4];
  assign N37 = N36 | \rof_6_.aggregate [5];
  assign N36 = \rof_6_.aggregate [7] | \rof_6_.aggregate [6];
  assign \rof_7_.aggregate [0] = a_i[0] & b_i[7];
  assign \rof_7_.aggregate [1] = a_i[1] & b_i[6];
  assign \rof_7_.aggregate [2] = a_i[2] & b_i[5];
  assign \rof_7_.aggregate [3] = a_i[3] & b_i[4];
  assign \rof_7_.aggregate [4] = a_i[4] & b_i[3];
  assign \rof_7_.aggregate [5] = a_i[5] & b_i[2];
  assign \rof_7_.aggregate [6] = a_i[6] & b_i[1];
  assign \rof_7_.aggregate [7] = a_i[7] & b_i[0];
  assign o[7] = N47 | \rof_7_.aggregate [0];
  assign N47 = N46 | \rof_7_.aggregate [1];
  assign N46 = N45 | \rof_7_.aggregate [2];
  assign N45 = N44 | \rof_7_.aggregate [3];
  assign N44 = N43 | \rof_7_.aggregate [4];
  assign N43 = N42 | \rof_7_.aggregate [5];
  assign N42 = \rof_7_.aggregate [7] | \rof_7_.aggregate [6];

endmodule



module bsg_mux_one_hot_00000040_00000008
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [511:0] data_i;
  input [7:0] sel_one_hot_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383;
  wire [511:0] data_masked;
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[1];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[1];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[1];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[2];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[2];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[2];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[2];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[2];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[2];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[2];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[2];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[2];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[2];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[2];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[2];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[2];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[2];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[2];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[2];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[2];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[2];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[2];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[2];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[2];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[2];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[2];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[2];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[2];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[2];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[2];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[2];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[2];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[2];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[2];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[2];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[2];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[2];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[2];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[2];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[2];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[2];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[2];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[2];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[2];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[2];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[2];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[2];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[2];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[2];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[2];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[2];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[2];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[2];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[2];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[2];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[2];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[2];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[2];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[2];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[2];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[2];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[2];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[2];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[2];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[2];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[2];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[2];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[3];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[3];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[3];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[3];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[3];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[3];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[3];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[3];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[3];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[3];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[3];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[3];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[3];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[3];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[3];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[3];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[3];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[3];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[3];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[3];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[3];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[3];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[3];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[3];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[3];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[3];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[3];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[3];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[3];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[3];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[3];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[3];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[3];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[3];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[3];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[3];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[3];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[3];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[3];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[3];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[3];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[3];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[3];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[3];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[3];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[3];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[3];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[3];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[3];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[3];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[3];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[3];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[3];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[3];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[3];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[3];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[3];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[3];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[3];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[3];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[3];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[3];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[3];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[3];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[4];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[4];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[4];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[4];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[4];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[4];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[4];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[4];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[4];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[4];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[4];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[4];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[4];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[4];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[4];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[4];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[4];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[4];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[4];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[4];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[4];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[4];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[4];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[4];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[4];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[4];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[4];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[4];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[4];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[4];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[4];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[4];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[4];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[4];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[4];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[4];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[4];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[4];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[4];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[4];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[4];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[4];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[4];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[4];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[4];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[4];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[4];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[4];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[4];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[4];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[4];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[4];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[4];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[4];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[4];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[4];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[4];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[4];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[4];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[4];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[4];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[4];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[4];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[4];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[5];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[5];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[5];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[5];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[5];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[5];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[5];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[5];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[5];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[5];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[5];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[5];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[5];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[5];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[5];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[5];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[5];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[5];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[5];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[5];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[5];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[5];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[5];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[5];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[5];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[5];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[5];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[5];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[5];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[5];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[5];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[5];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[5];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[5];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[5];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[5];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[5];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[5];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[5];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[5];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[5];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[5];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[5];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[5];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[5];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[5];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[5];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[5];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[5];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[5];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[5];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[5];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[5];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[5];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[5];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[5];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[5];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[5];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[5];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[5];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[5];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[5];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[5];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[5];
  assign data_masked[447] = data_i[447] & sel_one_hot_i[6];
  assign data_masked[446] = data_i[446] & sel_one_hot_i[6];
  assign data_masked[445] = data_i[445] & sel_one_hot_i[6];
  assign data_masked[444] = data_i[444] & sel_one_hot_i[6];
  assign data_masked[443] = data_i[443] & sel_one_hot_i[6];
  assign data_masked[442] = data_i[442] & sel_one_hot_i[6];
  assign data_masked[441] = data_i[441] & sel_one_hot_i[6];
  assign data_masked[440] = data_i[440] & sel_one_hot_i[6];
  assign data_masked[439] = data_i[439] & sel_one_hot_i[6];
  assign data_masked[438] = data_i[438] & sel_one_hot_i[6];
  assign data_masked[437] = data_i[437] & sel_one_hot_i[6];
  assign data_masked[436] = data_i[436] & sel_one_hot_i[6];
  assign data_masked[435] = data_i[435] & sel_one_hot_i[6];
  assign data_masked[434] = data_i[434] & sel_one_hot_i[6];
  assign data_masked[433] = data_i[433] & sel_one_hot_i[6];
  assign data_masked[432] = data_i[432] & sel_one_hot_i[6];
  assign data_masked[431] = data_i[431] & sel_one_hot_i[6];
  assign data_masked[430] = data_i[430] & sel_one_hot_i[6];
  assign data_masked[429] = data_i[429] & sel_one_hot_i[6];
  assign data_masked[428] = data_i[428] & sel_one_hot_i[6];
  assign data_masked[427] = data_i[427] & sel_one_hot_i[6];
  assign data_masked[426] = data_i[426] & sel_one_hot_i[6];
  assign data_masked[425] = data_i[425] & sel_one_hot_i[6];
  assign data_masked[424] = data_i[424] & sel_one_hot_i[6];
  assign data_masked[423] = data_i[423] & sel_one_hot_i[6];
  assign data_masked[422] = data_i[422] & sel_one_hot_i[6];
  assign data_masked[421] = data_i[421] & sel_one_hot_i[6];
  assign data_masked[420] = data_i[420] & sel_one_hot_i[6];
  assign data_masked[419] = data_i[419] & sel_one_hot_i[6];
  assign data_masked[418] = data_i[418] & sel_one_hot_i[6];
  assign data_masked[417] = data_i[417] & sel_one_hot_i[6];
  assign data_masked[416] = data_i[416] & sel_one_hot_i[6];
  assign data_masked[415] = data_i[415] & sel_one_hot_i[6];
  assign data_masked[414] = data_i[414] & sel_one_hot_i[6];
  assign data_masked[413] = data_i[413] & sel_one_hot_i[6];
  assign data_masked[412] = data_i[412] & sel_one_hot_i[6];
  assign data_masked[411] = data_i[411] & sel_one_hot_i[6];
  assign data_masked[410] = data_i[410] & sel_one_hot_i[6];
  assign data_masked[409] = data_i[409] & sel_one_hot_i[6];
  assign data_masked[408] = data_i[408] & sel_one_hot_i[6];
  assign data_masked[407] = data_i[407] & sel_one_hot_i[6];
  assign data_masked[406] = data_i[406] & sel_one_hot_i[6];
  assign data_masked[405] = data_i[405] & sel_one_hot_i[6];
  assign data_masked[404] = data_i[404] & sel_one_hot_i[6];
  assign data_masked[403] = data_i[403] & sel_one_hot_i[6];
  assign data_masked[402] = data_i[402] & sel_one_hot_i[6];
  assign data_masked[401] = data_i[401] & sel_one_hot_i[6];
  assign data_masked[400] = data_i[400] & sel_one_hot_i[6];
  assign data_masked[399] = data_i[399] & sel_one_hot_i[6];
  assign data_masked[398] = data_i[398] & sel_one_hot_i[6];
  assign data_masked[397] = data_i[397] & sel_one_hot_i[6];
  assign data_masked[396] = data_i[396] & sel_one_hot_i[6];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[6];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[6];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[6];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[6];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[6];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[6];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[6];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[6];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[6];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[6];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[6];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[6];
  assign data_masked[511] = data_i[511] & sel_one_hot_i[7];
  assign data_masked[510] = data_i[510] & sel_one_hot_i[7];
  assign data_masked[509] = data_i[509] & sel_one_hot_i[7];
  assign data_masked[508] = data_i[508] & sel_one_hot_i[7];
  assign data_masked[507] = data_i[507] & sel_one_hot_i[7];
  assign data_masked[506] = data_i[506] & sel_one_hot_i[7];
  assign data_masked[505] = data_i[505] & sel_one_hot_i[7];
  assign data_masked[504] = data_i[504] & sel_one_hot_i[7];
  assign data_masked[503] = data_i[503] & sel_one_hot_i[7];
  assign data_masked[502] = data_i[502] & sel_one_hot_i[7];
  assign data_masked[501] = data_i[501] & sel_one_hot_i[7];
  assign data_masked[500] = data_i[500] & sel_one_hot_i[7];
  assign data_masked[499] = data_i[499] & sel_one_hot_i[7];
  assign data_masked[498] = data_i[498] & sel_one_hot_i[7];
  assign data_masked[497] = data_i[497] & sel_one_hot_i[7];
  assign data_masked[496] = data_i[496] & sel_one_hot_i[7];
  assign data_masked[495] = data_i[495] & sel_one_hot_i[7];
  assign data_masked[494] = data_i[494] & sel_one_hot_i[7];
  assign data_masked[493] = data_i[493] & sel_one_hot_i[7];
  assign data_masked[492] = data_i[492] & sel_one_hot_i[7];
  assign data_masked[491] = data_i[491] & sel_one_hot_i[7];
  assign data_masked[490] = data_i[490] & sel_one_hot_i[7];
  assign data_masked[489] = data_i[489] & sel_one_hot_i[7];
  assign data_masked[488] = data_i[488] & sel_one_hot_i[7];
  assign data_masked[487] = data_i[487] & sel_one_hot_i[7];
  assign data_masked[486] = data_i[486] & sel_one_hot_i[7];
  assign data_masked[485] = data_i[485] & sel_one_hot_i[7];
  assign data_masked[484] = data_i[484] & sel_one_hot_i[7];
  assign data_masked[483] = data_i[483] & sel_one_hot_i[7];
  assign data_masked[482] = data_i[482] & sel_one_hot_i[7];
  assign data_masked[481] = data_i[481] & sel_one_hot_i[7];
  assign data_masked[480] = data_i[480] & sel_one_hot_i[7];
  assign data_masked[479] = data_i[479] & sel_one_hot_i[7];
  assign data_masked[478] = data_i[478] & sel_one_hot_i[7];
  assign data_masked[477] = data_i[477] & sel_one_hot_i[7];
  assign data_masked[476] = data_i[476] & sel_one_hot_i[7];
  assign data_masked[475] = data_i[475] & sel_one_hot_i[7];
  assign data_masked[474] = data_i[474] & sel_one_hot_i[7];
  assign data_masked[473] = data_i[473] & sel_one_hot_i[7];
  assign data_masked[472] = data_i[472] & sel_one_hot_i[7];
  assign data_masked[471] = data_i[471] & sel_one_hot_i[7];
  assign data_masked[470] = data_i[470] & sel_one_hot_i[7];
  assign data_masked[469] = data_i[469] & sel_one_hot_i[7];
  assign data_masked[468] = data_i[468] & sel_one_hot_i[7];
  assign data_masked[467] = data_i[467] & sel_one_hot_i[7];
  assign data_masked[466] = data_i[466] & sel_one_hot_i[7];
  assign data_masked[465] = data_i[465] & sel_one_hot_i[7];
  assign data_masked[464] = data_i[464] & sel_one_hot_i[7];
  assign data_masked[463] = data_i[463] & sel_one_hot_i[7];
  assign data_masked[462] = data_i[462] & sel_one_hot_i[7];
  assign data_masked[461] = data_i[461] & sel_one_hot_i[7];
  assign data_masked[460] = data_i[460] & sel_one_hot_i[7];
  assign data_masked[459] = data_i[459] & sel_one_hot_i[7];
  assign data_masked[458] = data_i[458] & sel_one_hot_i[7];
  assign data_masked[457] = data_i[457] & sel_one_hot_i[7];
  assign data_masked[456] = data_i[456] & sel_one_hot_i[7];
  assign data_masked[455] = data_i[455] & sel_one_hot_i[7];
  assign data_masked[454] = data_i[454] & sel_one_hot_i[7];
  assign data_masked[453] = data_i[453] & sel_one_hot_i[7];
  assign data_masked[452] = data_i[452] & sel_one_hot_i[7];
  assign data_masked[451] = data_i[451] & sel_one_hot_i[7];
  assign data_masked[450] = data_i[450] & sel_one_hot_i[7];
  assign data_masked[449] = data_i[449] & sel_one_hot_i[7];
  assign data_masked[448] = data_i[448] & sel_one_hot_i[7];
  assign data_o[0] = N5 | data_masked[0];
  assign N5 = N4 | data_masked[64];
  assign N4 = N3 | data_masked[128];
  assign N3 = N2 | data_masked[192];
  assign N2 = N1 | data_masked[256];
  assign N1 = N0 | data_masked[320];
  assign N0 = data_masked[448] | data_masked[384];
  assign data_o[1] = N11 | data_masked[1];
  assign N11 = N10 | data_masked[65];
  assign N10 = N9 | data_masked[129];
  assign N9 = N8 | data_masked[193];
  assign N8 = N7 | data_masked[257];
  assign N7 = N6 | data_masked[321];
  assign N6 = data_masked[449] | data_masked[385];
  assign data_o[2] = N17 | data_masked[2];
  assign N17 = N16 | data_masked[66];
  assign N16 = N15 | data_masked[130];
  assign N15 = N14 | data_masked[194];
  assign N14 = N13 | data_masked[258];
  assign N13 = N12 | data_masked[322];
  assign N12 = data_masked[450] | data_masked[386];
  assign data_o[3] = N23 | data_masked[3];
  assign N23 = N22 | data_masked[67];
  assign N22 = N21 | data_masked[131];
  assign N21 = N20 | data_masked[195];
  assign N20 = N19 | data_masked[259];
  assign N19 = N18 | data_masked[323];
  assign N18 = data_masked[451] | data_masked[387];
  assign data_o[4] = N29 | data_masked[4];
  assign N29 = N28 | data_masked[68];
  assign N28 = N27 | data_masked[132];
  assign N27 = N26 | data_masked[196];
  assign N26 = N25 | data_masked[260];
  assign N25 = N24 | data_masked[324];
  assign N24 = data_masked[452] | data_masked[388];
  assign data_o[5] = N35 | data_masked[5];
  assign N35 = N34 | data_masked[69];
  assign N34 = N33 | data_masked[133];
  assign N33 = N32 | data_masked[197];
  assign N32 = N31 | data_masked[261];
  assign N31 = N30 | data_masked[325];
  assign N30 = data_masked[453] | data_masked[389];
  assign data_o[6] = N41 | data_masked[6];
  assign N41 = N40 | data_masked[70];
  assign N40 = N39 | data_masked[134];
  assign N39 = N38 | data_masked[198];
  assign N38 = N37 | data_masked[262];
  assign N37 = N36 | data_masked[326];
  assign N36 = data_masked[454] | data_masked[390];
  assign data_o[7] = N47 | data_masked[7];
  assign N47 = N46 | data_masked[71];
  assign N46 = N45 | data_masked[135];
  assign N45 = N44 | data_masked[199];
  assign N44 = N43 | data_masked[263];
  assign N43 = N42 | data_masked[327];
  assign N42 = data_masked[455] | data_masked[391];
  assign data_o[8] = N53 | data_masked[8];
  assign N53 = N52 | data_masked[72];
  assign N52 = N51 | data_masked[136];
  assign N51 = N50 | data_masked[200];
  assign N50 = N49 | data_masked[264];
  assign N49 = N48 | data_masked[328];
  assign N48 = data_masked[456] | data_masked[392];
  assign data_o[9] = N59 | data_masked[9];
  assign N59 = N58 | data_masked[73];
  assign N58 = N57 | data_masked[137];
  assign N57 = N56 | data_masked[201];
  assign N56 = N55 | data_masked[265];
  assign N55 = N54 | data_masked[329];
  assign N54 = data_masked[457] | data_masked[393];
  assign data_o[10] = N65 | data_masked[10];
  assign N65 = N64 | data_masked[74];
  assign N64 = N63 | data_masked[138];
  assign N63 = N62 | data_masked[202];
  assign N62 = N61 | data_masked[266];
  assign N61 = N60 | data_masked[330];
  assign N60 = data_masked[458] | data_masked[394];
  assign data_o[11] = N71 | data_masked[11];
  assign N71 = N70 | data_masked[75];
  assign N70 = N69 | data_masked[139];
  assign N69 = N68 | data_masked[203];
  assign N68 = N67 | data_masked[267];
  assign N67 = N66 | data_masked[331];
  assign N66 = data_masked[459] | data_masked[395];
  assign data_o[12] = N77 | data_masked[12];
  assign N77 = N76 | data_masked[76];
  assign N76 = N75 | data_masked[140];
  assign N75 = N74 | data_masked[204];
  assign N74 = N73 | data_masked[268];
  assign N73 = N72 | data_masked[332];
  assign N72 = data_masked[460] | data_masked[396];
  assign data_o[13] = N83 | data_masked[13];
  assign N83 = N82 | data_masked[77];
  assign N82 = N81 | data_masked[141];
  assign N81 = N80 | data_masked[205];
  assign N80 = N79 | data_masked[269];
  assign N79 = N78 | data_masked[333];
  assign N78 = data_masked[461] | data_masked[397];
  assign data_o[14] = N89 | data_masked[14];
  assign N89 = N88 | data_masked[78];
  assign N88 = N87 | data_masked[142];
  assign N87 = N86 | data_masked[206];
  assign N86 = N85 | data_masked[270];
  assign N85 = N84 | data_masked[334];
  assign N84 = data_masked[462] | data_masked[398];
  assign data_o[15] = N95 | data_masked[15];
  assign N95 = N94 | data_masked[79];
  assign N94 = N93 | data_masked[143];
  assign N93 = N92 | data_masked[207];
  assign N92 = N91 | data_masked[271];
  assign N91 = N90 | data_masked[335];
  assign N90 = data_masked[463] | data_masked[399];
  assign data_o[16] = N101 | data_masked[16];
  assign N101 = N100 | data_masked[80];
  assign N100 = N99 | data_masked[144];
  assign N99 = N98 | data_masked[208];
  assign N98 = N97 | data_masked[272];
  assign N97 = N96 | data_masked[336];
  assign N96 = data_masked[464] | data_masked[400];
  assign data_o[17] = N107 | data_masked[17];
  assign N107 = N106 | data_masked[81];
  assign N106 = N105 | data_masked[145];
  assign N105 = N104 | data_masked[209];
  assign N104 = N103 | data_masked[273];
  assign N103 = N102 | data_masked[337];
  assign N102 = data_masked[465] | data_masked[401];
  assign data_o[18] = N113 | data_masked[18];
  assign N113 = N112 | data_masked[82];
  assign N112 = N111 | data_masked[146];
  assign N111 = N110 | data_masked[210];
  assign N110 = N109 | data_masked[274];
  assign N109 = N108 | data_masked[338];
  assign N108 = data_masked[466] | data_masked[402];
  assign data_o[19] = N119 | data_masked[19];
  assign N119 = N118 | data_masked[83];
  assign N118 = N117 | data_masked[147];
  assign N117 = N116 | data_masked[211];
  assign N116 = N115 | data_masked[275];
  assign N115 = N114 | data_masked[339];
  assign N114 = data_masked[467] | data_masked[403];
  assign data_o[20] = N125 | data_masked[20];
  assign N125 = N124 | data_masked[84];
  assign N124 = N123 | data_masked[148];
  assign N123 = N122 | data_masked[212];
  assign N122 = N121 | data_masked[276];
  assign N121 = N120 | data_masked[340];
  assign N120 = data_masked[468] | data_masked[404];
  assign data_o[21] = N131 | data_masked[21];
  assign N131 = N130 | data_masked[85];
  assign N130 = N129 | data_masked[149];
  assign N129 = N128 | data_masked[213];
  assign N128 = N127 | data_masked[277];
  assign N127 = N126 | data_masked[341];
  assign N126 = data_masked[469] | data_masked[405];
  assign data_o[22] = N137 | data_masked[22];
  assign N137 = N136 | data_masked[86];
  assign N136 = N135 | data_masked[150];
  assign N135 = N134 | data_masked[214];
  assign N134 = N133 | data_masked[278];
  assign N133 = N132 | data_masked[342];
  assign N132 = data_masked[470] | data_masked[406];
  assign data_o[23] = N143 | data_masked[23];
  assign N143 = N142 | data_masked[87];
  assign N142 = N141 | data_masked[151];
  assign N141 = N140 | data_masked[215];
  assign N140 = N139 | data_masked[279];
  assign N139 = N138 | data_masked[343];
  assign N138 = data_masked[471] | data_masked[407];
  assign data_o[24] = N149 | data_masked[24];
  assign N149 = N148 | data_masked[88];
  assign N148 = N147 | data_masked[152];
  assign N147 = N146 | data_masked[216];
  assign N146 = N145 | data_masked[280];
  assign N145 = N144 | data_masked[344];
  assign N144 = data_masked[472] | data_masked[408];
  assign data_o[25] = N155 | data_masked[25];
  assign N155 = N154 | data_masked[89];
  assign N154 = N153 | data_masked[153];
  assign N153 = N152 | data_masked[217];
  assign N152 = N151 | data_masked[281];
  assign N151 = N150 | data_masked[345];
  assign N150 = data_masked[473] | data_masked[409];
  assign data_o[26] = N161 | data_masked[26];
  assign N161 = N160 | data_masked[90];
  assign N160 = N159 | data_masked[154];
  assign N159 = N158 | data_masked[218];
  assign N158 = N157 | data_masked[282];
  assign N157 = N156 | data_masked[346];
  assign N156 = data_masked[474] | data_masked[410];
  assign data_o[27] = N167 | data_masked[27];
  assign N167 = N166 | data_masked[91];
  assign N166 = N165 | data_masked[155];
  assign N165 = N164 | data_masked[219];
  assign N164 = N163 | data_masked[283];
  assign N163 = N162 | data_masked[347];
  assign N162 = data_masked[475] | data_masked[411];
  assign data_o[28] = N173 | data_masked[28];
  assign N173 = N172 | data_masked[92];
  assign N172 = N171 | data_masked[156];
  assign N171 = N170 | data_masked[220];
  assign N170 = N169 | data_masked[284];
  assign N169 = N168 | data_masked[348];
  assign N168 = data_masked[476] | data_masked[412];
  assign data_o[29] = N179 | data_masked[29];
  assign N179 = N178 | data_masked[93];
  assign N178 = N177 | data_masked[157];
  assign N177 = N176 | data_masked[221];
  assign N176 = N175 | data_masked[285];
  assign N175 = N174 | data_masked[349];
  assign N174 = data_masked[477] | data_masked[413];
  assign data_o[30] = N185 | data_masked[30];
  assign N185 = N184 | data_masked[94];
  assign N184 = N183 | data_masked[158];
  assign N183 = N182 | data_masked[222];
  assign N182 = N181 | data_masked[286];
  assign N181 = N180 | data_masked[350];
  assign N180 = data_masked[478] | data_masked[414];
  assign data_o[31] = N191 | data_masked[31];
  assign N191 = N190 | data_masked[95];
  assign N190 = N189 | data_masked[159];
  assign N189 = N188 | data_masked[223];
  assign N188 = N187 | data_masked[287];
  assign N187 = N186 | data_masked[351];
  assign N186 = data_masked[479] | data_masked[415];
  assign data_o[32] = N197 | data_masked[32];
  assign N197 = N196 | data_masked[96];
  assign N196 = N195 | data_masked[160];
  assign N195 = N194 | data_masked[224];
  assign N194 = N193 | data_masked[288];
  assign N193 = N192 | data_masked[352];
  assign N192 = data_masked[480] | data_masked[416];
  assign data_o[33] = N203 | data_masked[33];
  assign N203 = N202 | data_masked[97];
  assign N202 = N201 | data_masked[161];
  assign N201 = N200 | data_masked[225];
  assign N200 = N199 | data_masked[289];
  assign N199 = N198 | data_masked[353];
  assign N198 = data_masked[481] | data_masked[417];
  assign data_o[34] = N209 | data_masked[34];
  assign N209 = N208 | data_masked[98];
  assign N208 = N207 | data_masked[162];
  assign N207 = N206 | data_masked[226];
  assign N206 = N205 | data_masked[290];
  assign N205 = N204 | data_masked[354];
  assign N204 = data_masked[482] | data_masked[418];
  assign data_o[35] = N215 | data_masked[35];
  assign N215 = N214 | data_masked[99];
  assign N214 = N213 | data_masked[163];
  assign N213 = N212 | data_masked[227];
  assign N212 = N211 | data_masked[291];
  assign N211 = N210 | data_masked[355];
  assign N210 = data_masked[483] | data_masked[419];
  assign data_o[36] = N221 | data_masked[36];
  assign N221 = N220 | data_masked[100];
  assign N220 = N219 | data_masked[164];
  assign N219 = N218 | data_masked[228];
  assign N218 = N217 | data_masked[292];
  assign N217 = N216 | data_masked[356];
  assign N216 = data_masked[484] | data_masked[420];
  assign data_o[37] = N227 | data_masked[37];
  assign N227 = N226 | data_masked[101];
  assign N226 = N225 | data_masked[165];
  assign N225 = N224 | data_masked[229];
  assign N224 = N223 | data_masked[293];
  assign N223 = N222 | data_masked[357];
  assign N222 = data_masked[485] | data_masked[421];
  assign data_o[38] = N233 | data_masked[38];
  assign N233 = N232 | data_masked[102];
  assign N232 = N231 | data_masked[166];
  assign N231 = N230 | data_masked[230];
  assign N230 = N229 | data_masked[294];
  assign N229 = N228 | data_masked[358];
  assign N228 = data_masked[486] | data_masked[422];
  assign data_o[39] = N239 | data_masked[39];
  assign N239 = N238 | data_masked[103];
  assign N238 = N237 | data_masked[167];
  assign N237 = N236 | data_masked[231];
  assign N236 = N235 | data_masked[295];
  assign N235 = N234 | data_masked[359];
  assign N234 = data_masked[487] | data_masked[423];
  assign data_o[40] = N245 | data_masked[40];
  assign N245 = N244 | data_masked[104];
  assign N244 = N243 | data_masked[168];
  assign N243 = N242 | data_masked[232];
  assign N242 = N241 | data_masked[296];
  assign N241 = N240 | data_masked[360];
  assign N240 = data_masked[488] | data_masked[424];
  assign data_o[41] = N251 | data_masked[41];
  assign N251 = N250 | data_masked[105];
  assign N250 = N249 | data_masked[169];
  assign N249 = N248 | data_masked[233];
  assign N248 = N247 | data_masked[297];
  assign N247 = N246 | data_masked[361];
  assign N246 = data_masked[489] | data_masked[425];
  assign data_o[42] = N257 | data_masked[42];
  assign N257 = N256 | data_masked[106];
  assign N256 = N255 | data_masked[170];
  assign N255 = N254 | data_masked[234];
  assign N254 = N253 | data_masked[298];
  assign N253 = N252 | data_masked[362];
  assign N252 = data_masked[490] | data_masked[426];
  assign data_o[43] = N263 | data_masked[43];
  assign N263 = N262 | data_masked[107];
  assign N262 = N261 | data_masked[171];
  assign N261 = N260 | data_masked[235];
  assign N260 = N259 | data_masked[299];
  assign N259 = N258 | data_masked[363];
  assign N258 = data_masked[491] | data_masked[427];
  assign data_o[44] = N269 | data_masked[44];
  assign N269 = N268 | data_masked[108];
  assign N268 = N267 | data_masked[172];
  assign N267 = N266 | data_masked[236];
  assign N266 = N265 | data_masked[300];
  assign N265 = N264 | data_masked[364];
  assign N264 = data_masked[492] | data_masked[428];
  assign data_o[45] = N275 | data_masked[45];
  assign N275 = N274 | data_masked[109];
  assign N274 = N273 | data_masked[173];
  assign N273 = N272 | data_masked[237];
  assign N272 = N271 | data_masked[301];
  assign N271 = N270 | data_masked[365];
  assign N270 = data_masked[493] | data_masked[429];
  assign data_o[46] = N281 | data_masked[46];
  assign N281 = N280 | data_masked[110];
  assign N280 = N279 | data_masked[174];
  assign N279 = N278 | data_masked[238];
  assign N278 = N277 | data_masked[302];
  assign N277 = N276 | data_masked[366];
  assign N276 = data_masked[494] | data_masked[430];
  assign data_o[47] = N287 | data_masked[47];
  assign N287 = N286 | data_masked[111];
  assign N286 = N285 | data_masked[175];
  assign N285 = N284 | data_masked[239];
  assign N284 = N283 | data_masked[303];
  assign N283 = N282 | data_masked[367];
  assign N282 = data_masked[495] | data_masked[431];
  assign data_o[48] = N293 | data_masked[48];
  assign N293 = N292 | data_masked[112];
  assign N292 = N291 | data_masked[176];
  assign N291 = N290 | data_masked[240];
  assign N290 = N289 | data_masked[304];
  assign N289 = N288 | data_masked[368];
  assign N288 = data_masked[496] | data_masked[432];
  assign data_o[49] = N299 | data_masked[49];
  assign N299 = N298 | data_masked[113];
  assign N298 = N297 | data_masked[177];
  assign N297 = N296 | data_masked[241];
  assign N296 = N295 | data_masked[305];
  assign N295 = N294 | data_masked[369];
  assign N294 = data_masked[497] | data_masked[433];
  assign data_o[50] = N305 | data_masked[50];
  assign N305 = N304 | data_masked[114];
  assign N304 = N303 | data_masked[178];
  assign N303 = N302 | data_masked[242];
  assign N302 = N301 | data_masked[306];
  assign N301 = N300 | data_masked[370];
  assign N300 = data_masked[498] | data_masked[434];
  assign data_o[51] = N311 | data_masked[51];
  assign N311 = N310 | data_masked[115];
  assign N310 = N309 | data_masked[179];
  assign N309 = N308 | data_masked[243];
  assign N308 = N307 | data_masked[307];
  assign N307 = N306 | data_masked[371];
  assign N306 = data_masked[499] | data_masked[435];
  assign data_o[52] = N317 | data_masked[52];
  assign N317 = N316 | data_masked[116];
  assign N316 = N315 | data_masked[180];
  assign N315 = N314 | data_masked[244];
  assign N314 = N313 | data_masked[308];
  assign N313 = N312 | data_masked[372];
  assign N312 = data_masked[500] | data_masked[436];
  assign data_o[53] = N323 | data_masked[53];
  assign N323 = N322 | data_masked[117];
  assign N322 = N321 | data_masked[181];
  assign N321 = N320 | data_masked[245];
  assign N320 = N319 | data_masked[309];
  assign N319 = N318 | data_masked[373];
  assign N318 = data_masked[501] | data_masked[437];
  assign data_o[54] = N329 | data_masked[54];
  assign N329 = N328 | data_masked[118];
  assign N328 = N327 | data_masked[182];
  assign N327 = N326 | data_masked[246];
  assign N326 = N325 | data_masked[310];
  assign N325 = N324 | data_masked[374];
  assign N324 = data_masked[502] | data_masked[438];
  assign data_o[55] = N335 | data_masked[55];
  assign N335 = N334 | data_masked[119];
  assign N334 = N333 | data_masked[183];
  assign N333 = N332 | data_masked[247];
  assign N332 = N331 | data_masked[311];
  assign N331 = N330 | data_masked[375];
  assign N330 = data_masked[503] | data_masked[439];
  assign data_o[56] = N341 | data_masked[56];
  assign N341 = N340 | data_masked[120];
  assign N340 = N339 | data_masked[184];
  assign N339 = N338 | data_masked[248];
  assign N338 = N337 | data_masked[312];
  assign N337 = N336 | data_masked[376];
  assign N336 = data_masked[504] | data_masked[440];
  assign data_o[57] = N347 | data_masked[57];
  assign N347 = N346 | data_masked[121];
  assign N346 = N345 | data_masked[185];
  assign N345 = N344 | data_masked[249];
  assign N344 = N343 | data_masked[313];
  assign N343 = N342 | data_masked[377];
  assign N342 = data_masked[505] | data_masked[441];
  assign data_o[58] = N353 | data_masked[58];
  assign N353 = N352 | data_masked[122];
  assign N352 = N351 | data_masked[186];
  assign N351 = N350 | data_masked[250];
  assign N350 = N349 | data_masked[314];
  assign N349 = N348 | data_masked[378];
  assign N348 = data_masked[506] | data_masked[442];
  assign data_o[59] = N359 | data_masked[59];
  assign N359 = N358 | data_masked[123];
  assign N358 = N357 | data_masked[187];
  assign N357 = N356 | data_masked[251];
  assign N356 = N355 | data_masked[315];
  assign N355 = N354 | data_masked[379];
  assign N354 = data_masked[507] | data_masked[443];
  assign data_o[60] = N365 | data_masked[60];
  assign N365 = N364 | data_masked[124];
  assign N364 = N363 | data_masked[188];
  assign N363 = N362 | data_masked[252];
  assign N362 = N361 | data_masked[316];
  assign N361 = N360 | data_masked[380];
  assign N360 = data_masked[508] | data_masked[444];
  assign data_o[61] = N371 | data_masked[61];
  assign N371 = N370 | data_masked[125];
  assign N370 = N369 | data_masked[189];
  assign N369 = N368 | data_masked[253];
  assign N368 = N367 | data_masked[317];
  assign N367 = N366 | data_masked[381];
  assign N366 = data_masked[509] | data_masked[445];
  assign data_o[62] = N377 | data_masked[62];
  assign N377 = N376 | data_masked[126];
  assign N376 = N375 | data_masked[190];
  assign N375 = N374 | data_masked[254];
  assign N374 = N373 | data_masked[318];
  assign N373 = N372 | data_masked[382];
  assign N372 = data_masked[510] | data_masked[446];
  assign data_o[63] = N383 | data_masked[63];
  assign N383 = N382 | data_masked[127];
  assign N382 = N381 | data_masked[191];
  assign N381 = N380 | data_masked[255];
  assign N380 = N379 | data_masked[319];
  assign N379 = N378 | data_masked[383];
  assign N378 = data_masked[511] | data_masked[447];

endmodule



module bsg_mux_00000040_00000001
(
  data_i,
  sel_i,
  data_o
);

  input [63:0] data_i;
  input [0:0] sel_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  assign data_o[63] = data_i[63];
  assign data_o[62] = data_i[62];
  assign data_o[61] = data_i[61];
  assign data_o[60] = data_i[60];
  assign data_o[59] = data_i[59];
  assign data_o[58] = data_i[58];
  assign data_o[57] = data_i[57];
  assign data_o[56] = data_i[56];
  assign data_o[55] = data_i[55];
  assign data_o[54] = data_i[54];
  assign data_o[53] = data_i[53];
  assign data_o[52] = data_i[52];
  assign data_o[51] = data_i[51];
  assign data_o[50] = data_i[50];
  assign data_o[49] = data_i[49];
  assign data_o[48] = data_i[48];
  assign data_o[47] = data_i[47];
  assign data_o[46] = data_i[46];
  assign data_o[45] = data_i[45];
  assign data_o[44] = data_i[44];
  assign data_o[43] = data_i[43];
  assign data_o[42] = data_i[42];
  assign data_o[41] = data_i[41];
  assign data_o[40] = data_i[40];
  assign data_o[39] = data_i[39];
  assign data_o[38] = data_i[38];
  assign data_o[37] = data_i[37];
  assign data_o[36] = data_i[36];
  assign data_o[35] = data_i[35];
  assign data_o[34] = data_i[34];
  assign data_o[33] = data_i[33];
  assign data_o[32] = data_i[32];
  assign data_o[31] = data_i[31];
  assign data_o[30] = data_i[30];
  assign data_o[29] = data_i[29];
  assign data_o[28] = data_i[28];
  assign data_o[27] = data_i[27];
  assign data_o[26] = data_i[26];
  assign data_o[25] = data_i[25];
  assign data_o[24] = data_i[24];
  assign data_o[23] = data_i[23];
  assign data_o[22] = data_i[22];
  assign data_o[21] = data_i[21];
  assign data_o[20] = data_i[20];
  assign data_o[19] = data_i[19];
  assign data_o[18] = data_i[18];
  assign data_o[17] = data_i[17];
  assign data_o[16] = data_i[16];
  assign data_o[15] = data_i[15];
  assign data_o[14] = data_i[14];
  assign data_o[13] = data_i[13];
  assign data_o[12] = data_i[12];
  assign data_o[11] = data_i[11];
  assign data_o[10] = data_i[10];
  assign data_o[9] = data_i[9];
  assign data_o[8] = data_i[8];
  assign data_o[7] = data_i[7];
  assign data_o[6] = data_i[6];
  assign data_o[5] = data_i[5];
  assign data_o[4] = data_i[4];
  assign data_o[3] = data_i[3];
  assign data_o[2] = data_i[2];
  assign data_o[1] = data_i[1];
  assign data_o[0] = data_i[0];

endmodule



module bsg_mem_1rw_sync_mask_write_bit_0000000f_00000040_1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [14:0] data_i;
  input [5:0] addr_i;
  input [14:0] w_mask_i;
  output [14:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [14:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_mux_width_p1_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [1:0] data_i;
  input [0:0] sel_i;
  output [0:0] data_o;
  wire [0:0] data_o;
  wire N0,N1;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[1] : 1'b0;
  assign N0 = sel_i[0];
  assign N1 = ~sel_i[0];

endmodule



module bsg_mux_width_p1_els_p4
(
  data_i,
  sel_i,
  data_o
);

  input [3:0] data_i;
  input [1:0] sel_i;
  output [0:0] data_o;
  wire [0:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[1] : 
                     (N3)? data_i[2] : 
                     (N5)? data_i[3] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_lru_pseudo_tree_encode_00000008
(
  lru_i,
  way_id_o
);

  input [6:0] lru_i;
  output [2:0] way_id_o;
  wire [2:0] way_id_o;
  wire way_id_o_2_;
  assign way_id_o_2_ = lru_i[0];
  assign way_id_o[2] = way_id_o_2_;

  bsg_mux_width_p1_els_p2
  \lru.rank_1_.nz.mux 
  (
    .data_i(lru_i[2:1]),
    .sel_i(way_id_o_2_),
    .data_o(way_id_o[1])
  );


  bsg_mux_width_p1_els_p4
  \lru.rank_2_.nz.mux 
  (
    .data_i(lru_i[6:3]),
    .sel_i({ way_id_o_2_, way_id_o[1:1] }),
    .data_o(way_id_o[0])
  );


endmodule



module bsg_expand_bitmask_in_width_p8_expand_p1
(
  i,
  o
);

  input [7:0] i;
  output [7:0] o;
  wire [7:0] o;
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_decode_num_out_p4
(
  i,
  o
);

  input [1:0] i;
  output [3:0] o;
  wire [3:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_expand_bitmask_in_width_p4_expand_p2
(
  i,
  o
);

  input [3:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire o_7_,o_5_,o_3_,o_1_;
  assign o_7_ = i[3];
  assign o[6] = o_7_;
  assign o[7] = o_7_;
  assign o_5_ = i[2];
  assign o[4] = o_5_;
  assign o[5] = o_5_;
  assign o_3_ = i[1];
  assign o[2] = o_3_;
  assign o[3] = o_3_;
  assign o_1_ = i[0];
  assign o[0] = o_1_;
  assign o[1] = o_1_;

endmodule



module bsg_decode_num_out_p2
(
  i,
  o
);

  input [0:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o = { 1'b0, 1'b1 } << i[0];

endmodule



module bsg_expand_bitmask_in_width_p2_expand_p4
(
  i,
  o
);

  input [1:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire o_7_,o_3_;
  assign o_7_ = i[1];
  assign o[4] = o_7_;
  assign o[5] = o_7_;
  assign o[6] = o_7_;
  assign o[7] = o_7_;
  assign o_3_ = i[0];
  assign o[0] = o_3_;
  assign o[1] = o_3_;
  assign o[2] = o_3_;
  assign o[3] = o_3_;

endmodule



module bsg_decode_num_out_p1
(
  i,
  o
);

  input [0:0] i;
  output [0:0] o;
  wire [0:0] o;
  assign o[0] = 1'b1;

endmodule



module bsg_expand_bitmask_in_width_p1_expand_p8
(
  i,
  o
);

  input [0:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire o_7_;
  assign o_7_ = i[0];
  assign o[0] = o_7_;
  assign o[1] = o_7_;
  assign o[2] = o_7_;
  assign o[3] = o_7_;
  assign o[4] = o_7_;
  assign o[5] = o_7_;
  assign o[6] = o_7_;
  assign o[7] = o_7_;

endmodule



module bsg_mux_one_hot_width_p64_els_p4
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [255:0] data_i;
  input [3:0] sel_one_hot_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127;
  wire [255:0] data_masked;
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[1];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[1];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[1];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[2];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[2];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[2];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[2];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[2];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[2];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[2];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[2];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[2];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[2];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[2];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[2];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[2];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[2];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[2];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[2];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[2];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[2];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[2];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[2];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[2];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[2];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[2];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[2];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[2];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[2];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[2];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[2];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[2];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[2];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[2];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[2];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[2];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[2];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[2];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[2];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[2];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[2];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[2];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[2];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[2];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[2];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[2];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[2];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[2];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[2];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[2];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[2];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[2];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[2];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[2];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[2];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[2];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[2];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[2];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[2];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[2];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[2];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[2];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[2];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[2];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[2];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[2];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[2];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[3];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[3];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[3];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[3];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[3];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[3];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[3];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[3];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[3];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[3];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[3];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[3];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[3];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[3];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[3];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[3];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[3];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[3];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[3];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[3];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[3];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[3];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[3];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[3];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[3];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[3];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[3];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[3];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[3];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[3];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[3];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[3];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[3];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[3];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[3];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[3];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[3];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[3];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[3];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[3];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[3];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[3];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[3];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[3];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[3];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[3];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[3];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[3];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[3];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[3];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[3];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[3];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[3];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[3];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[3];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[3];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[3];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[3];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[3];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[3];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[3];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[3];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[3];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[3];
  assign data_o[0] = N1 | data_masked[0];
  assign N1 = N0 | data_masked[64];
  assign N0 = data_masked[192] | data_masked[128];
  assign data_o[1] = N3 | data_masked[1];
  assign N3 = N2 | data_masked[65];
  assign N2 = data_masked[193] | data_masked[129];
  assign data_o[2] = N5 | data_masked[2];
  assign N5 = N4 | data_masked[66];
  assign N4 = data_masked[194] | data_masked[130];
  assign data_o[3] = N7 | data_masked[3];
  assign N7 = N6 | data_masked[67];
  assign N6 = data_masked[195] | data_masked[131];
  assign data_o[4] = N9 | data_masked[4];
  assign N9 = N8 | data_masked[68];
  assign N8 = data_masked[196] | data_masked[132];
  assign data_o[5] = N11 | data_masked[5];
  assign N11 = N10 | data_masked[69];
  assign N10 = data_masked[197] | data_masked[133];
  assign data_o[6] = N13 | data_masked[6];
  assign N13 = N12 | data_masked[70];
  assign N12 = data_masked[198] | data_masked[134];
  assign data_o[7] = N15 | data_masked[7];
  assign N15 = N14 | data_masked[71];
  assign N14 = data_masked[199] | data_masked[135];
  assign data_o[8] = N17 | data_masked[8];
  assign N17 = N16 | data_masked[72];
  assign N16 = data_masked[200] | data_masked[136];
  assign data_o[9] = N19 | data_masked[9];
  assign N19 = N18 | data_masked[73];
  assign N18 = data_masked[201] | data_masked[137];
  assign data_o[10] = N21 | data_masked[10];
  assign N21 = N20 | data_masked[74];
  assign N20 = data_masked[202] | data_masked[138];
  assign data_o[11] = N23 | data_masked[11];
  assign N23 = N22 | data_masked[75];
  assign N22 = data_masked[203] | data_masked[139];
  assign data_o[12] = N25 | data_masked[12];
  assign N25 = N24 | data_masked[76];
  assign N24 = data_masked[204] | data_masked[140];
  assign data_o[13] = N27 | data_masked[13];
  assign N27 = N26 | data_masked[77];
  assign N26 = data_masked[205] | data_masked[141];
  assign data_o[14] = N29 | data_masked[14];
  assign N29 = N28 | data_masked[78];
  assign N28 = data_masked[206] | data_masked[142];
  assign data_o[15] = N31 | data_masked[15];
  assign N31 = N30 | data_masked[79];
  assign N30 = data_masked[207] | data_masked[143];
  assign data_o[16] = N33 | data_masked[16];
  assign N33 = N32 | data_masked[80];
  assign N32 = data_masked[208] | data_masked[144];
  assign data_o[17] = N35 | data_masked[17];
  assign N35 = N34 | data_masked[81];
  assign N34 = data_masked[209] | data_masked[145];
  assign data_o[18] = N37 | data_masked[18];
  assign N37 = N36 | data_masked[82];
  assign N36 = data_masked[210] | data_masked[146];
  assign data_o[19] = N39 | data_masked[19];
  assign N39 = N38 | data_masked[83];
  assign N38 = data_masked[211] | data_masked[147];
  assign data_o[20] = N41 | data_masked[20];
  assign N41 = N40 | data_masked[84];
  assign N40 = data_masked[212] | data_masked[148];
  assign data_o[21] = N43 | data_masked[21];
  assign N43 = N42 | data_masked[85];
  assign N42 = data_masked[213] | data_masked[149];
  assign data_o[22] = N45 | data_masked[22];
  assign N45 = N44 | data_masked[86];
  assign N44 = data_masked[214] | data_masked[150];
  assign data_o[23] = N47 | data_masked[23];
  assign N47 = N46 | data_masked[87];
  assign N46 = data_masked[215] | data_masked[151];
  assign data_o[24] = N49 | data_masked[24];
  assign N49 = N48 | data_masked[88];
  assign N48 = data_masked[216] | data_masked[152];
  assign data_o[25] = N51 | data_masked[25];
  assign N51 = N50 | data_masked[89];
  assign N50 = data_masked[217] | data_masked[153];
  assign data_o[26] = N53 | data_masked[26];
  assign N53 = N52 | data_masked[90];
  assign N52 = data_masked[218] | data_masked[154];
  assign data_o[27] = N55 | data_masked[27];
  assign N55 = N54 | data_masked[91];
  assign N54 = data_masked[219] | data_masked[155];
  assign data_o[28] = N57 | data_masked[28];
  assign N57 = N56 | data_masked[92];
  assign N56 = data_masked[220] | data_masked[156];
  assign data_o[29] = N59 | data_masked[29];
  assign N59 = N58 | data_masked[93];
  assign N58 = data_masked[221] | data_masked[157];
  assign data_o[30] = N61 | data_masked[30];
  assign N61 = N60 | data_masked[94];
  assign N60 = data_masked[222] | data_masked[158];
  assign data_o[31] = N63 | data_masked[31];
  assign N63 = N62 | data_masked[95];
  assign N62 = data_masked[223] | data_masked[159];
  assign data_o[32] = N65 | data_masked[32];
  assign N65 = N64 | data_masked[96];
  assign N64 = data_masked[224] | data_masked[160];
  assign data_o[33] = N67 | data_masked[33];
  assign N67 = N66 | data_masked[97];
  assign N66 = data_masked[225] | data_masked[161];
  assign data_o[34] = N69 | data_masked[34];
  assign N69 = N68 | data_masked[98];
  assign N68 = data_masked[226] | data_masked[162];
  assign data_o[35] = N71 | data_masked[35];
  assign N71 = N70 | data_masked[99];
  assign N70 = data_masked[227] | data_masked[163];
  assign data_o[36] = N73 | data_masked[36];
  assign N73 = N72 | data_masked[100];
  assign N72 = data_masked[228] | data_masked[164];
  assign data_o[37] = N75 | data_masked[37];
  assign N75 = N74 | data_masked[101];
  assign N74 = data_masked[229] | data_masked[165];
  assign data_o[38] = N77 | data_masked[38];
  assign N77 = N76 | data_masked[102];
  assign N76 = data_masked[230] | data_masked[166];
  assign data_o[39] = N79 | data_masked[39];
  assign N79 = N78 | data_masked[103];
  assign N78 = data_masked[231] | data_masked[167];
  assign data_o[40] = N81 | data_masked[40];
  assign N81 = N80 | data_masked[104];
  assign N80 = data_masked[232] | data_masked[168];
  assign data_o[41] = N83 | data_masked[41];
  assign N83 = N82 | data_masked[105];
  assign N82 = data_masked[233] | data_masked[169];
  assign data_o[42] = N85 | data_masked[42];
  assign N85 = N84 | data_masked[106];
  assign N84 = data_masked[234] | data_masked[170];
  assign data_o[43] = N87 | data_masked[43];
  assign N87 = N86 | data_masked[107];
  assign N86 = data_masked[235] | data_masked[171];
  assign data_o[44] = N89 | data_masked[44];
  assign N89 = N88 | data_masked[108];
  assign N88 = data_masked[236] | data_masked[172];
  assign data_o[45] = N91 | data_masked[45];
  assign N91 = N90 | data_masked[109];
  assign N90 = data_masked[237] | data_masked[173];
  assign data_o[46] = N93 | data_masked[46];
  assign N93 = N92 | data_masked[110];
  assign N92 = data_masked[238] | data_masked[174];
  assign data_o[47] = N95 | data_masked[47];
  assign N95 = N94 | data_masked[111];
  assign N94 = data_masked[239] | data_masked[175];
  assign data_o[48] = N97 | data_masked[48];
  assign N97 = N96 | data_masked[112];
  assign N96 = data_masked[240] | data_masked[176];
  assign data_o[49] = N99 | data_masked[49];
  assign N99 = N98 | data_masked[113];
  assign N98 = data_masked[241] | data_masked[177];
  assign data_o[50] = N101 | data_masked[50];
  assign N101 = N100 | data_masked[114];
  assign N100 = data_masked[242] | data_masked[178];
  assign data_o[51] = N103 | data_masked[51];
  assign N103 = N102 | data_masked[115];
  assign N102 = data_masked[243] | data_masked[179];
  assign data_o[52] = N105 | data_masked[52];
  assign N105 = N104 | data_masked[116];
  assign N104 = data_masked[244] | data_masked[180];
  assign data_o[53] = N107 | data_masked[53];
  assign N107 = N106 | data_masked[117];
  assign N106 = data_masked[245] | data_masked[181];
  assign data_o[54] = N109 | data_masked[54];
  assign N109 = N108 | data_masked[118];
  assign N108 = data_masked[246] | data_masked[182];
  assign data_o[55] = N111 | data_masked[55];
  assign N111 = N110 | data_masked[119];
  assign N110 = data_masked[247] | data_masked[183];
  assign data_o[56] = N113 | data_masked[56];
  assign N113 = N112 | data_masked[120];
  assign N112 = data_masked[248] | data_masked[184];
  assign data_o[57] = N115 | data_masked[57];
  assign N115 = N114 | data_masked[121];
  assign N114 = data_masked[249] | data_masked[185];
  assign data_o[58] = N117 | data_masked[58];
  assign N117 = N116 | data_masked[122];
  assign N116 = data_masked[250] | data_masked[186];
  assign data_o[59] = N119 | data_masked[59];
  assign N119 = N118 | data_masked[123];
  assign N118 = data_masked[251] | data_masked[187];
  assign data_o[60] = N121 | data_masked[60];
  assign N121 = N120 | data_masked[124];
  assign N120 = data_masked[252] | data_masked[188];
  assign data_o[61] = N123 | data_masked[61];
  assign N123 = N122 | data_masked[125];
  assign N122 = data_masked[253] | data_masked[189];
  assign data_o[62] = N125 | data_masked[62];
  assign N125 = N124 | data_masked[126];
  assign N124 = data_masked[254] | data_masked[190];
  assign data_o[63] = N127 | data_masked[63];
  assign N127 = N126 | data_masked[127];
  assign N126 = data_masked[255] | data_masked[191];

endmodule



module bsg_mux_one_hot_00000008_4
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [31:0] data_i;
  input [3:0] sel_one_hot_i;
  output [7:0] data_o;
  wire [7:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;
  wire [31:0] data_masked;
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[1];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[1];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[1];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[1];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[1];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[1];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[1];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[1];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[2];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[2];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[2];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[2];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[2];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[2];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[2];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[2];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[3];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[3];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[3];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[3];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[3];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[3];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[3];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[3];
  assign data_o[0] = N1 | data_masked[0];
  assign N1 = N0 | data_masked[8];
  assign N0 = data_masked[24] | data_masked[16];
  assign data_o[1] = N3 | data_masked[1];
  assign N3 = N2 | data_masked[9];
  assign N2 = data_masked[25] | data_masked[17];
  assign data_o[2] = N5 | data_masked[2];
  assign N5 = N4 | data_masked[10];
  assign N4 = data_masked[26] | data_masked[18];
  assign data_o[3] = N7 | data_masked[3];
  assign N7 = N6 | data_masked[11];
  assign N6 = data_masked[27] | data_masked[19];
  assign data_o[4] = N9 | data_masked[4];
  assign N9 = N8 | data_masked[12];
  assign N8 = data_masked[28] | data_masked[20];
  assign data_o[5] = N11 | data_masked[5];
  assign N11 = N10 | data_masked[13];
  assign N10 = data_masked[29] | data_masked[21];
  assign data_o[6] = N13 | data_masked[6];
  assign N13 = N12 | data_masked[14];
  assign N12 = data_masked[30] | data_masked[22];
  assign data_o[7] = N15 | data_masked[7];
  assign N15 = N14 | data_masked[15];
  assign N14 = data_masked[31] | data_masked[23];

endmodule



module bsg_counter_up_down_max_val_p2_init_val_p0_max_step_p1
(
  clk_i,
  reset_i,
  up_i,
  down_i,
  count_o
);

  input [0:0] up_i;
  input [0:0] down_i;
  output [1:0] count_o;
  input clk_i;
  input reset_i;
  wire [1:0] count_o;
  wire N0,N1,N2,N3,N4;
  reg count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign { N2, N1 } = count_o - down_i[0];
  assign { N4, N3 } = { N2, N1 } + up_i[0];
  assign N0 = ~reset_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      count_o_1_sv2v_reg <= 1'b0;
      count_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      count_o_1_sv2v_reg <= N4;
      count_o_0_sv2v_reg <= N3;
    end 
  end


endmodule



module bsg_dff_en_width_p113
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [112:0] data_i;
  output [112:0] data_o;
  input clk_i;
  input en_i;
  wire [112:0] data_o;
  reg data_o_112_sv2v_reg,data_o_111_sv2v_reg,data_o_110_sv2v_reg,data_o_109_sv2v_reg,
  data_o_108_sv2v_reg,data_o_107_sv2v_reg,data_o_106_sv2v_reg,data_o_105_sv2v_reg,
  data_o_104_sv2v_reg,data_o_103_sv2v_reg,data_o_102_sv2v_reg,data_o_101_sv2v_reg,
  data_o_100_sv2v_reg,data_o_99_sv2v_reg,data_o_98_sv2v_reg,data_o_97_sv2v_reg,
  data_o_96_sv2v_reg,data_o_95_sv2v_reg,data_o_94_sv2v_reg,data_o_93_sv2v_reg,
  data_o_92_sv2v_reg,data_o_91_sv2v_reg,data_o_90_sv2v_reg,data_o_89_sv2v_reg,
  data_o_88_sv2v_reg,data_o_87_sv2v_reg,data_o_86_sv2v_reg,data_o_85_sv2v_reg,
  data_o_84_sv2v_reg,data_o_83_sv2v_reg,data_o_82_sv2v_reg,data_o_81_sv2v_reg,data_o_80_sv2v_reg,
  data_o_79_sv2v_reg,data_o_78_sv2v_reg,data_o_77_sv2v_reg,data_o_76_sv2v_reg,
  data_o_75_sv2v_reg,data_o_74_sv2v_reg,data_o_73_sv2v_reg,data_o_72_sv2v_reg,
  data_o_71_sv2v_reg,data_o_70_sv2v_reg,data_o_69_sv2v_reg,data_o_68_sv2v_reg,
  data_o_67_sv2v_reg,data_o_66_sv2v_reg,data_o_65_sv2v_reg,data_o_64_sv2v_reg,
  data_o_63_sv2v_reg,data_o_62_sv2v_reg,data_o_61_sv2v_reg,data_o_60_sv2v_reg,data_o_59_sv2v_reg,
  data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,data_o_55_sv2v_reg,
  data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,data_o_51_sv2v_reg,
  data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,data_o_47_sv2v_reg,
  data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,data_o_43_sv2v_reg,
  data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,
  data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,
  data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,
  data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,
  data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,
  data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,
  data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,
  data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,
  data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[112] = data_o_112_sv2v_reg;
  assign data_o[111] = data_o_111_sv2v_reg;
  assign data_o[110] = data_o_110_sv2v_reg;
  assign data_o[109] = data_o_109_sv2v_reg;
  assign data_o[108] = data_o_108_sv2v_reg;
  assign data_o[107] = data_o_107_sv2v_reg;
  assign data_o[106] = data_o_106_sv2v_reg;
  assign data_o[105] = data_o_105_sv2v_reg;
  assign data_o[104] = data_o_104_sv2v_reg;
  assign data_o[103] = data_o_103_sv2v_reg;
  assign data_o[102] = data_o_102_sv2v_reg;
  assign data_o[101] = data_o_101_sv2v_reg;
  assign data_o[100] = data_o_100_sv2v_reg;
  assign data_o[99] = data_o_99_sv2v_reg;
  assign data_o[98] = data_o_98_sv2v_reg;
  assign data_o[97] = data_o_97_sv2v_reg;
  assign data_o[96] = data_o_96_sv2v_reg;
  assign data_o[95] = data_o_95_sv2v_reg;
  assign data_o[94] = data_o_94_sv2v_reg;
  assign data_o[93] = data_o_93_sv2v_reg;
  assign data_o[92] = data_o_92_sv2v_reg;
  assign data_o[91] = data_o_91_sv2v_reg;
  assign data_o[90] = data_o_90_sv2v_reg;
  assign data_o[89] = data_o_89_sv2v_reg;
  assign data_o[88] = data_o_88_sv2v_reg;
  assign data_o[87] = data_o_87_sv2v_reg;
  assign data_o[86] = data_o_86_sv2v_reg;
  assign data_o[85] = data_o_85_sv2v_reg;
  assign data_o[84] = data_o_84_sv2v_reg;
  assign data_o[83] = data_o_83_sv2v_reg;
  assign data_o[82] = data_o_82_sv2v_reg;
  assign data_o[81] = data_o_81_sv2v_reg;
  assign data_o[80] = data_o_80_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_112_sv2v_reg <= data_i[112];
      data_o_111_sv2v_reg <= data_i[111];
      data_o_110_sv2v_reg <= data_i[110];
      data_o_109_sv2v_reg <= data_i[109];
      data_o_108_sv2v_reg <= data_i[108];
      data_o_107_sv2v_reg <= data_i[107];
      data_o_106_sv2v_reg <= data_i[106];
      data_o_105_sv2v_reg <= data_i[105];
      data_o_104_sv2v_reg <= data_i[104];
      data_o_103_sv2v_reg <= data_i[103];
      data_o_102_sv2v_reg <= data_i[102];
      data_o_101_sv2v_reg <= data_i[101];
      data_o_100_sv2v_reg <= data_i[100];
      data_o_99_sv2v_reg <= data_i[99];
      data_o_98_sv2v_reg <= data_i[98];
      data_o_97_sv2v_reg <= data_i[97];
      data_o_96_sv2v_reg <= data_i[96];
      data_o_95_sv2v_reg <= data_i[95];
      data_o_94_sv2v_reg <= data_i[94];
      data_o_93_sv2v_reg <= data_i[93];
      data_o_92_sv2v_reg <= data_i[92];
      data_o_91_sv2v_reg <= data_i[91];
      data_o_90_sv2v_reg <= data_i[90];
      data_o_89_sv2v_reg <= data_i[89];
      data_o_88_sv2v_reg <= data_i[88];
      data_o_87_sv2v_reg <= data_i[87];
      data_o_86_sv2v_reg <= data_i[86];
      data_o_85_sv2v_reg <= data_i[85];
      data_o_84_sv2v_reg <= data_i[84];
      data_o_83_sv2v_reg <= data_i[83];
      data_o_82_sv2v_reg <= data_i[82];
      data_o_81_sv2v_reg <= data_i[81];
      data_o_80_sv2v_reg <= data_i[80];
      data_o_79_sv2v_reg <= data_i[79];
      data_o_78_sv2v_reg <= data_i[78];
      data_o_77_sv2v_reg <= data_i[77];
      data_o_76_sv2v_reg <= data_i[76];
      data_o_75_sv2v_reg <= data_i[75];
      data_o_74_sv2v_reg <= data_i[74];
      data_o_73_sv2v_reg <= data_i[73];
      data_o_72_sv2v_reg <= data_i[72];
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mux_segmented_segments_p8_segment_width_p8
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [63:0] data0_i;
  input [63:0] data1_i;
  input [7:0] sel_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;
  assign data_o[7:0] = (N0)? data1_i[7:0] : 
                       (N8)? data0_i[7:0] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[15:8] = (N1)? data1_i[15:8] : 
                        (N9)? data0_i[15:8] : 1'b0;
  assign N1 = sel_i[1];
  assign data_o[23:16] = (N2)? data1_i[23:16] : 
                         (N10)? data0_i[23:16] : 1'b0;
  assign N2 = sel_i[2];
  assign data_o[31:24] = (N3)? data1_i[31:24] : 
                         (N11)? data0_i[31:24] : 1'b0;
  assign N3 = sel_i[3];
  assign data_o[39:32] = (N4)? data1_i[39:32] : 
                         (N12)? data0_i[39:32] : 1'b0;
  assign N4 = sel_i[4];
  assign data_o[47:40] = (N5)? data1_i[47:40] : 
                         (N13)? data0_i[47:40] : 1'b0;
  assign N5 = sel_i[5];
  assign data_o[55:48] = (N6)? data1_i[55:48] : 
                         (N14)? data0_i[55:48] : 1'b0;
  assign N6 = sel_i[6];
  assign data_o[63:56] = (N7)? data1_i[63:56] : 
                         (N15)? data0_i[63:56] : 1'b0;
  assign N7 = sel_i[7];
  assign N8 = ~sel_i[0];
  assign N9 = ~sel_i[1];
  assign N10 = ~sel_i[2];
  assign N11 = ~sel_i[3];
  assign N12 = ~sel_i[4];
  assign N13 = ~sel_i[5];
  assign N14 = ~sel_i[6];
  assign N15 = ~sel_i[7];

endmodule



module bsg_dff_reset_width_p72
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [71:0] data_i;
  output [71:0] data_o;
  input clk_i;
  input reset_i;
  wire [71:0] data_o;
  reg data_o_71_sv2v_reg,data_o_70_sv2v_reg,data_o_69_sv2v_reg,data_o_68_sv2v_reg,
  data_o_67_sv2v_reg,data_o_66_sv2v_reg,data_o_65_sv2v_reg,data_o_64_sv2v_reg,
  data_o_63_sv2v_reg,data_o_62_sv2v_reg,data_o_61_sv2v_reg,data_o_60_sv2v_reg,
  data_o_59_sv2v_reg,data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,
  data_o_55_sv2v_reg,data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,data_o_51_sv2v_reg,
  data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,data_o_47_sv2v_reg,
  data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,data_o_43_sv2v_reg,
  data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,
  data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,
  data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,
  data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,
  data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,
  data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,
  data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,
  data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_71_sv2v_reg <= 1'b0;
      data_o_70_sv2v_reg <= 1'b0;
      data_o_69_sv2v_reg <= 1'b0;
      data_o_68_sv2v_reg <= 1'b0;
      data_o_67_sv2v_reg <= 1'b0;
      data_o_66_sv2v_reg <= 1'b0;
      data_o_65_sv2v_reg <= 1'b0;
      data_o_64_sv2v_reg <= 1'b0;
      data_o_63_sv2v_reg <= 1'b0;
      data_o_62_sv2v_reg <= 1'b0;
      data_o_61_sv2v_reg <= 1'b0;
      data_o_60_sv2v_reg <= 1'b0;
      data_o_59_sv2v_reg <= 1'b0;
      data_o_58_sv2v_reg <= 1'b0;
      data_o_57_sv2v_reg <= 1'b0;
      data_o_56_sv2v_reg <= 1'b0;
      data_o_55_sv2v_reg <= 1'b0;
      data_o_54_sv2v_reg <= 1'b0;
      data_o_53_sv2v_reg <= 1'b0;
      data_o_52_sv2v_reg <= 1'b0;
      data_o_51_sv2v_reg <= 1'b0;
      data_o_50_sv2v_reg <= 1'b0;
      data_o_49_sv2v_reg <= 1'b0;
      data_o_48_sv2v_reg <= 1'b0;
      data_o_47_sv2v_reg <= 1'b0;
      data_o_46_sv2v_reg <= 1'b0;
      data_o_45_sv2v_reg <= 1'b0;
      data_o_44_sv2v_reg <= 1'b0;
      data_o_43_sv2v_reg <= 1'b0;
      data_o_42_sv2v_reg <= 1'b0;
      data_o_41_sv2v_reg <= 1'b0;
      data_o_40_sv2v_reg <= 1'b0;
      data_o_39_sv2v_reg <= 1'b0;
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bp_be_dcache_wbuf_00_00000040_00000008_00000200_00000080_00000014
(
  clk_i,
  reset_i,
  wbuf_entry_i,
  v_i,
  wbuf_entry_o,
  v_o,
  force_o,
  yumi_i,
  data_mem_pkt_i,
  data_mem_pkt_v_i,
  tag_mem_pkt_i,
  tag_mem_pkt_v_i,
  stat_mem_pkt_i,
  stat_mem_pkt_v_i,
  snoop_match_o,
  v_tl_i,
  addr_tl_i,
  data_tv_i,
  data_merged_o
);

  input [112:0] wbuf_entry_i;
  output [112:0] wbuf_entry_o;
  input [142:0] data_mem_pkt_i;
  input [34:0] tag_mem_pkt_i;
  input [10:0] stat_mem_pkt_i;
  input [31:0] addr_tl_i;
  input [63:0] data_tv_i;
  output [63:0] data_merged_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input data_mem_pkt_v_i;
  input tag_mem_pkt_v_i;
  input stat_mem_pkt_v_i;
  input v_tl_i;
  output v_o;
  output force_o;
  output snoop_match_o;
  wire [112:0] wbuf_entry_o,wbuf_entry_el0_r,wbuf_entry_el1_n,wbuf_entry_el1_r;
  wire [63:0] data_merged_o,el0or1_data,bypass_data_n,bypass_data_r;
  wire v_o,force_o,snoop_match_o,N0,N1,N2,N3,N4,N5,N6,N7,el0_valid,el1_valid,
  el0_enable,N8,el1_enable,mux1_sel,N9,N10,N11,N12,N13,N14,N15,N16,tag_hit0_n,tag_hit1_n,
  tag_hit2_n,_2_net__7_,_2_net__6_,_2_net__5_,_2_net__4_,_2_net__3_,_2_net__2_,
  _2_net__1_,_2_net__0_,_4_net__7_,_4_net__6_,_4_net__5_,_4_net__4_,_4_net__3_,
  _4_net__2_,_4_net__1_,_4_net__0_,N17,snoop_tag_match,N18,snoop_stat_match,N19,
  snoop_el0_match,N20,snoop_el1_match,N21,snoop_el2_match,N22,N23,N24,N25,N26,N27,N28,N29,
  N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,
  N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,
  N70,N71,N72,N73,N74,N75;
  wire [1:0] num_els_r;
  wire [7:7] tag_hit0x4,tag_hit1x4,tag_hit2x4;
  wire [7:0] bypass_mask_n,bypass_mask_r;

  bsg_counter_up_down_max_val_p2_init_val_p0_max_step_p1
  num_els_counter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .up_i(v_i),
    .down_i(yumi_i),
    .count_o(num_els_r)
  );


  bsg_dff_en_width_p113
  wbuf_entry0_reg
  (
    .clk_i(clk_i),
    .data_i(wbuf_entry_i),
    .en_i(el0_enable),
    .data_o(wbuf_entry_el0_r)
  );


  bsg_dff_en_width_p113
  wbuf_entry1_reg
  (
    .clk_i(clk_i),
    .data_i(wbuf_entry_el1_n),
    .en_i(el1_enable),
    .data_o(wbuf_entry_el1_r)
  );

  assign tag_hit0_n = addr_tl_i[31:3] == wbuf_entry_el0_r[31:3];
  assign tag_hit1_n = addr_tl_i[31:3] == wbuf_entry_el1_r[31:3];
  assign tag_hit2_n = addr_tl_i[31:3] == wbuf_entry_i[31:3];

  bsg_mux_segmented_segments_p8_segment_width_p8
  mux_segmented_merge0
  (
    .data0_i(wbuf_entry_el1_r[95:32]),
    .data1_i(wbuf_entry_el0_r[95:32]),
    .sel_i({ _2_net__7_, _2_net__6_, _2_net__5_, _2_net__4_, _2_net__3_, _2_net__2_, _2_net__1_, _2_net__0_ }),
    .data_o(el0or1_data)
  );


  bsg_mux_segmented_segments_p8_segment_width_p8
  mux_segmented_merge1
  (
    .data0_i(el0or1_data),
    .data1_i(wbuf_entry_i[95:32]),
    .sel_i({ _4_net__7_, _4_net__6_, _4_net__5_, _4_net__4_, _4_net__3_, _4_net__2_, _4_net__1_, _4_net__0_ }),
    .data_o(bypass_data_n)
  );


  bsg_dff_reset_width_p72
  bypass_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ bypass_mask_n, bypass_data_n }),
    .data_o({ bypass_mask_r, bypass_data_r })
  );


  bsg_mux_segmented_segments_p8_segment_width_p8
  bypass_mux_segmented
  (
    .data0_i(data_tv_i),
    .data1_i(bypass_data_r),
    .sel_i(bypass_mask_r),
    .data_o(data_merged_o)
  );

  assign N17 = addr_tl_i[11:6] == tag_mem_pkt_i[34:29];
  assign N18 = addr_tl_i[11:6] == stat_mem_pkt_i[10:5];
  assign N19 = wbuf_entry_el0_r[11:6] == data_mem_pkt_i[142:137];
  assign N20 = wbuf_entry_el1_r[11:6] == data_mem_pkt_i[142:137];
  assign N21 = wbuf_entry_i[11:6] == data_mem_pkt_i[142:137];
  assign N22 = ~num_els_r[1];
  assign N23 = num_els_r[0] | N22;
  assign N24 = ~N23;
  assign N11 = (N0)? v_i : 
               (N1)? 1'b1 : 1'b0;
  assign N0 = N7;
  assign N1 = num_els_r[0];
  assign N12 = (N0)? 1'b0 : 
               (N1)? N9 : 1'b0;
  assign N13 = (N0)? N8 : 
               (N1)? N10 : 1'b0;
  assign mux1_sel = (N2)? num_els_r[0] : 
                    (N3)? 1'b1 : 1'b0;
  assign N2 = N22;
  assign N3 = el0_valid;
  assign v_o = (N2)? N11 : 
               (N3)? 1'b1 : 1'b0;
  assign el1_valid = (N2)? num_els_r[0] : 
                     (N3)? 1'b1 : 1'b0;
  assign el0_enable = (N2)? N12 : 
                      (N3)? N14 : 1'b0;
  assign el1_enable = (N2)? N13 : 
                      (N3)? yumi_i : 1'b0;
  assign wbuf_entry_el1_n = (N3)? wbuf_entry_el0_r : 
                            (N4)? wbuf_entry_i : 1'b0;
  assign N4 = N15;
  assign wbuf_entry_o = (N5)? wbuf_entry_el1_r : 
                        (N6)? wbuf_entry_i : 1'b0;
  assign N5 = mux1_sel;
  assign N6 = N16;
  assign el0_valid = num_els_r[1];
  assign N7 = ~num_els_r[0];
  assign N8 = v_i & N25;
  assign N25 = ~yumi_i;
  assign N9 = v_i & N26;
  assign N26 = ~yumi_i;
  assign N10 = v_i & yumi_i;
  assign N14 = v_i & yumi_i;
  assign force_o = v_i & N24;
  assign N15 = ~el0_valid;
  assign N16 = ~mux1_sel;
  assign tag_hit0x4[7] = N27 & el0_valid;
  assign N27 = v_tl_i & tag_hit0_n;
  assign tag_hit1x4[7] = N28 & el1_valid;
  assign N28 = v_tl_i & tag_hit1_n;
  assign tag_hit2x4[7] = N29 & v_i;
  assign N29 = v_tl_i & tag_hit2_n;
  assign _2_net__7_ = tag_hit0x4[7] & wbuf_entry_el0_r[103];
  assign _2_net__6_ = tag_hit0x4[7] & wbuf_entry_el0_r[102];
  assign _2_net__5_ = tag_hit0x4[7] & wbuf_entry_el0_r[101];
  assign _2_net__4_ = tag_hit0x4[7] & wbuf_entry_el0_r[100];
  assign _2_net__3_ = tag_hit0x4[7] & wbuf_entry_el0_r[99];
  assign _2_net__2_ = tag_hit0x4[7] & wbuf_entry_el0_r[98];
  assign _2_net__1_ = tag_hit0x4[7] & wbuf_entry_el0_r[97];
  assign _2_net__0_ = tag_hit0x4[7] & wbuf_entry_el0_r[96];
  assign _4_net__7_ = tag_hit2x4[7] & wbuf_entry_i[103];
  assign _4_net__6_ = tag_hit2x4[7] & wbuf_entry_i[102];
  assign _4_net__5_ = tag_hit2x4[7] & wbuf_entry_i[101];
  assign _4_net__4_ = tag_hit2x4[7] & wbuf_entry_i[100];
  assign _4_net__3_ = tag_hit2x4[7] & wbuf_entry_i[99];
  assign _4_net__2_ = tag_hit2x4[7] & wbuf_entry_i[98];
  assign _4_net__1_ = tag_hit2x4[7] & wbuf_entry_i[97];
  assign _4_net__0_ = tag_hit2x4[7] & wbuf_entry_i[96];
  assign bypass_mask_n[7] = N32 | N33;
  assign N32 = N30 | N31;
  assign N30 = tag_hit0x4[7] & wbuf_entry_el0_r[103];
  assign N31 = tag_hit1x4[7] & wbuf_entry_el1_r[103];
  assign N33 = tag_hit2x4[7] & wbuf_entry_i[103];
  assign bypass_mask_n[6] = N36 | N37;
  assign N36 = N34 | N35;
  assign N34 = tag_hit0x4[7] & wbuf_entry_el0_r[102];
  assign N35 = tag_hit1x4[7] & wbuf_entry_el1_r[102];
  assign N37 = tag_hit2x4[7] & wbuf_entry_i[102];
  assign bypass_mask_n[5] = N40 | N41;
  assign N40 = N38 | N39;
  assign N38 = tag_hit0x4[7] & wbuf_entry_el0_r[101];
  assign N39 = tag_hit1x4[7] & wbuf_entry_el1_r[101];
  assign N41 = tag_hit2x4[7] & wbuf_entry_i[101];
  assign bypass_mask_n[4] = N44 | N45;
  assign N44 = N42 | N43;
  assign N42 = tag_hit0x4[7] & wbuf_entry_el0_r[100];
  assign N43 = tag_hit1x4[7] & wbuf_entry_el1_r[100];
  assign N45 = tag_hit2x4[7] & wbuf_entry_i[100];
  assign bypass_mask_n[3] = N48 | N49;
  assign N48 = N46 | N47;
  assign N46 = tag_hit0x4[7] & wbuf_entry_el0_r[99];
  assign N47 = tag_hit1x4[7] & wbuf_entry_el1_r[99];
  assign N49 = tag_hit2x4[7] & wbuf_entry_i[99];
  assign bypass_mask_n[2] = N52 | N53;
  assign N52 = N50 | N51;
  assign N50 = tag_hit0x4[7] & wbuf_entry_el0_r[98];
  assign N51 = tag_hit1x4[7] & wbuf_entry_el1_r[98];
  assign N53 = tag_hit2x4[7] & wbuf_entry_i[98];
  assign bypass_mask_n[1] = N56 | N57;
  assign N56 = N54 | N55;
  assign N54 = tag_hit0x4[7] & wbuf_entry_el0_r[97];
  assign N55 = tag_hit1x4[7] & wbuf_entry_el1_r[97];
  assign N57 = tag_hit2x4[7] & wbuf_entry_i[97];
  assign bypass_mask_n[0] = N60 | N61;
  assign N60 = N58 | N59;
  assign N58 = tag_hit0x4[7] & wbuf_entry_el0_r[96];
  assign N59 = tag_hit1x4[7] & wbuf_entry_el1_r[96];
  assign N61 = tag_hit2x4[7] & wbuf_entry_i[96];
  assign snoop_tag_match = N62 & N17;
  assign N62 = v_tl_i & tag_mem_pkt_v_i;
  assign snoop_stat_match = N63 & N18;
  assign N63 = v_tl_i & stat_mem_pkt_v_i;
  assign snoop_el0_match = N66 & N19;
  assign N66 = N65 & data_mem_pkt_v_i;
  assign N65 = el0_valid & N64;
  assign N64 = ~wbuf_entry_i[112];
  assign snoop_el1_match = N69 & N20;
  assign N69 = N68 & data_mem_pkt_v_i;
  assign N68 = el1_valid & N67;
  assign N67 = ~wbuf_entry_el1_r[112];
  assign snoop_el2_match = N72 & N21;
  assign N72 = N71 & data_mem_pkt_v_i;
  assign N71 = v_i & N70;
  assign N70 = ~wbuf_entry_i[112];
  assign snoop_match_o = N75 | snoop_el2_match;
  assign N75 = N74 | snoop_el1_match;
  assign N74 = N73 | snoop_el0_match;
  assign N73 = snoop_tag_match | snoop_stat_match;

endmodule



module bsg_dff_0000000c
(
  clk_i,
  data_i,
  data_o
);

  input [11:0] data_i;
  output [11:0] data_o;
  input clk_i;
  wire [11:0] data_o;
  reg data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,
  data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_scan_00000008_1_1
(
  i,
  o
);

  input [7:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__7_,t_1__6_,
  t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__7_ = i[0] | 1'b0;
  assign t_1__6_ = i[1] | i[0];
  assign t_1__5_ = i[2] | i[1];
  assign t_1__4_ = i[3] | i[2];
  assign t_1__3_ = i[4] | i[3];
  assign t_1__2_ = i[5] | i[4];
  assign t_1__1_ = i[6] | i[5];
  assign t_1__0_ = i[7] | i[6];
  assign t_2__7_ = t_1__7_ | 1'b0;
  assign t_2__6_ = t_1__6_ | 1'b0;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign o[0] = t_2__7_ | 1'b0;
  assign o[1] = t_2__6_ | 1'b0;
  assign o[2] = t_2__5_ | 1'b0;
  assign o[3] = t_2__4_ | 1'b0;
  assign o[4] = t_2__3_ | t_2__7_;
  assign o[5] = t_2__2_ | t_2__6_;
  assign o[6] = t_2__1_ | t_2__5_;
  assign o[7] = t_2__0_ | t_2__4_;

endmodule



module bsg_priority_encode_one_hot_out_00000008_1
(
  i,
  o,
  v_o
);

  input [7:0] i;
  output [7:0] o;
  output v_o;
  wire [7:0] o;
  wire v_o,N0,N1,N2,N3,N4,N5,N6;
  wire [6:1] scan_lo;

  bsg_scan_00000008_1_1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, scan_lo, o[0:0] })
  );

  assign o[7] = v_o & N0;
  assign N0 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N1;
  assign N1 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N2;
  assign N2 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N3;
  assign N3 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N4;
  assign N4 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N5;
  assign N5 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N6;
  assign N6 = ~o[0];

endmodule



module bsg_priority_encode_00000008_1
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [7:0] enc_lo;

  bsg_priority_encode_one_hot_out_00000008_1
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_00000008_1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o)
  );


endmodule



module bsg_dff_00000003
(
  clk_i,
  data_i,
  data_o
);

  input [2:0] data_i;
  output [2:0] data_o;
  input clk_i;
  wire [2:0] data_o;
  reg data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_rotate_left_00000008
(
  data_i,
  rot_i,
  o
);

  input [7:0] data_i;
  input [2:0] rot_i;
  output [7:0] o;
  wire [7:0] o;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7;
  assign { o, sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7 } = { data_i, data_i[7:1] } << rot_i;

endmodule



module bsg_rotate_left_00000080
(
  data_i,
  rot_i,
  o
);

  input [127:0] data_i;
  input [6:0] rot_i;
  output [127:0] o;
  wire [127:0] o;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,
  sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,
  sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,sv2v_dc_21,sv2v_dc_22,
  sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,sv2v_dc_27,sv2v_dc_28,sv2v_dc_29,
  sv2v_dc_30,sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,sv2v_dc_34,sv2v_dc_35,sv2v_dc_36,sv2v_dc_37,
  sv2v_dc_38,sv2v_dc_39,sv2v_dc_40,sv2v_dc_41,sv2v_dc_42,sv2v_dc_43,sv2v_dc_44,
  sv2v_dc_45,sv2v_dc_46,sv2v_dc_47,sv2v_dc_48,sv2v_dc_49,sv2v_dc_50,sv2v_dc_51,
  sv2v_dc_52,sv2v_dc_53,sv2v_dc_54,sv2v_dc_55,sv2v_dc_56,sv2v_dc_57,sv2v_dc_58,sv2v_dc_59,
  sv2v_dc_60,sv2v_dc_61,sv2v_dc_62,sv2v_dc_63,sv2v_dc_64,sv2v_dc_65,sv2v_dc_66,
  sv2v_dc_67,sv2v_dc_68,sv2v_dc_69,sv2v_dc_70,sv2v_dc_71,sv2v_dc_72,sv2v_dc_73,
  sv2v_dc_74,sv2v_dc_75,sv2v_dc_76,sv2v_dc_77,sv2v_dc_78,sv2v_dc_79,sv2v_dc_80,
  sv2v_dc_81,sv2v_dc_82,sv2v_dc_83,sv2v_dc_84,sv2v_dc_85,sv2v_dc_86,sv2v_dc_87,sv2v_dc_88,
  sv2v_dc_89,sv2v_dc_90,sv2v_dc_91,sv2v_dc_92,sv2v_dc_93,sv2v_dc_94,sv2v_dc_95,
  sv2v_dc_96,sv2v_dc_97,sv2v_dc_98,sv2v_dc_99,sv2v_dc_100,sv2v_dc_101,sv2v_dc_102,
  sv2v_dc_103,sv2v_dc_104,sv2v_dc_105,sv2v_dc_106,sv2v_dc_107,sv2v_dc_108,sv2v_dc_109,
  sv2v_dc_110,sv2v_dc_111,sv2v_dc_112,sv2v_dc_113,sv2v_dc_114,sv2v_dc_115,
  sv2v_dc_116,sv2v_dc_117,sv2v_dc_118,sv2v_dc_119,sv2v_dc_120,sv2v_dc_121,sv2v_dc_122,
  sv2v_dc_123,sv2v_dc_124,sv2v_dc_125,sv2v_dc_126,sv2v_dc_127;
  assign { o, sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36, sv2v_dc_37, sv2v_dc_38, sv2v_dc_39, sv2v_dc_40, sv2v_dc_41, sv2v_dc_42, sv2v_dc_43, sv2v_dc_44, sv2v_dc_45, sv2v_dc_46, sv2v_dc_47, sv2v_dc_48, sv2v_dc_49, sv2v_dc_50, sv2v_dc_51, sv2v_dc_52, sv2v_dc_53, sv2v_dc_54, sv2v_dc_55, sv2v_dc_56, sv2v_dc_57, sv2v_dc_58, sv2v_dc_59, sv2v_dc_60, sv2v_dc_61, sv2v_dc_62, sv2v_dc_63, sv2v_dc_64, sv2v_dc_65, sv2v_dc_66, sv2v_dc_67, sv2v_dc_68, sv2v_dc_69, sv2v_dc_70, sv2v_dc_71, sv2v_dc_72, sv2v_dc_73, sv2v_dc_74, sv2v_dc_75, sv2v_dc_76, sv2v_dc_77, sv2v_dc_78, sv2v_dc_79, sv2v_dc_80, sv2v_dc_81, sv2v_dc_82, sv2v_dc_83, sv2v_dc_84, sv2v_dc_85, sv2v_dc_86, sv2v_dc_87, sv2v_dc_88, sv2v_dc_89, sv2v_dc_90, sv2v_dc_91, sv2v_dc_92, sv2v_dc_93, sv2v_dc_94, sv2v_dc_95, sv2v_dc_96, sv2v_dc_97, sv2v_dc_98, sv2v_dc_99, sv2v_dc_100, sv2v_dc_101, sv2v_dc_102, sv2v_dc_103, sv2v_dc_104, sv2v_dc_105, sv2v_dc_106, sv2v_dc_107, sv2v_dc_108, sv2v_dc_109, sv2v_dc_110, sv2v_dc_111, sv2v_dc_112, sv2v_dc_113, sv2v_dc_114, sv2v_dc_115, sv2v_dc_116, sv2v_dc_117, sv2v_dc_118, sv2v_dc_119, sv2v_dc_120, sv2v_dc_121, sv2v_dc_122, sv2v_dc_123, sv2v_dc_124, sv2v_dc_125, sv2v_dc_126, sv2v_dc_127 } = { data_i, data_i[127:1] } << rot_i;

endmodule



module bsg_rotate_right_00000200
(
  data_i,
  rot_i,
  o
);

  input [511:0] data_i;
  input [8:0] rot_i;
  output [511:0] o;
  wire [511:0] o;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,
  sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,
  sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,sv2v_dc_21,sv2v_dc_22,
  sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,sv2v_dc_27,sv2v_dc_28,sv2v_dc_29,
  sv2v_dc_30,sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,sv2v_dc_34,sv2v_dc_35,sv2v_dc_36,sv2v_dc_37,
  sv2v_dc_38,sv2v_dc_39,sv2v_dc_40,sv2v_dc_41,sv2v_dc_42,sv2v_dc_43,sv2v_dc_44,
  sv2v_dc_45,sv2v_dc_46,sv2v_dc_47,sv2v_dc_48,sv2v_dc_49,sv2v_dc_50,sv2v_dc_51,
  sv2v_dc_52,sv2v_dc_53,sv2v_dc_54,sv2v_dc_55,sv2v_dc_56,sv2v_dc_57,sv2v_dc_58,sv2v_dc_59,
  sv2v_dc_60,sv2v_dc_61,sv2v_dc_62,sv2v_dc_63,sv2v_dc_64,sv2v_dc_65,sv2v_dc_66,
  sv2v_dc_67,sv2v_dc_68,sv2v_dc_69,sv2v_dc_70,sv2v_dc_71,sv2v_dc_72,sv2v_dc_73,
  sv2v_dc_74,sv2v_dc_75,sv2v_dc_76,sv2v_dc_77,sv2v_dc_78,sv2v_dc_79,sv2v_dc_80,
  sv2v_dc_81,sv2v_dc_82,sv2v_dc_83,sv2v_dc_84,sv2v_dc_85,sv2v_dc_86,sv2v_dc_87,sv2v_dc_88,
  sv2v_dc_89,sv2v_dc_90,sv2v_dc_91,sv2v_dc_92,sv2v_dc_93,sv2v_dc_94,sv2v_dc_95,
  sv2v_dc_96,sv2v_dc_97,sv2v_dc_98,sv2v_dc_99,sv2v_dc_100,sv2v_dc_101,sv2v_dc_102,
  sv2v_dc_103,sv2v_dc_104,sv2v_dc_105,sv2v_dc_106,sv2v_dc_107,sv2v_dc_108,sv2v_dc_109,
  sv2v_dc_110,sv2v_dc_111,sv2v_dc_112,sv2v_dc_113,sv2v_dc_114,sv2v_dc_115,
  sv2v_dc_116,sv2v_dc_117,sv2v_dc_118,sv2v_dc_119,sv2v_dc_120,sv2v_dc_121,sv2v_dc_122,
  sv2v_dc_123,sv2v_dc_124,sv2v_dc_125,sv2v_dc_126,sv2v_dc_127,sv2v_dc_128,sv2v_dc_129,
  sv2v_dc_130,sv2v_dc_131,sv2v_dc_132,sv2v_dc_133,sv2v_dc_134,sv2v_dc_135,
  sv2v_dc_136,sv2v_dc_137,sv2v_dc_138,sv2v_dc_139,sv2v_dc_140,sv2v_dc_141,sv2v_dc_142,
  sv2v_dc_143,sv2v_dc_144,sv2v_dc_145,sv2v_dc_146,sv2v_dc_147,sv2v_dc_148,sv2v_dc_149,
  sv2v_dc_150,sv2v_dc_151,sv2v_dc_152,sv2v_dc_153,sv2v_dc_154,sv2v_dc_155,
  sv2v_dc_156,sv2v_dc_157,sv2v_dc_158,sv2v_dc_159,sv2v_dc_160,sv2v_dc_161,sv2v_dc_162,
  sv2v_dc_163,sv2v_dc_164,sv2v_dc_165,sv2v_dc_166,sv2v_dc_167,sv2v_dc_168,sv2v_dc_169,
  sv2v_dc_170,sv2v_dc_171,sv2v_dc_172,sv2v_dc_173,sv2v_dc_174,sv2v_dc_175,
  sv2v_dc_176,sv2v_dc_177,sv2v_dc_178,sv2v_dc_179,sv2v_dc_180,sv2v_dc_181,sv2v_dc_182,
  sv2v_dc_183,sv2v_dc_184,sv2v_dc_185,sv2v_dc_186,sv2v_dc_187,sv2v_dc_188,sv2v_dc_189,
  sv2v_dc_190,sv2v_dc_191,sv2v_dc_192,sv2v_dc_193,sv2v_dc_194,sv2v_dc_195,
  sv2v_dc_196,sv2v_dc_197,sv2v_dc_198,sv2v_dc_199,sv2v_dc_200,sv2v_dc_201,sv2v_dc_202,
  sv2v_dc_203,sv2v_dc_204,sv2v_dc_205,sv2v_dc_206,sv2v_dc_207,sv2v_dc_208,sv2v_dc_209,
  sv2v_dc_210,sv2v_dc_211,sv2v_dc_212,sv2v_dc_213,sv2v_dc_214,sv2v_dc_215,
  sv2v_dc_216,sv2v_dc_217,sv2v_dc_218,sv2v_dc_219,sv2v_dc_220,sv2v_dc_221,sv2v_dc_222,
  sv2v_dc_223,sv2v_dc_224,sv2v_dc_225,sv2v_dc_226,sv2v_dc_227,sv2v_dc_228,sv2v_dc_229,
  sv2v_dc_230,sv2v_dc_231,sv2v_dc_232,sv2v_dc_233,sv2v_dc_234,sv2v_dc_235,
  sv2v_dc_236,sv2v_dc_237,sv2v_dc_238,sv2v_dc_239,sv2v_dc_240,sv2v_dc_241,sv2v_dc_242,
  sv2v_dc_243,sv2v_dc_244,sv2v_dc_245,sv2v_dc_246,sv2v_dc_247,sv2v_dc_248,sv2v_dc_249,
  sv2v_dc_250,sv2v_dc_251,sv2v_dc_252,sv2v_dc_253,sv2v_dc_254,sv2v_dc_255,
  sv2v_dc_256,sv2v_dc_257,sv2v_dc_258,sv2v_dc_259,sv2v_dc_260,sv2v_dc_261,sv2v_dc_262,
  sv2v_dc_263,sv2v_dc_264,sv2v_dc_265,sv2v_dc_266,sv2v_dc_267,sv2v_dc_268,sv2v_dc_269,
  sv2v_dc_270,sv2v_dc_271,sv2v_dc_272,sv2v_dc_273,sv2v_dc_274,sv2v_dc_275,
  sv2v_dc_276,sv2v_dc_277,sv2v_dc_278,sv2v_dc_279,sv2v_dc_280,sv2v_dc_281,sv2v_dc_282,
  sv2v_dc_283,sv2v_dc_284,sv2v_dc_285,sv2v_dc_286,sv2v_dc_287,sv2v_dc_288,sv2v_dc_289,
  sv2v_dc_290,sv2v_dc_291,sv2v_dc_292,sv2v_dc_293,sv2v_dc_294,sv2v_dc_295,
  sv2v_dc_296,sv2v_dc_297,sv2v_dc_298,sv2v_dc_299,sv2v_dc_300,sv2v_dc_301,sv2v_dc_302,
  sv2v_dc_303,sv2v_dc_304,sv2v_dc_305,sv2v_dc_306,sv2v_dc_307,sv2v_dc_308,sv2v_dc_309,
  sv2v_dc_310,sv2v_dc_311,sv2v_dc_312,sv2v_dc_313,sv2v_dc_314,sv2v_dc_315,
  sv2v_dc_316,sv2v_dc_317,sv2v_dc_318,sv2v_dc_319,sv2v_dc_320,sv2v_dc_321,sv2v_dc_322,
  sv2v_dc_323,sv2v_dc_324,sv2v_dc_325,sv2v_dc_326,sv2v_dc_327,sv2v_dc_328,sv2v_dc_329,
  sv2v_dc_330,sv2v_dc_331,sv2v_dc_332,sv2v_dc_333,sv2v_dc_334,sv2v_dc_335,
  sv2v_dc_336,sv2v_dc_337,sv2v_dc_338,sv2v_dc_339,sv2v_dc_340,sv2v_dc_341,sv2v_dc_342,
  sv2v_dc_343,sv2v_dc_344,sv2v_dc_345,sv2v_dc_346,sv2v_dc_347,sv2v_dc_348,sv2v_dc_349,
  sv2v_dc_350,sv2v_dc_351,sv2v_dc_352,sv2v_dc_353,sv2v_dc_354,sv2v_dc_355,
  sv2v_dc_356,sv2v_dc_357,sv2v_dc_358,sv2v_dc_359,sv2v_dc_360,sv2v_dc_361,sv2v_dc_362,
  sv2v_dc_363,sv2v_dc_364,sv2v_dc_365,sv2v_dc_366,sv2v_dc_367,sv2v_dc_368,sv2v_dc_369,
  sv2v_dc_370,sv2v_dc_371,sv2v_dc_372,sv2v_dc_373,sv2v_dc_374,sv2v_dc_375,
  sv2v_dc_376,sv2v_dc_377,sv2v_dc_378,sv2v_dc_379,sv2v_dc_380,sv2v_dc_381,sv2v_dc_382,
  sv2v_dc_383,sv2v_dc_384,sv2v_dc_385,sv2v_dc_386,sv2v_dc_387,sv2v_dc_388,sv2v_dc_389,
  sv2v_dc_390,sv2v_dc_391,sv2v_dc_392,sv2v_dc_393,sv2v_dc_394,sv2v_dc_395,
  sv2v_dc_396,sv2v_dc_397,sv2v_dc_398,sv2v_dc_399,sv2v_dc_400,sv2v_dc_401,sv2v_dc_402,
  sv2v_dc_403,sv2v_dc_404,sv2v_dc_405,sv2v_dc_406,sv2v_dc_407,sv2v_dc_408,sv2v_dc_409,
  sv2v_dc_410,sv2v_dc_411,sv2v_dc_412,sv2v_dc_413,sv2v_dc_414,sv2v_dc_415,
  sv2v_dc_416,sv2v_dc_417,sv2v_dc_418,sv2v_dc_419,sv2v_dc_420,sv2v_dc_421,sv2v_dc_422,
  sv2v_dc_423,sv2v_dc_424,sv2v_dc_425,sv2v_dc_426,sv2v_dc_427,sv2v_dc_428,sv2v_dc_429,
  sv2v_dc_430,sv2v_dc_431,sv2v_dc_432,sv2v_dc_433,sv2v_dc_434,sv2v_dc_435,
  sv2v_dc_436,sv2v_dc_437,sv2v_dc_438,sv2v_dc_439,sv2v_dc_440,sv2v_dc_441,sv2v_dc_442,
  sv2v_dc_443,sv2v_dc_444,sv2v_dc_445,sv2v_dc_446,sv2v_dc_447,sv2v_dc_448,sv2v_dc_449,
  sv2v_dc_450,sv2v_dc_451,sv2v_dc_452,sv2v_dc_453,sv2v_dc_454,sv2v_dc_455,
  sv2v_dc_456,sv2v_dc_457,sv2v_dc_458,sv2v_dc_459,sv2v_dc_460,sv2v_dc_461,sv2v_dc_462,
  sv2v_dc_463,sv2v_dc_464,sv2v_dc_465,sv2v_dc_466,sv2v_dc_467,sv2v_dc_468,sv2v_dc_469,
  sv2v_dc_470,sv2v_dc_471,sv2v_dc_472,sv2v_dc_473,sv2v_dc_474,sv2v_dc_475,
  sv2v_dc_476,sv2v_dc_477,sv2v_dc_478,sv2v_dc_479,sv2v_dc_480,sv2v_dc_481,sv2v_dc_482,
  sv2v_dc_483,sv2v_dc_484,sv2v_dc_485,sv2v_dc_486,sv2v_dc_487,sv2v_dc_488,sv2v_dc_489,
  sv2v_dc_490,sv2v_dc_491,sv2v_dc_492,sv2v_dc_493,sv2v_dc_494,sv2v_dc_495,
  sv2v_dc_496,sv2v_dc_497,sv2v_dc_498,sv2v_dc_499,sv2v_dc_500,sv2v_dc_501,sv2v_dc_502,
  sv2v_dc_503,sv2v_dc_504,sv2v_dc_505,sv2v_dc_506,sv2v_dc_507,sv2v_dc_508,sv2v_dc_509,
  sv2v_dc_510,sv2v_dc_511;
  assign { sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36, sv2v_dc_37, sv2v_dc_38, sv2v_dc_39, sv2v_dc_40, sv2v_dc_41, sv2v_dc_42, sv2v_dc_43, sv2v_dc_44, sv2v_dc_45, sv2v_dc_46, sv2v_dc_47, sv2v_dc_48, sv2v_dc_49, sv2v_dc_50, sv2v_dc_51, sv2v_dc_52, sv2v_dc_53, sv2v_dc_54, sv2v_dc_55, sv2v_dc_56, sv2v_dc_57, sv2v_dc_58, sv2v_dc_59, sv2v_dc_60, sv2v_dc_61, sv2v_dc_62, sv2v_dc_63, sv2v_dc_64, sv2v_dc_65, sv2v_dc_66, sv2v_dc_67, sv2v_dc_68, sv2v_dc_69, sv2v_dc_70, sv2v_dc_71, sv2v_dc_72, sv2v_dc_73, sv2v_dc_74, sv2v_dc_75, sv2v_dc_76, sv2v_dc_77, sv2v_dc_78, sv2v_dc_79, sv2v_dc_80, sv2v_dc_81, sv2v_dc_82, sv2v_dc_83, sv2v_dc_84, sv2v_dc_85, sv2v_dc_86, sv2v_dc_87, sv2v_dc_88, sv2v_dc_89, sv2v_dc_90, sv2v_dc_91, sv2v_dc_92, sv2v_dc_93, sv2v_dc_94, sv2v_dc_95, sv2v_dc_96, sv2v_dc_97, sv2v_dc_98, sv2v_dc_99, sv2v_dc_100, sv2v_dc_101, sv2v_dc_102, sv2v_dc_103, sv2v_dc_104, sv2v_dc_105, sv2v_dc_106, sv2v_dc_107, sv2v_dc_108, sv2v_dc_109, sv2v_dc_110, sv2v_dc_111, sv2v_dc_112, sv2v_dc_113, sv2v_dc_114, sv2v_dc_115, sv2v_dc_116, sv2v_dc_117, sv2v_dc_118, sv2v_dc_119, sv2v_dc_120, sv2v_dc_121, sv2v_dc_122, sv2v_dc_123, sv2v_dc_124, sv2v_dc_125, sv2v_dc_126, sv2v_dc_127, sv2v_dc_128, sv2v_dc_129, sv2v_dc_130, sv2v_dc_131, sv2v_dc_132, sv2v_dc_133, sv2v_dc_134, sv2v_dc_135, sv2v_dc_136, sv2v_dc_137, sv2v_dc_138, sv2v_dc_139, sv2v_dc_140, sv2v_dc_141, sv2v_dc_142, sv2v_dc_143, sv2v_dc_144, sv2v_dc_145, sv2v_dc_146, sv2v_dc_147, sv2v_dc_148, sv2v_dc_149, sv2v_dc_150, sv2v_dc_151, sv2v_dc_152, sv2v_dc_153, sv2v_dc_154, sv2v_dc_155, sv2v_dc_156, sv2v_dc_157, sv2v_dc_158, sv2v_dc_159, sv2v_dc_160, sv2v_dc_161, sv2v_dc_162, sv2v_dc_163, sv2v_dc_164, sv2v_dc_165, sv2v_dc_166, sv2v_dc_167, sv2v_dc_168, sv2v_dc_169, sv2v_dc_170, sv2v_dc_171, sv2v_dc_172, sv2v_dc_173, sv2v_dc_174, sv2v_dc_175, sv2v_dc_176, sv2v_dc_177, sv2v_dc_178, sv2v_dc_179, sv2v_dc_180, sv2v_dc_181, sv2v_dc_182, sv2v_dc_183, sv2v_dc_184, sv2v_dc_185, sv2v_dc_186, sv2v_dc_187, sv2v_dc_188, sv2v_dc_189, sv2v_dc_190, sv2v_dc_191, sv2v_dc_192, sv2v_dc_193, sv2v_dc_194, sv2v_dc_195, sv2v_dc_196, sv2v_dc_197, sv2v_dc_198, sv2v_dc_199, sv2v_dc_200, sv2v_dc_201, sv2v_dc_202, sv2v_dc_203, sv2v_dc_204, sv2v_dc_205, sv2v_dc_206, sv2v_dc_207, sv2v_dc_208, sv2v_dc_209, sv2v_dc_210, sv2v_dc_211, sv2v_dc_212, sv2v_dc_213, sv2v_dc_214, sv2v_dc_215, sv2v_dc_216, sv2v_dc_217, sv2v_dc_218, sv2v_dc_219, sv2v_dc_220, sv2v_dc_221, sv2v_dc_222, sv2v_dc_223, sv2v_dc_224, sv2v_dc_225, sv2v_dc_226, sv2v_dc_227, sv2v_dc_228, sv2v_dc_229, sv2v_dc_230, sv2v_dc_231, sv2v_dc_232, sv2v_dc_233, sv2v_dc_234, sv2v_dc_235, sv2v_dc_236, sv2v_dc_237, sv2v_dc_238, sv2v_dc_239, sv2v_dc_240, sv2v_dc_241, sv2v_dc_242, sv2v_dc_243, sv2v_dc_244, sv2v_dc_245, sv2v_dc_246, sv2v_dc_247, sv2v_dc_248, sv2v_dc_249, sv2v_dc_250, sv2v_dc_251, sv2v_dc_252, sv2v_dc_253, sv2v_dc_254, sv2v_dc_255, sv2v_dc_256, sv2v_dc_257, sv2v_dc_258, sv2v_dc_259, sv2v_dc_260, sv2v_dc_261, sv2v_dc_262, sv2v_dc_263, sv2v_dc_264, sv2v_dc_265, sv2v_dc_266, sv2v_dc_267, sv2v_dc_268, sv2v_dc_269, sv2v_dc_270, sv2v_dc_271, sv2v_dc_272, sv2v_dc_273, sv2v_dc_274, sv2v_dc_275, sv2v_dc_276, sv2v_dc_277, sv2v_dc_278, sv2v_dc_279, sv2v_dc_280, sv2v_dc_281, sv2v_dc_282, sv2v_dc_283, sv2v_dc_284, sv2v_dc_285, sv2v_dc_286, sv2v_dc_287, sv2v_dc_288, sv2v_dc_289, sv2v_dc_290, sv2v_dc_291, sv2v_dc_292, sv2v_dc_293, sv2v_dc_294, sv2v_dc_295, sv2v_dc_296, sv2v_dc_297, sv2v_dc_298, sv2v_dc_299, sv2v_dc_300, sv2v_dc_301, sv2v_dc_302, sv2v_dc_303, sv2v_dc_304, sv2v_dc_305, sv2v_dc_306, sv2v_dc_307, sv2v_dc_308, sv2v_dc_309, sv2v_dc_310, sv2v_dc_311, sv2v_dc_312, sv2v_dc_313, sv2v_dc_314, sv2v_dc_315, sv2v_dc_316, sv2v_dc_317, sv2v_dc_318, sv2v_dc_319, sv2v_dc_320, sv2v_dc_321, sv2v_dc_322, sv2v_dc_323, sv2v_dc_324, sv2v_dc_325, sv2v_dc_326, sv2v_dc_327, sv2v_dc_328, sv2v_dc_329, sv2v_dc_330, sv2v_dc_331, sv2v_dc_332, sv2v_dc_333, sv2v_dc_334, sv2v_dc_335, sv2v_dc_336, sv2v_dc_337, sv2v_dc_338, sv2v_dc_339, sv2v_dc_340, sv2v_dc_341, sv2v_dc_342, sv2v_dc_343, sv2v_dc_344, sv2v_dc_345, sv2v_dc_346, sv2v_dc_347, sv2v_dc_348, sv2v_dc_349, sv2v_dc_350, sv2v_dc_351, sv2v_dc_352, sv2v_dc_353, sv2v_dc_354, sv2v_dc_355, sv2v_dc_356, sv2v_dc_357, sv2v_dc_358, sv2v_dc_359, sv2v_dc_360, sv2v_dc_361, sv2v_dc_362, sv2v_dc_363, sv2v_dc_364, sv2v_dc_365, sv2v_dc_366, sv2v_dc_367, sv2v_dc_368, sv2v_dc_369, sv2v_dc_370, sv2v_dc_371, sv2v_dc_372, sv2v_dc_373, sv2v_dc_374, sv2v_dc_375, sv2v_dc_376, sv2v_dc_377, sv2v_dc_378, sv2v_dc_379, sv2v_dc_380, sv2v_dc_381, sv2v_dc_382, sv2v_dc_383, sv2v_dc_384, sv2v_dc_385, sv2v_dc_386, sv2v_dc_387, sv2v_dc_388, sv2v_dc_389, sv2v_dc_390, sv2v_dc_391, sv2v_dc_392, sv2v_dc_393, sv2v_dc_394, sv2v_dc_395, sv2v_dc_396, sv2v_dc_397, sv2v_dc_398, sv2v_dc_399, sv2v_dc_400, sv2v_dc_401, sv2v_dc_402, sv2v_dc_403, sv2v_dc_404, sv2v_dc_405, sv2v_dc_406, sv2v_dc_407, sv2v_dc_408, sv2v_dc_409, sv2v_dc_410, sv2v_dc_411, sv2v_dc_412, sv2v_dc_413, sv2v_dc_414, sv2v_dc_415, sv2v_dc_416, sv2v_dc_417, sv2v_dc_418, sv2v_dc_419, sv2v_dc_420, sv2v_dc_421, sv2v_dc_422, sv2v_dc_423, sv2v_dc_424, sv2v_dc_425, sv2v_dc_426, sv2v_dc_427, sv2v_dc_428, sv2v_dc_429, sv2v_dc_430, sv2v_dc_431, sv2v_dc_432, sv2v_dc_433, sv2v_dc_434, sv2v_dc_435, sv2v_dc_436, sv2v_dc_437, sv2v_dc_438, sv2v_dc_439, sv2v_dc_440, sv2v_dc_441, sv2v_dc_442, sv2v_dc_443, sv2v_dc_444, sv2v_dc_445, sv2v_dc_446, sv2v_dc_447, sv2v_dc_448, sv2v_dc_449, sv2v_dc_450, sv2v_dc_451, sv2v_dc_452, sv2v_dc_453, sv2v_dc_454, sv2v_dc_455, sv2v_dc_456, sv2v_dc_457, sv2v_dc_458, sv2v_dc_459, sv2v_dc_460, sv2v_dc_461, sv2v_dc_462, sv2v_dc_463, sv2v_dc_464, sv2v_dc_465, sv2v_dc_466, sv2v_dc_467, sv2v_dc_468, sv2v_dc_469, sv2v_dc_470, sv2v_dc_471, sv2v_dc_472, sv2v_dc_473, sv2v_dc_474, sv2v_dc_475, sv2v_dc_476, sv2v_dc_477, sv2v_dc_478, sv2v_dc_479, sv2v_dc_480, sv2v_dc_481, sv2v_dc_482, sv2v_dc_483, sv2v_dc_484, sv2v_dc_485, sv2v_dc_486, sv2v_dc_487, sv2v_dc_488, sv2v_dc_489, sv2v_dc_490, sv2v_dc_491, sv2v_dc_492, sv2v_dc_493, sv2v_dc_494, sv2v_dc_495, sv2v_dc_496, sv2v_dc_497, sv2v_dc_498, sv2v_dc_499, sv2v_dc_500, sv2v_dc_501, sv2v_dc_502, sv2v_dc_503, sv2v_dc_504, sv2v_dc_505, sv2v_dc_506, sv2v_dc_507, sv2v_dc_508, sv2v_dc_509, sv2v_dc_510, sv2v_dc_511, o } = { data_i[510:0], data_i } >> rot_i;

endmodule



module bsg_lru_pseudo_tree_decode_00000008
(
  way_id_i,
  data_o,
  mask_o
);

  input [2:0] way_id_i;
  output [6:0] data_o;
  output [6:0] mask_o;
  wire [6:0] data_o,mask_o;
  wire N0,N1,N2;
  assign mask_o[0] = 1'b1;
  assign data_o[0] = 1'b1 & N0;
  assign N0 = ~way_id_i[2];
  assign mask_o[1] = 1'b1 & N0;
  assign data_o[1] = mask_o[1] & N1;
  assign N1 = ~way_id_i[1];
  assign mask_o[2] = 1'b1 & way_id_i[2];
  assign data_o[2] = mask_o[2] & N1;
  assign mask_o[3] = mask_o[1] & N1;
  assign data_o[3] = mask_o[3] & N2;
  assign N2 = ~way_id_i[0];
  assign mask_o[4] = mask_o[1] & way_id_i[1];
  assign data_o[4] = mask_o[4] & N2;
  assign mask_o[5] = mask_o[2] & N1;
  assign data_o[5] = mask_o[5] & N2;
  assign mask_o[6] = mask_o[2] & way_id_i[1];
  assign data_o[6] = mask_o[6] & N2;

endmodule



module bsg_decode_with_v_00000008
(
  i,
  v_i,
  o
);

  input [2:0] i;
  output [7:0] o;
  input v_i;
  wire [7:0] o,lo;

  bsg_decode_00000008
  bd
  (
    .i(i),
    .o(lo)
  );

  assign o[7] = v_i & lo[7];
  assign o[6] = v_i & lo[6];
  assign o[5] = v_i & lo[5];
  assign o[4] = v_i & lo[4];
  assign o[3] = v_i & lo[3];
  assign o[2] = v_i & lo[2];
  assign o[1] = v_i & lo[1];
  assign o[0] = v_i & lo[0];

endmodule



module bsg_dff_reset_set_clear_width_p1_clear_over_set_p1
(
  clk_i,
  reset_i,
  set_i,
  clear_i,
  data_o
);

  input [0:0] set_i;
  input [0:0] clear_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  wire [0:0] data_o;
  wire N0,N1,N2;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N0 = N1 & N2;
  assign N1 = data_o[0] | set_i[0];
  assign N2 = ~clear_i[0];

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_0_sv2v_reg <= N0;
    end 
  end


endmodule



module bsg_dff_en_0000001a
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [25:0] data_i;
  output [25:0] data_o;
  input clk_i;
  input en_i;
  wire [25:0] data_o;
  reg data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,
  data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,
  data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_counter_clear_up_max_val_p15_init_val_p0_disable_overflow_warning_p1
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [3:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire [3:0] count_o;
  wire N0,N1,N4,N5,N6,N8,N9,N10,N11,N12,N13,N14,N15,N16,N2,N3,N7,N30,N17;
  reg count_o_3_sv2v_reg,count_o_2_sv2v_reg,count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[3] = count_o_3_sv2v_reg;
  assign count_o[2] = count_o_2_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign N17 = reset_i | clear_i;
  assign { N9, N8, N6, N5 } = count_o + 1'b1;
  assign N10 = (N0)? 1'b1 : 
               (N7)? 1'b1 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = clear_i;
  assign N12 = (N1)? 1'b1 : 
               (N30)? 1'b0 : 1'b0;
  assign N1 = up_i;
  assign N11 = (N0)? up_i : 
               (N7)? N5 : 1'b0;
  assign N4 = N16;
  assign N13 = ~reset_i;
  assign N14 = ~clear_i;
  assign N15 = N13 & N14;
  assign N16 = up_i & N15;
  assign N2 = up_i | clear_i;
  assign N3 = ~N2;
  assign N7 = up_i & N14;
  assign N30 = ~up_i;

  always @(posedge clk_i) begin
    if(N17) begin
      count_o_3_sv2v_reg <= 1'b0;
      count_o_2_sv2v_reg <= 1'b0;
      count_o_1_sv2v_reg <= 1'b0;
    end else if(N12) begin
      count_o_3_sv2v_reg <= N9;
      count_o_2_sv2v_reg <= N8;
      count_o_1_sv2v_reg <= N6;
    end 
    if(reset_i) begin
      count_o_0_sv2v_reg <= 1'b0;
    end else if(N10) begin
      count_o_0_sv2v_reg <= N11;
    end 
  end


endmodule



module bsg_dff_en_0000008a
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [137:0] data_i;
  output [137:0] data_o;
  input clk_i;
  input en_i;
  wire [137:0] data_o;
  reg data_o_137_sv2v_reg,data_o_136_sv2v_reg,data_o_135_sv2v_reg,data_o_134_sv2v_reg,
  data_o_133_sv2v_reg,data_o_132_sv2v_reg,data_o_131_sv2v_reg,data_o_130_sv2v_reg,
  data_o_129_sv2v_reg,data_o_128_sv2v_reg,data_o_127_sv2v_reg,data_o_126_sv2v_reg,
  data_o_125_sv2v_reg,data_o_124_sv2v_reg,data_o_123_sv2v_reg,data_o_122_sv2v_reg,
  data_o_121_sv2v_reg,data_o_120_sv2v_reg,data_o_119_sv2v_reg,data_o_118_sv2v_reg,
  data_o_117_sv2v_reg,data_o_116_sv2v_reg,data_o_115_sv2v_reg,data_o_114_sv2v_reg,
  data_o_113_sv2v_reg,data_o_112_sv2v_reg,data_o_111_sv2v_reg,data_o_110_sv2v_reg,
  data_o_109_sv2v_reg,data_o_108_sv2v_reg,data_o_107_sv2v_reg,data_o_106_sv2v_reg,
  data_o_105_sv2v_reg,data_o_104_sv2v_reg,data_o_103_sv2v_reg,data_o_102_sv2v_reg,
  data_o_101_sv2v_reg,data_o_100_sv2v_reg,data_o_99_sv2v_reg,data_o_98_sv2v_reg,
  data_o_97_sv2v_reg,data_o_96_sv2v_reg,data_o_95_sv2v_reg,data_o_94_sv2v_reg,
  data_o_93_sv2v_reg,data_o_92_sv2v_reg,data_o_91_sv2v_reg,data_o_90_sv2v_reg,
  data_o_89_sv2v_reg,data_o_88_sv2v_reg,data_o_87_sv2v_reg,data_o_86_sv2v_reg,
  data_o_85_sv2v_reg,data_o_84_sv2v_reg,data_o_83_sv2v_reg,data_o_82_sv2v_reg,
  data_o_81_sv2v_reg,data_o_80_sv2v_reg,data_o_79_sv2v_reg,data_o_78_sv2v_reg,data_o_77_sv2v_reg,
  data_o_76_sv2v_reg,data_o_75_sv2v_reg,data_o_74_sv2v_reg,data_o_73_sv2v_reg,
  data_o_72_sv2v_reg,data_o_71_sv2v_reg,data_o_70_sv2v_reg,data_o_69_sv2v_reg,
  data_o_68_sv2v_reg,data_o_67_sv2v_reg,data_o_66_sv2v_reg,data_o_65_sv2v_reg,
  data_o_64_sv2v_reg,data_o_63_sv2v_reg,data_o_62_sv2v_reg,data_o_61_sv2v_reg,data_o_60_sv2v_reg,
  data_o_59_sv2v_reg,data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,
  data_o_55_sv2v_reg,data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,
  data_o_51_sv2v_reg,data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,
  data_o_47_sv2v_reg,data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,
  data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,
  data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,
  data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,
  data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,
  data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,
  data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,
  data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[137] = data_o_137_sv2v_reg;
  assign data_o[136] = data_o_136_sv2v_reg;
  assign data_o[135] = data_o_135_sv2v_reg;
  assign data_o[134] = data_o_134_sv2v_reg;
  assign data_o[133] = data_o_133_sv2v_reg;
  assign data_o[132] = data_o_132_sv2v_reg;
  assign data_o[131] = data_o_131_sv2v_reg;
  assign data_o[130] = data_o_130_sv2v_reg;
  assign data_o[129] = data_o_129_sv2v_reg;
  assign data_o[128] = data_o_128_sv2v_reg;
  assign data_o[127] = data_o_127_sv2v_reg;
  assign data_o[126] = data_o_126_sv2v_reg;
  assign data_o[125] = data_o_125_sv2v_reg;
  assign data_o[124] = data_o_124_sv2v_reg;
  assign data_o[123] = data_o_123_sv2v_reg;
  assign data_o[122] = data_o_122_sv2v_reg;
  assign data_o[121] = data_o_121_sv2v_reg;
  assign data_o[120] = data_o_120_sv2v_reg;
  assign data_o[119] = data_o_119_sv2v_reg;
  assign data_o[118] = data_o_118_sv2v_reg;
  assign data_o[117] = data_o_117_sv2v_reg;
  assign data_o[116] = data_o_116_sv2v_reg;
  assign data_o[115] = data_o_115_sv2v_reg;
  assign data_o[114] = data_o_114_sv2v_reg;
  assign data_o[113] = data_o_113_sv2v_reg;
  assign data_o[112] = data_o_112_sv2v_reg;
  assign data_o[111] = data_o_111_sv2v_reg;
  assign data_o[110] = data_o_110_sv2v_reg;
  assign data_o[109] = data_o_109_sv2v_reg;
  assign data_o[108] = data_o_108_sv2v_reg;
  assign data_o[107] = data_o_107_sv2v_reg;
  assign data_o[106] = data_o_106_sv2v_reg;
  assign data_o[105] = data_o_105_sv2v_reg;
  assign data_o[104] = data_o_104_sv2v_reg;
  assign data_o[103] = data_o_103_sv2v_reg;
  assign data_o[102] = data_o_102_sv2v_reg;
  assign data_o[101] = data_o_101_sv2v_reg;
  assign data_o[100] = data_o_100_sv2v_reg;
  assign data_o[99] = data_o_99_sv2v_reg;
  assign data_o[98] = data_o_98_sv2v_reg;
  assign data_o[97] = data_o_97_sv2v_reg;
  assign data_o[96] = data_o_96_sv2v_reg;
  assign data_o[95] = data_o_95_sv2v_reg;
  assign data_o[94] = data_o_94_sv2v_reg;
  assign data_o[93] = data_o_93_sv2v_reg;
  assign data_o[92] = data_o_92_sv2v_reg;
  assign data_o[91] = data_o_91_sv2v_reg;
  assign data_o[90] = data_o_90_sv2v_reg;
  assign data_o[89] = data_o_89_sv2v_reg;
  assign data_o[88] = data_o_88_sv2v_reg;
  assign data_o[87] = data_o_87_sv2v_reg;
  assign data_o[86] = data_o_86_sv2v_reg;
  assign data_o[85] = data_o_85_sv2v_reg;
  assign data_o[84] = data_o_84_sv2v_reg;
  assign data_o[83] = data_o_83_sv2v_reg;
  assign data_o[82] = data_o_82_sv2v_reg;
  assign data_o[81] = data_o_81_sv2v_reg;
  assign data_o[80] = data_o_80_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_137_sv2v_reg <= data_i[137];
      data_o_136_sv2v_reg <= data_i[136];
      data_o_135_sv2v_reg <= data_i[135];
      data_o_134_sv2v_reg <= data_i[134];
      data_o_133_sv2v_reg <= data_i[133];
      data_o_132_sv2v_reg <= data_i[132];
      data_o_131_sv2v_reg <= data_i[131];
      data_o_130_sv2v_reg <= data_i[130];
      data_o_129_sv2v_reg <= data_i[129];
      data_o_128_sv2v_reg <= data_i[128];
      data_o_127_sv2v_reg <= data_i[127];
      data_o_126_sv2v_reg <= data_i[126];
      data_o_125_sv2v_reg <= data_i[125];
      data_o_124_sv2v_reg <= data_i[124];
      data_o_123_sv2v_reg <= data_i[123];
      data_o_122_sv2v_reg <= data_i[122];
      data_o_121_sv2v_reg <= data_i[121];
      data_o_120_sv2v_reg <= data_i[120];
      data_o_119_sv2v_reg <= data_i[119];
      data_o_118_sv2v_reg <= data_i[118];
      data_o_117_sv2v_reg <= data_i[117];
      data_o_116_sv2v_reg <= data_i[116];
      data_o_115_sv2v_reg <= data_i[115];
      data_o_114_sv2v_reg <= data_i[114];
      data_o_113_sv2v_reg <= data_i[113];
      data_o_112_sv2v_reg <= data_i[112];
      data_o_111_sv2v_reg <= data_i[111];
      data_o_110_sv2v_reg <= data_i[110];
      data_o_109_sv2v_reg <= data_i[109];
      data_o_108_sv2v_reg <= data_i[108];
      data_o_107_sv2v_reg <= data_i[107];
      data_o_106_sv2v_reg <= data_i[106];
      data_o_105_sv2v_reg <= data_i[105];
      data_o_104_sv2v_reg <= data_i[104];
      data_o_103_sv2v_reg <= data_i[103];
      data_o_102_sv2v_reg <= data_i[102];
      data_o_101_sv2v_reg <= data_i[101];
      data_o_100_sv2v_reg <= data_i[100];
      data_o_99_sv2v_reg <= data_i[99];
      data_o_98_sv2v_reg <= data_i[98];
      data_o_97_sv2v_reg <= data_i[97];
      data_o_96_sv2v_reg <= data_i[96];
      data_o_95_sv2v_reg <= data_i[95];
      data_o_94_sv2v_reg <= data_i[94];
      data_o_93_sv2v_reg <= data_i[93];
      data_o_92_sv2v_reg <= data_i[92];
      data_o_91_sv2v_reg <= data_i[91];
      data_o_90_sv2v_reg <= data_i[90];
      data_o_89_sv2v_reg <= data_i[89];
      data_o_88_sv2v_reg <= data_i[88];
      data_o_87_sv2v_reg <= data_i[87];
      data_o_86_sv2v_reg <= data_i[86];
      data_o_85_sv2v_reg <= data_i[85];
      data_o_84_sv2v_reg <= data_i[84];
      data_o_83_sv2v_reg <= data_i[83];
      data_o_82_sv2v_reg <= data_i[82];
      data_o_81_sv2v_reg <= data_i[81];
      data_o_80_sv2v_reg <= data_i[80];
      data_o_79_sv2v_reg <= data_i[79];
      data_o_78_sv2v_reg <= data_i[78];
      data_o_77_sv2v_reg <= data_i[77];
      data_o_76_sv2v_reg <= data_i[76];
      data_o_75_sv2v_reg <= data_i[75];
      data_o_74_sv2v_reg <= data_i[74];
      data_o_73_sv2v_reg <= data_i[73];
      data_o_72_sv2v_reg <= data_i[72];
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_en_00000010
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [15:0] data_i;
  output [15:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [15:0] data_o;
  wire N0,N1,N2;
  reg data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,
  data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,
  data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bp_be_dcache
(
  clk_i,
  reset_i,
  cfg_bus_i,
  busy_o,
  ordered_o,
  dcache_pkt_i,
  v_i,
  ptag_i,
  ptag_v_i,
  ptag_uncached_i,
  ptag_dram_i,
  st_data_i,
  flush_i,
  v_o,
  data_o,
  rd_addr_o,
  tag_o,
  unsigned_o,
  int_o,
  float_o,
  ptw_o,
  ret_o,
  late_o,
  cache_req_o,
  cache_req_v_o,
  cache_req_yumi_i,
  cache_req_lock_i,
  cache_req_metadata_o,
  cache_req_metadata_v_o,
  cache_req_id_i,
  cache_req_critical_i,
  cache_req_last_i,
  cache_req_credits_full_i,
  cache_req_credits_empty_i,
  data_mem_pkt_v_i,
  data_mem_pkt_i,
  data_mem_pkt_yumi_o,
  data_mem_o,
  tag_mem_pkt_v_i,
  tag_mem_pkt_i,
  tag_mem_pkt_yumi_o,
  tag_mem_o,
  stat_mem_pkt_v_i,
  stat_mem_pkt_i,
  stat_mem_pkt_yumi_o,
  stat_mem_o
);

  input [60:0] cfg_bus_i;
  input [22:0] dcache_pkt_i;
  input [27:0] ptag_i;
  input [63:0] st_data_i;
  output [63:0] data_o;
  output [4:0] rd_addr_o;
  output [1:0] tag_o;
  output [116:0] cache_req_o;
  output [3:0] cache_req_metadata_o;
  input [0:0] cache_req_id_i;
  input [142:0] data_mem_pkt_i;
  output [511:0] data_mem_o;
  input [34:0] tag_mem_pkt_i;
  output [22:0] tag_mem_o;
  input [10:0] stat_mem_pkt_i;
  output [14:0] stat_mem_o;
  input clk_i;
  input reset_i;
  input v_i;
  input ptag_v_i;
  input ptag_uncached_i;
  input ptag_dram_i;
  input flush_i;
  input cache_req_yumi_i;
  input cache_req_lock_i;
  input cache_req_critical_i;
  input cache_req_last_i;
  input cache_req_credits_full_i;
  input cache_req_credits_empty_i;
  input data_mem_pkt_v_i;
  input tag_mem_pkt_v_i;
  input stat_mem_pkt_v_i;
  output busy_o;
  output ordered_o;
  output v_o;
  output unsigned_o;
  output int_o;
  output float_o;
  output ptw_o;
  output ret_o;
  output late_o;
  output cache_req_v_o;
  output cache_req_metadata_v_o;
  output data_mem_pkt_yumi_o;
  output tag_mem_pkt_yumi_o;
  output stat_mem_pkt_yumi_o;
  wire [63:0] data_o,data_mem_mask_li,st_data_tv_n,snoop_st_data,ld_data_way_picked,
  ld_data_dword_raw,ld_data_dword_merged,final_data_tv,atomic_reg_data,atomic_mem_data,
  atomic_alu_result,atomic_result,\wbuf_in_3_.slice_data ;
  wire [4:0] rd_addr_o;
  wire [1:0] tag_o,state_r,\wbuf_in_2_.addr_dec ,state_n;
  wire [116:0] cache_req_o;
  wire [3:0] cache_req_metadata_o,\wbuf_in_1_.addr_dec ,\l1_lrsc.lrsc_lock_cnt ;
  wire [511:0] data_mem_o,data_mem_data_li,data_mem_data_lo,ld_data_tv_n,ld_data_tv_r;
  wire [22:0] tag_mem_o;
  wire [14:0] stat_mem_o,stat_mem_data_li,stat_mem_mask_li;
  wire busy_o,ordered_o,v_o,unsigned_o,int_o,float_o,ptw_o,ret_o,late_o,cache_req_v_o,
  cache_req_metadata_v_o,data_mem_pkt_yumi_o,tag_mem_pkt_yumi_o,
  stat_mem_pkt_yumi_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,blocking_hazard,nonblocking_hazard,fill_hazard,
  flush_tv,data_mem_write_hazard,flush_tl,critical_recv,complete_recv,tag_mem_v_li,
  tag_mem_w_li,safe_tl_we,tl_we,v_tl_r,N89,\tag_comp_tl_0_.tag_match_tl ,N90,N91,N92,
  N93,N94,N95,N96,N97,N98,N99,\tag_comp_tl_1_.tag_match_tl ,N100,N101,N102,N103,
  N104,N105,N106,N107,N108,N109,\tag_comp_tl_2_.tag_match_tl ,N110,N111,N112,N113,
  N114,N115,N116,N117,N118,N119,\tag_comp_tl_3_.tag_match_tl ,N120,N121,N122,N123,
  N124,N125,N126,N127,N128,N129,\tag_comp_tl_4_.tag_match_tl ,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,\tag_comp_tl_5_.tag_match_tl ,N140,N141,N142,N143,
  N144,N145,N146,N147,N148,N149,\tag_comp_tl_6_.tag_match_tl ,N150,N151,N152,N153,
  N154,N155,N156,N157,N158,N159,\tag_comp_tl_7_.tag_match_tl ,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,uncached_tl,safe_tv_we,tv_we,_2_net_,v_tv_r,uncached_tv_n,
  snoop_paddr_5,snoop_paddr_4,snoop_paddr_3,snoop_paddr_2,snoop_paddr_1,
  snoop_paddr_0,snoop_uncached,decode_tv_r_load_op_,decode_tv_r_store_op_,
  decode_tv_r_signed_op_,decode_tv_r_cache_op_,decode_tv_r_block_op_,decode_tv_r_double_op_,
  decode_tv_r_word_op_,decode_tv_r_half_op_,decode_tv_r_byte_op_,decode_tv_r_uncached_op_,
  decode_tv_r_lr_op_,decode_tv_r_sc_op_,decode_tv_r_amo_op_,decode_tv_r_clean_op_,
  decode_tv_r_inval_op_,decode_tv_r_bclean_op_,decode_tv_r_binval_op_,
  decode_tv_r_bzero_op_,decode_tv_r_amo_subop__3_,decode_tv_r_amo_subop__2_,
  decode_tv_r_amo_subop__1_,decode_tv_r_amo_subop__0_,uncached_tv_r,store_hit_tv,sc_fail_tv,
  nonblocking_req,store_miss_tv,load_miss_tv,blocking_miss_tv,nonblocking_miss_tv,
  engine_miss_tv,any_miss_tv,sc_success_tv,N169,N170,N171,N172,N173,stat_mem_v_li,
  stat_mem_w_li,wbuf_v_li,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
  N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,
  N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,
  N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,
  N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,
  N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,
  N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,
  N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,
  N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,
  N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,
  N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,
  N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,
  N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,
  N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,
  N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,
  N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,
  N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,
  N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,
  N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,
  N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,
  N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,
  N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,
  N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,
  N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,
  N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,
  N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,
  N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,
  N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,
  N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,
  N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,
  N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,
  N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,
  N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,
  N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,
  N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,
  N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,
  N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,
  N763,N764,N765,N766,N767,N768,wbuf_entry_in_bank_sel__7_,
  wbuf_entry_in_bank_sel__6_,wbuf_entry_in_bank_sel__5_,wbuf_entry_in_bank_sel__4_,
  wbuf_entry_in_bank_sel__3_,wbuf_entry_in_bank_sel__2_,wbuf_entry_in_bank_sel__1_,
  wbuf_entry_in_bank_sel__0_,wbuf_entry_in_mask__7_,wbuf_entry_in_mask__6_,wbuf_entry_in_mask__5_,
  wbuf_entry_in_mask__4_,wbuf_entry_in_mask__3_,wbuf_entry_in_mask__2_,
  wbuf_entry_in_mask__1_,wbuf_entry_in_mask__0_,wbuf_entry_in_data__63_,wbuf_entry_in_data__62_,
  wbuf_entry_in_data__61_,wbuf_entry_in_data__60_,wbuf_entry_in_data__59_,
  wbuf_entry_in_data__58_,wbuf_entry_in_data__57_,wbuf_entry_in_data__56_,
  wbuf_entry_in_data__55_,wbuf_entry_in_data__54_,wbuf_entry_in_data__53_,wbuf_entry_in_data__52_,
  wbuf_entry_in_data__51_,wbuf_entry_in_data__50_,wbuf_entry_in_data__49_,
  wbuf_entry_in_data__48_,wbuf_entry_in_data__47_,wbuf_entry_in_data__46_,
  wbuf_entry_in_data__45_,wbuf_entry_in_data__44_,wbuf_entry_in_data__43_,wbuf_entry_in_data__42_,
  wbuf_entry_in_data__41_,wbuf_entry_in_data__40_,wbuf_entry_in_data__39_,
  wbuf_entry_in_data__38_,wbuf_entry_in_data__37_,wbuf_entry_in_data__36_,
  wbuf_entry_in_data__35_,wbuf_entry_in_data__34_,wbuf_entry_in_data__33_,wbuf_entry_in_data__32_,
  wbuf_entry_in_data__31_,wbuf_entry_in_data__30_,wbuf_entry_in_data__29_,
  wbuf_entry_in_data__28_,wbuf_entry_in_data__27_,wbuf_entry_in_data__26_,
  wbuf_entry_in_data__25_,wbuf_entry_in_data__24_,wbuf_entry_in_data__23_,wbuf_entry_in_data__22_,
  wbuf_entry_in_data__21_,wbuf_entry_in_data__20_,wbuf_entry_in_data__19_,
  wbuf_entry_in_data__18_,wbuf_entry_in_data__17_,wbuf_entry_in_data__16_,
  wbuf_entry_in_data__15_,wbuf_entry_in_data__14_,wbuf_entry_in_data__13_,wbuf_entry_in_data__12_,
  wbuf_entry_in_data__11_,wbuf_entry_in_data__10_,wbuf_entry_in_data__9_,
  wbuf_entry_in_data__8_,wbuf_entry_in_data__7_,wbuf_entry_in_data__6_,
  wbuf_entry_in_data__5_,wbuf_entry_in_data__4_,wbuf_entry_in_data__3_,wbuf_entry_in_data__2_,
  wbuf_entry_in_data__1_,wbuf_entry_in_data__0_,wbuf_v_lo,wbuf_force_lo,wbuf_yumi_li,
  wbuf_entry_out_snoop_,wbuf_entry_out_bank_sel__7_,wbuf_entry_out_bank_sel__6_,
  wbuf_entry_out_bank_sel__5_,wbuf_entry_out_bank_sel__4_,wbuf_entry_out_bank_sel__3_,
  wbuf_entry_out_bank_sel__2_,wbuf_entry_out_bank_sel__1_,wbuf_entry_out_bank_sel__0_,
  wbuf_entry_out_data__63_,wbuf_entry_out_data__62_,wbuf_entry_out_data__61_,
  wbuf_entry_out_data__60_,wbuf_entry_out_data__59_,wbuf_entry_out_data__58_,
  wbuf_entry_out_data__57_,wbuf_entry_out_data__56_,wbuf_entry_out_data__55_,
  wbuf_entry_out_data__54_,wbuf_entry_out_data__53_,wbuf_entry_out_data__52_,
  wbuf_entry_out_data__51_,wbuf_entry_out_data__50_,wbuf_entry_out_data__49_,wbuf_entry_out_data__48_,
  wbuf_entry_out_data__47_,wbuf_entry_out_data__46_,wbuf_entry_out_data__45_,
  wbuf_entry_out_data__44_,wbuf_entry_out_data__43_,wbuf_entry_out_data__42_,
  wbuf_entry_out_data__41_,wbuf_entry_out_data__40_,wbuf_entry_out_data__39_,
  wbuf_entry_out_data__38_,wbuf_entry_out_data__37_,wbuf_entry_out_data__36_,
  wbuf_entry_out_data__35_,wbuf_entry_out_data__34_,wbuf_entry_out_data__33_,wbuf_entry_out_data__32_,
  wbuf_entry_out_data__31_,wbuf_entry_out_data__30_,wbuf_entry_out_data__29_,
  wbuf_entry_out_data__28_,wbuf_entry_out_data__27_,wbuf_entry_out_data__26_,
  wbuf_entry_out_data__25_,wbuf_entry_out_data__24_,wbuf_entry_out_data__23_,
  wbuf_entry_out_data__22_,wbuf_entry_out_data__21_,wbuf_entry_out_data__20_,
  wbuf_entry_out_data__19_,wbuf_entry_out_data__18_,wbuf_entry_out_data__17_,wbuf_entry_out_data__16_,
  wbuf_entry_out_data__15_,wbuf_entry_out_data__14_,wbuf_entry_out_data__13_,
  wbuf_entry_out_data__12_,wbuf_entry_out_data__11_,wbuf_entry_out_data__10_,
  wbuf_entry_out_data__9_,wbuf_entry_out_data__8_,wbuf_entry_out_data__7_,
  wbuf_entry_out_data__6_,wbuf_entry_out_data__5_,wbuf_entry_out_data__4_,wbuf_entry_out_data__3_,
  wbuf_entry_out_data__2_,wbuf_entry_out_data__1_,wbuf_entry_out_data__0_,
  wbuf_entry_out_caddr__31_,wbuf_entry_out_caddr__30_,wbuf_entry_out_caddr__29_,
  wbuf_entry_out_caddr__28_,wbuf_entry_out_caddr__27_,wbuf_entry_out_caddr__26_,
  wbuf_entry_out_caddr__25_,wbuf_entry_out_caddr__24_,wbuf_entry_out_caddr__23_,
  wbuf_entry_out_caddr__22_,wbuf_entry_out_caddr__21_,wbuf_entry_out_caddr__20_,
  wbuf_entry_out_caddr__19_,wbuf_entry_out_caddr__18_,wbuf_entry_out_caddr__17_,
  wbuf_entry_out_caddr__16_,wbuf_entry_out_caddr__15_,wbuf_entry_out_caddr__14_,
  wbuf_entry_out_caddr__13_,wbuf_entry_out_caddr__12_,wbuf_entry_out_caddr__11_,
  wbuf_entry_out_caddr__10_,wbuf_entry_out_caddr__9_,wbuf_entry_out_caddr__8_,wbuf_entry_out_caddr__7_,
  wbuf_entry_out_caddr__6_,wbuf_entry_out_caddr__5_,wbuf_entry_out_caddr__4_,
  wbuf_entry_out_caddr__3_,wbuf_entry_out_caddr__2_,wbuf_entry_out_caddr__1_,
  wbuf_entry_out_caddr__0_,wbuf_snoop_match_lo,load_req,store_req,uncached_amo_req,
  uncached_load_req,uncached_store_req,bclean_req,inval_req,clean_req,flush_req,blocking_sent,
  N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,
  N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,
  N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,
  N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,
  N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,
  N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,
  N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,
  metadata_hit_r,_14_net__7_,_14_net__6_,_14_net__5_,_14_net__4_,_14_net__3_,
  _14_net__2_,_14_net__1_,_14_net__0_,metadata_invalid_exist,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,tag_mem_fast_read,
  tag_mem_slow_read,tag_mem_slow_write,tag_mem_fast_write,N897,N898,N899,N900,N901,N902,
  N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,N918,
  N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,N934,
  N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,N950,
  N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,N966,
  N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,N982,
  N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,N998,
  N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012,
  N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,N1025,
  N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038,
  N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,
  N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,N1065,
  N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,
  N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091,N1092,
  N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,N1105,
  N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118,
  N1119,N1120,N1121,N1122,N1123,stat_mem_fast_read,stat_mem_fast_write,
  stat_mem_slow_write,stat_mem_slow_read,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  \tdm.dirty_mask_v_li ,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,
  N1143,\l1_lrsc.set_reservation ,\l1_lrsc.load_reserved_v_r ,N1144,N1145,
  \l1_lrsc.clear_reservation ,N1146,N1147,\l1_lrsc.load_reservation_match_tv ,
  \l1_lrsc.lrsc_lock_up ,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,
  N1159,N1160,\hum.fill_v ,\hum.fill_recv ,N1161,N1162,N1163,N1164,N1165,N1166,N1167,
  N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,_25_net_,N1178,
  N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,
  N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,
  N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,
  N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,
  N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,
  N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,
  N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,
  N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,
  N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,
  N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,
  N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,
  N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,
  N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,
  N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,
  N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,
  N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,
  N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,
  N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,
  N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,
  N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,
  N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,
  N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,
  N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,
  N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,
  N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,
  N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,
  N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
  N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,
  N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,
  N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,
  N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,
  N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,
  N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,
  N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,
  N1633,N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,
  N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,
  N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,
  N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,
  N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,
  N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,
  N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,
  N1726,N1727,N1728,N1729,N1730;
  wire [32:0] decode_lo,decode_tl_r,decode_tv_n,snoop_decode;
  wire [5:0] tag_mem_addr_li,stat_mem_addr_li,\l1_lrsc.load_reserved_index_r ,
  \hum.fill_index ;
  wire [183:0] tag_mem_data_li,tag_mem_mask_li,tag_mem_data_lo;
  wire [7:0] data_mem_v_li,data_mem_w_li,load_hit_tl,store_hit_tl,bank_sel_one_hot_tl,
  way_v_tv_n,store_hit_tv_n,load_hit_tv_n,bank_sel_one_hot_tv_n,snoop_bank_sel_one_hot,
  way_v_tv_r,store_hit_v_tv_r,load_hit_v_tv_r,bank_sel_one_hot_tv_r,
  ld_data_way_select_tv,\wbuf_in_0_.addr_dec ,metadata_way_v_r,tag_mem_way_one_hot,
  data_mem_pkt_fill_mask_expanded,data_mem_write_bank_mask,wbuf_data_mem_mask,
  data_mem_force_write,data_mem_slow_write,data_mem_slow_read,data_mem_fast_write,dirty_mask_lo,
  \hum.fill_bank_mask_r ,\hum.fill_bank_mask_n ,\hum.fill_hit_n ,\hum.fill_hit_r ,
  pseudo_hit;
  wire [71:0] data_mem_addr_li;
  wire [11:0] paddr_tl;
  wire [39:0] paddr_tv_n;
  wire [39:12] snoop_paddr;
  wire [2:0] store_hit_way_tv,load_hit_way_tv,lru_encode,metadata_hit_index_r,
  metadata_invalid_way,lru_way_li,tag_mem_pkt_way_r,\data_mem_lines_0_.data_mem_pkt_offset ,
  \data_mem_lines_1_.data_mem_pkt_offset ,\data_mem_lines_2_.data_mem_pkt_offset ,
  \data_mem_lines_3_.data_mem_pkt_offset ,\data_mem_lines_4_.data_mem_pkt_offset ,
  \data_mem_lines_5_.data_mem_pkt_offset ,\data_mem_lines_6_.data_mem_pkt_offset ,
  \data_mem_lines_7_.data_mem_pkt_offset ,data_mem_pkt_way_r,lru_decode_way_li,
  \tdm.dirty_mask_way_li ,stat_mem_pkt_way_r;
  wire [63:32] amo32_reg_in,amo64_reg_in;
  wire [31:0] wbuf_data_mem_mask_in,\wbuf_in_2_.slice_data ;
  wire [0:0] \wbuf_in_3_.addr_dec ,data_mem_fast_read;
  wire [127:0] data_mem_pkt_fill_data_li;
  wire [6:0] lru_decode_data_lo,lru_decode_mask_lo;
  wire [19:0] \l1_lrsc.load_reserved_tag_r ;
  reg state_r_1_sv2v_reg,state_r_0_sv2v_reg;
  assign state_r[1] = state_r_1_sv2v_reg;
  assign state_r[0] = state_r_0_sv2v_reg;
  assign cache_req_o[116] = 1'b0;

  bp_be_dcache_decoder_00_00000ffe
  pkt_decoder
  (
    .pkt_i(dcache_pkt_i),
    .decode_o(decode_lo)
  );


  bsg_mem_1rw_sync_mask_write_bit_000000b8_00000040_1
  tag_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(tag_mem_data_li),
    .addr_i(tag_mem_addr_li),
    .v_i(tag_mem_v_li),
    .w_mask_i(tag_mem_mask_li),
    .w_i(tag_mem_w_li),
    .data_o(tag_mem_data_lo)
  );


  bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
  \d_0_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li[0]),
    .w_i(data_mem_w_li[0]),
    .addr_i(data_mem_addr_li[8:0]),
    .data_i(data_mem_data_li[63:0]),
    .write_mask_i(data_mem_mask_li[7:0]),
    .data_o(data_mem_data_lo[63:0])
  );


  bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
  \d_1_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li[1]),
    .w_i(data_mem_w_li[1]),
    .addr_i(data_mem_addr_li[17:9]),
    .data_i(data_mem_data_li[127:64]),
    .write_mask_i(data_mem_mask_li[15:8]),
    .data_o(data_mem_data_lo[127:64])
  );


  bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
  \d_2_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li[2]),
    .w_i(data_mem_w_li[2]),
    .addr_i(data_mem_addr_li[26:18]),
    .data_i(data_mem_data_li[191:128]),
    .write_mask_i(data_mem_mask_li[23:16]),
    .data_o(data_mem_data_lo[191:128])
  );


  bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
  \d_3_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li[3]),
    .w_i(data_mem_w_li[3]),
    .addr_i(data_mem_addr_li[35:27]),
    .data_i(data_mem_data_li[255:192]),
    .write_mask_i(data_mem_mask_li[31:24]),
    .data_o(data_mem_data_lo[255:192])
  );


  bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
  \d_4_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li[4]),
    .w_i(data_mem_w_li[4]),
    .addr_i(data_mem_addr_li[44:36]),
    .data_i(data_mem_data_li[319:256]),
    .write_mask_i(data_mem_mask_li[39:32]),
    .data_o(data_mem_data_lo[319:256])
  );


  bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
  \d_5_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li[5]),
    .w_i(data_mem_w_li[5]),
    .addr_i(data_mem_addr_li[53:45]),
    .data_i(data_mem_data_li[383:320]),
    .write_mask_i(data_mem_mask_li[47:40]),
    .data_o(data_mem_data_lo[383:320])
  );


  bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
  \d_6_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li[6]),
    .w_i(data_mem_w_li[6]),
    .addr_i(data_mem_addr_li[62:54]),
    .data_i(data_mem_data_li[447:384]),
    .write_mask_i(data_mem_mask_li[55:48]),
    .data_o(data_mem_data_lo[447:384])
  );


  bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
  \d_7_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li[7]),
    .w_i(data_mem_w_li[7]),
    .addr_i(data_mem_addr_li[71:63]),
    .data_i(data_mem_data_li[511:448]),
    .write_mask_i(data_mem_mask_li[63:56]),
    .data_o(data_mem_data_lo[511:448])
  );


  bsg_dff_reset_width_p1
  v_tl_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(tl_we),
    .data_o(v_tl_r)
  );


  bsg_dff_width_p45
  tl_stage_reg
  (
    .clk_i(clk_i),
    .data_i({ dcache_pkt_i[11:0], decode_lo }),
    .data_o({ paddr_tl, decode_tl_r })
  );

  assign N89 = ptag_i[19:0] == tag_mem_data_lo[19:0];
  assign N90 = ~tag_mem_data_lo[22];
  assign N91 = ~tag_mem_data_lo[21];
  assign N92 = N91 | N90;
  assign N93 = tag_mem_data_lo[20] | N92;
  assign N94 = ~N93;
  assign N95 = N91 | tag_mem_data_lo[22];
  assign N96 = tag_mem_data_lo[20] | N95;
  assign N97 = ~N96;
  assign N98 = N94 | N97;
  assign N99 = ptag_i[19:0] == tag_mem_data_lo[42:23];
  assign N100 = ~tag_mem_data_lo[45];
  assign N101 = ~tag_mem_data_lo[44];
  assign N102 = N101 | N100;
  assign N103 = tag_mem_data_lo[43] | N102;
  assign N104 = ~N103;
  assign N105 = N101 | tag_mem_data_lo[45];
  assign N106 = tag_mem_data_lo[43] | N105;
  assign N107 = ~N106;
  assign N108 = N104 | N107;
  assign N109 = ptag_i[19:0] == tag_mem_data_lo[65:46];
  assign N110 = ~tag_mem_data_lo[68];
  assign N111 = ~tag_mem_data_lo[67];
  assign N112 = N111 | N110;
  assign N113 = tag_mem_data_lo[66] | N112;
  assign N114 = ~N113;
  assign N115 = N111 | tag_mem_data_lo[68];
  assign N116 = tag_mem_data_lo[66] | N115;
  assign N117 = ~N116;
  assign N118 = N114 | N117;
  assign N119 = ptag_i[19:0] == tag_mem_data_lo[88:69];
  assign N120 = ~tag_mem_data_lo[91];
  assign N121 = ~tag_mem_data_lo[90];
  assign N122 = N121 | N120;
  assign N123 = tag_mem_data_lo[89] | N122;
  assign N124 = ~N123;
  assign N125 = N121 | tag_mem_data_lo[91];
  assign N126 = tag_mem_data_lo[89] | N125;
  assign N127 = ~N126;
  assign N128 = N124 | N127;
  assign N129 = ptag_i[19:0] == tag_mem_data_lo[111:92];
  assign N130 = ~tag_mem_data_lo[114];
  assign N131 = ~tag_mem_data_lo[113];
  assign N132 = N131 | N130;
  assign N133 = tag_mem_data_lo[112] | N132;
  assign N134 = ~N133;
  assign N135 = N131 | tag_mem_data_lo[114];
  assign N136 = tag_mem_data_lo[112] | N135;
  assign N137 = ~N136;
  assign N138 = N134 | N137;
  assign N139 = ptag_i[19:0] == tag_mem_data_lo[134:115];
  assign N140 = ~tag_mem_data_lo[137];
  assign N141 = ~tag_mem_data_lo[136];
  assign N142 = N141 | N140;
  assign N143 = tag_mem_data_lo[135] | N142;
  assign N144 = ~N143;
  assign N145 = N141 | tag_mem_data_lo[137];
  assign N146 = tag_mem_data_lo[135] | N145;
  assign N147 = ~N146;
  assign N148 = N144 | N147;
  assign N149 = ptag_i[19:0] == tag_mem_data_lo[157:138];
  assign N150 = ~tag_mem_data_lo[160];
  assign N151 = ~tag_mem_data_lo[159];
  assign N152 = N151 | N150;
  assign N153 = tag_mem_data_lo[158] | N152;
  assign N154 = ~N153;
  assign N155 = N151 | tag_mem_data_lo[160];
  assign N156 = tag_mem_data_lo[158] | N155;
  assign N157 = ~N156;
  assign N158 = N154 | N157;
  assign N159 = ptag_i[19:0] == tag_mem_data_lo[180:161];
  assign N160 = ~tag_mem_data_lo[183];
  assign N161 = ~tag_mem_data_lo[182];
  assign N162 = N161 | N160;
  assign N163 = tag_mem_data_lo[181] | N162;
  assign N164 = ~N163;
  assign N165 = N161 | tag_mem_data_lo[183];
  assign N166 = tag_mem_data_lo[181] | N165;
  assign N167 = ~N166;
  assign N168 = N164 | N167;

  bsg_decode_00000008
  offset_decode
  (
    .i(paddr_tl[5:3]),
    .o(bank_sel_one_hot_tl)
  );


  bsg_dff_reset_width_p1
  v_tv_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(_2_net_),
    .data_o(v_tv_r)
  );


  bsg_mux_000002aa_2
  tv_snoop_mux
  (
    .data_i({ pseudo_hit, pseudo_hit, pseudo_hit, data_mem_data_li, snoop_st_data, snoop_paddr, \hum.fill_index , snoop_paddr_5, snoop_paddr_4, snoop_paddr_3, snoop_paddr_2, snoop_paddr_1, snoop_paddr_0, snoop_bank_sel_one_hot, snoop_uncached, snoop_decode, N1196, N1198, N1200, N1202, N1204, N1206, N1208, N1210, store_hit_tl, load_hit_tl, data_mem_data_lo, st_data_i, ptag_i, paddr_tl, bank_sel_one_hot_tl, uncached_tl, decode_tl_r }),
    .sel_i(critical_recv),
    .data_o({ way_v_tv_n, store_hit_tv_n, load_hit_tv_n, ld_data_tv_n, st_data_tv_n, paddr_tv_n, bank_sel_one_hot_tv_n, uncached_tv_n, decode_tv_n })
  );


  bsg_dff_000002ab
  tv_stage_reg
  (
    .clk_i(clk_i),
    .data_i({ critical_recv, way_v_tv_n, store_hit_tv_n, load_hit_tv_n, paddr_tv_n, ld_data_tv_n, st_data_tv_n, bank_sel_one_hot_tv_n, uncached_tv_n, decode_tv_n }),
    .data_o({ late_o, way_v_tv_r, store_hit_v_tv_r, load_hit_v_tv_r, cache_req_o[47:8], ld_data_tv_r, amo64_reg_in, amo32_reg_in, bank_sel_one_hot_tv_r, uncached_tv_r, tag_o, decode_tv_r_load_op_, ret_o, decode_tv_r_store_op_, decode_tv_r_signed_op_, float_o, int_o, ptw_o, decode_tv_r_cache_op_, decode_tv_r_block_op_, decode_tv_r_double_op_, decode_tv_r_word_op_, decode_tv_r_half_op_, decode_tv_r_byte_op_, decode_tv_r_uncached_op_, decode_tv_r_lr_op_, decode_tv_r_sc_op_, decode_tv_r_amo_op_, decode_tv_r_clean_op_, decode_tv_r_inval_op_, decode_tv_r_bclean_op_, decode_tv_r_binval_op_, decode_tv_r_bzero_op_, decode_tv_r_amo_subop__3_, decode_tv_r_amo_subop__2_, decode_tv_r_amo_subop__1_, decode_tv_r_amo_subop__0_, rd_addr_o })
  );


  bsg_encode_one_hot_00000008_1
  store_hit_index_encoder
  (
    .i(store_hit_v_tv_r),
    .addr_o(store_hit_way_tv),
    .v_o(store_hit_tv)
  );


  bsg_encode_one_hot_00000008_1
  load_hit_index_encoder
  (
    .i(load_hit_v_tv_r),
    .addr_o(load_hit_way_tv),
    .v_o(cache_req_o[115])
  );


  bsg_adder_one_hot_00000008
  select_adder
  (
    .a_i(load_hit_v_tv_r),
    .b_i(bank_sel_one_hot_tv_r),
    .o(ld_data_way_select_tv)
  );


  bsg_mux_one_hot_00000040_00000008
  ld_data_set_select_mux
  (
    .data_i(ld_data_tv_r),
    .sel_one_hot_i(ld_data_way_select_tv),
    .data_o(ld_data_way_picked)
  );


  bsg_mux_00000040_00000001
  dword_mux
  (
    .data_i(ld_data_way_picked),
    .sel_i(cache_req_o[11]),
    .data_o(ld_data_dword_raw)
  );

  assign final_data_tv = ld_data_dword_merged >> { cache_req_o[10:8], 1'b0, 1'b0, 1'b0 };

  bsg_mem_1rw_sync_mask_write_bit_0000000f_00000040_1
  stat_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(stat_mem_data_li),
    .addr_i(stat_mem_addr_li),
    .v_i(stat_mem_v_li),
    .w_mask_i(stat_mem_mask_li),
    .w_i(stat_mem_w_li),
    .data_o(stat_mem_o)
  );


  bsg_lru_pseudo_tree_encode_00000008
  lru_encoder
  (
    .lru_i(stat_mem_o[14:8]),
    .way_id_o(lru_encode)
  );

  assign N438 = $signed(atomic_reg_data) < $signed(atomic_mem_data);
  assign N504 = $signed(atomic_reg_data) > $signed(atomic_mem_data);
  assign N570 = atomic_reg_data < atomic_mem_data;
  assign N636 = atomic_reg_data > atomic_mem_data;

  bsg_decode_00000008
  \wbuf_in_0_.decode 
  (
    .i(cache_req_o[10:8]),
    .o(\wbuf_in_0_.addr_dec )
  );


  bsg_expand_bitmask_in_width_p8_expand_p1
  \wbuf_in_0_.expand 
  (
    .i(\wbuf_in_0_.addr_dec ),
    .o(wbuf_data_mem_mask_in[7:0])
  );


  bsg_decode_num_out_p4
  \wbuf_in_1_.decode 
  (
    .i(cache_req_o[10:9]),
    .o(\wbuf_in_1_.addr_dec )
  );


  bsg_expand_bitmask_in_width_p4_expand_p2
  \wbuf_in_1_.expand 
  (
    .i(\wbuf_in_1_.addr_dec ),
    .o(wbuf_data_mem_mask_in[15:8])
  );


  bsg_decode_num_out_p2
  \wbuf_in_2_.decode 
  (
    .i(cache_req_o[10]),
    .o(\wbuf_in_2_.addr_dec )
  );


  bsg_expand_bitmask_in_width_p2_expand_p4
  \wbuf_in_2_.expand 
  (
    .i(\wbuf_in_2_.addr_dec ),
    .o(wbuf_data_mem_mask_in[23:16])
  );


  bsg_decode_num_out_p1
  \wbuf_in_3_.decode 
  (
    .i(cache_req_o[11]),
    .o(\wbuf_in_3_.addr_dec [0])
  );


  bsg_expand_bitmask_in_width_p1_expand_p8
  \wbuf_in_3_.expand 
  (
    .i(\wbuf_in_3_.addr_dec [0]),
    .o(wbuf_data_mem_mask_in[31:24])
  );


  bsg_mux_one_hot_width_p64_els_p4
  wbuf_data_in_mux
  (
    .data_i({ \wbuf_in_3_.slice_data , \wbuf_in_2_.slice_data , \wbuf_in_2_.slice_data , amo32_reg_in[47:32], amo32_reg_in[47:32], amo32_reg_in[47:32], amo32_reg_in[47:32], amo32_reg_in[39:32], amo32_reg_in[39:32], amo32_reg_in[39:32], amo32_reg_in[39:32], amo32_reg_in[39:32], amo32_reg_in[39:32], amo32_reg_in[39:32], amo32_reg_in[39:32] }),
    .sel_one_hot_i({ decode_tv_r_double_op_, decode_tv_r_word_op_, decode_tv_r_half_op_, decode_tv_r_byte_op_ }),
    .data_o({ wbuf_entry_in_data__63_, wbuf_entry_in_data__62_, wbuf_entry_in_data__61_, wbuf_entry_in_data__60_, wbuf_entry_in_data__59_, wbuf_entry_in_data__58_, wbuf_entry_in_data__57_, wbuf_entry_in_data__56_, wbuf_entry_in_data__55_, wbuf_entry_in_data__54_, wbuf_entry_in_data__53_, wbuf_entry_in_data__52_, wbuf_entry_in_data__51_, wbuf_entry_in_data__50_, wbuf_entry_in_data__49_, wbuf_entry_in_data__48_, wbuf_entry_in_data__47_, wbuf_entry_in_data__46_, wbuf_entry_in_data__45_, wbuf_entry_in_data__44_, wbuf_entry_in_data__43_, wbuf_entry_in_data__42_, wbuf_entry_in_data__41_, wbuf_entry_in_data__40_, wbuf_entry_in_data__39_, wbuf_entry_in_data__38_, wbuf_entry_in_data__37_, wbuf_entry_in_data__36_, wbuf_entry_in_data__35_, wbuf_entry_in_data__34_, wbuf_entry_in_data__33_, wbuf_entry_in_data__32_, wbuf_entry_in_data__31_, wbuf_entry_in_data__30_, wbuf_entry_in_data__29_, wbuf_entry_in_data__28_, wbuf_entry_in_data__27_, wbuf_entry_in_data__26_, wbuf_entry_in_data__25_, wbuf_entry_in_data__24_, wbuf_entry_in_data__23_, wbuf_entry_in_data__22_, wbuf_entry_in_data__21_, wbuf_entry_in_data__20_, wbuf_entry_in_data__19_, wbuf_entry_in_data__18_, wbuf_entry_in_data__17_, wbuf_entry_in_data__16_, wbuf_entry_in_data__15_, wbuf_entry_in_data__14_, wbuf_entry_in_data__13_, wbuf_entry_in_data__12_, wbuf_entry_in_data__11_, wbuf_entry_in_data__10_, wbuf_entry_in_data__9_, wbuf_entry_in_data__8_, wbuf_entry_in_data__7_, wbuf_entry_in_data__6_, wbuf_entry_in_data__5_, wbuf_entry_in_data__4_, wbuf_entry_in_data__3_, wbuf_entry_in_data__2_, wbuf_entry_in_data__1_, wbuf_entry_in_data__0_ })
  );


  bsg_mux_one_hot_00000008_4
  wbuf_data_mem_mask_in_mux
  (
    .data_i(wbuf_data_mem_mask_in),
    .sel_one_hot_i({ decode_tv_r_double_op_, decode_tv_r_word_op_, decode_tv_r_half_op_, decode_tv_r_byte_op_ }),
    .data_o({ wbuf_entry_in_mask__7_, wbuf_entry_in_mask__6_, wbuf_entry_in_mask__5_, wbuf_entry_in_mask__4_, wbuf_entry_in_mask__3_, wbuf_entry_in_mask__2_, wbuf_entry_in_mask__1_, wbuf_entry_in_mask__0_ })
  );


  bp_be_dcache_wbuf_00_00000040_00000008_00000200_00000080_00000014
  wbuf
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .wbuf_entry_i({ late_o, wbuf_entry_in_bank_sel__7_, wbuf_entry_in_bank_sel__6_, wbuf_entry_in_bank_sel__5_, wbuf_entry_in_bank_sel__4_, wbuf_entry_in_bank_sel__3_, wbuf_entry_in_bank_sel__2_, wbuf_entry_in_bank_sel__1_, wbuf_entry_in_bank_sel__0_, wbuf_entry_in_mask__7_, wbuf_entry_in_mask__6_, wbuf_entry_in_mask__5_, wbuf_entry_in_mask__4_, wbuf_entry_in_mask__3_, wbuf_entry_in_mask__2_, wbuf_entry_in_mask__1_, wbuf_entry_in_mask__0_, wbuf_entry_in_data__63_, wbuf_entry_in_data__62_, wbuf_entry_in_data__61_, wbuf_entry_in_data__60_, wbuf_entry_in_data__59_, wbuf_entry_in_data__58_, wbuf_entry_in_data__57_, wbuf_entry_in_data__56_, wbuf_entry_in_data__55_, wbuf_entry_in_data__54_, wbuf_entry_in_data__53_, wbuf_entry_in_data__52_, wbuf_entry_in_data__51_, wbuf_entry_in_data__50_, wbuf_entry_in_data__49_, wbuf_entry_in_data__48_, wbuf_entry_in_data__47_, wbuf_entry_in_data__46_, wbuf_entry_in_data__45_, wbuf_entry_in_data__44_, wbuf_entry_in_data__43_, wbuf_entry_in_data__42_, wbuf_entry_in_data__41_, wbuf_entry_in_data__40_, wbuf_entry_in_data__39_, wbuf_entry_in_data__38_, wbuf_entry_in_data__37_, wbuf_entry_in_data__36_, wbuf_entry_in_data__35_, wbuf_entry_in_data__34_, wbuf_entry_in_data__33_, wbuf_entry_in_data__32_, wbuf_entry_in_data__31_, wbuf_entry_in_data__30_, wbuf_entry_in_data__29_, wbuf_entry_in_data__28_, wbuf_entry_in_data__27_, wbuf_entry_in_data__26_, wbuf_entry_in_data__25_, wbuf_entry_in_data__24_, wbuf_entry_in_data__23_, wbuf_entry_in_data__22_, wbuf_entry_in_data__21_, wbuf_entry_in_data__20_, wbuf_entry_in_data__19_, wbuf_entry_in_data__18_, wbuf_entry_in_data__17_, wbuf_entry_in_data__16_, wbuf_entry_in_data__15_, wbuf_entry_in_data__14_, wbuf_entry_in_data__13_, wbuf_entry_in_data__12_, wbuf_entry_in_data__11_, wbuf_entry_in_data__10_, wbuf_entry_in_data__9_, wbuf_entry_in_data__8_, wbuf_entry_in_data__7_, wbuf_entry_in_data__6_, wbuf_entry_in_data__5_, wbuf_entry_in_data__4_, wbuf_entry_in_data__3_, wbuf_entry_in_data__2_, wbuf_entry_in_data__1_, wbuf_entry_in_data__0_, cache_req_o[39:8] }),
    .v_i(wbuf_v_li),
    .wbuf_entry_o({ wbuf_entry_out_snoop_, wbuf_entry_out_bank_sel__7_, wbuf_entry_out_bank_sel__6_, wbuf_entry_out_bank_sel__5_, wbuf_entry_out_bank_sel__4_, wbuf_entry_out_bank_sel__3_, wbuf_entry_out_bank_sel__2_, wbuf_entry_out_bank_sel__1_, wbuf_entry_out_bank_sel__0_, wbuf_data_mem_mask, wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_, wbuf_entry_out_caddr__31_, wbuf_entry_out_caddr__30_, wbuf_entry_out_caddr__29_, wbuf_entry_out_caddr__28_, wbuf_entry_out_caddr__27_, wbuf_entry_out_caddr__26_, wbuf_entry_out_caddr__25_, wbuf_entry_out_caddr__24_, wbuf_entry_out_caddr__23_, wbuf_entry_out_caddr__22_, wbuf_entry_out_caddr__21_, wbuf_entry_out_caddr__20_, wbuf_entry_out_caddr__19_, wbuf_entry_out_caddr__18_, wbuf_entry_out_caddr__17_, wbuf_entry_out_caddr__16_, wbuf_entry_out_caddr__15_, wbuf_entry_out_caddr__14_, wbuf_entry_out_caddr__13_, wbuf_entry_out_caddr__12_, wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_, wbuf_entry_out_caddr__2_, wbuf_entry_out_caddr__1_, wbuf_entry_out_caddr__0_ }),
    .v_o(wbuf_v_lo),
    .force_o(wbuf_force_lo),
    .yumi_i(wbuf_yumi_li),
    .data_mem_pkt_i(data_mem_pkt_i),
    .data_mem_pkt_v_i(data_mem_pkt_v_i),
    .tag_mem_pkt_i(tag_mem_pkt_i),
    .tag_mem_pkt_v_i(tag_mem_pkt_v_i),
    .stat_mem_pkt_i(stat_mem_pkt_i),
    .stat_mem_pkt_v_i(stat_mem_pkt_v_i),
    .snoop_match_o(wbuf_snoop_match_lo),
    .v_tl_i(v_tl_r),
    .addr_tl_i({ ptag_i[19:0], paddr_tl }),
    .data_tv_i(ld_data_dword_raw),
    .data_merged_o(ld_data_dword_merged)
  );

  assign N784 = decode_tv_r_amo_subop__3_ | decode_tv_r_amo_subop__2_;
  assign N785 = decode_tv_r_amo_subop__1_ | N783;
  assign N786 = N784 | N785;
  assign N789 = N788 | decode_tv_r_amo_subop__0_;
  assign N790 = N784 | N789;
  assign N792 = N788 | N783;
  assign N793 = N784 | N792;
  assign N796 = decode_tv_r_amo_subop__3_ | N795;
  assign N797 = decode_tv_r_amo_subop__1_ | decode_tv_r_amo_subop__0_;
  assign N798 = N796 | N797;
  assign N800 = N796 | N785;
  assign N802 = N796 | N789;
  assign N804 = N796 | N792;
  assign N807 = N806 | decode_tv_r_amo_subop__2_;
  assign N808 = N807 | N797;
  assign N810 = N807 | N785;
  assign N812 = N807 | N789;
  assign N814 = N807 | N792;
  assign N816 = decode_tv_r_amo_subop__3_ & decode_tv_r_amo_subop__2_;
  assign N817 = N806 & N795;
  assign N818 = N788 & N783;
  assign N819 = N817 & N818;

  bsg_dff_reset_width_p1
  cache_req_v_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(cache_req_yumi_i),
    .data_o(cache_req_metadata_v_o)
  );


  bsg_dff_0000000c
  cached_hit_reg
  (
    .clk_i(clk_i),
    .data_i({ way_v_tv_r, cache_req_o[115:115], load_hit_way_tv }),
    .data_o({ metadata_way_v_r, metadata_hit_r, metadata_hit_index_r })
  );


  bsg_priority_encode_00000008_1
  pe_invalid
  (
    .i({ _14_net__7_, _14_net__6_, _14_net__5_, _14_net__4_, _14_net__3_, _14_net__2_, _14_net__1_, _14_net__0_ }),
    .addr_o(metadata_invalid_way),
    .v_o(metadata_invalid_exist)
  );

  assign cache_req_metadata_o[0] = (N889)? stat_mem_o[0] : 
                                   (N891)? stat_mem_o[1] : 
                                   (N893)? stat_mem_o[2] : 
                                   (N895)? stat_mem_o[3] : 
                                   (N890)? stat_mem_o[4] : 
                                   (N892)? stat_mem_o[5] : 
                                   (N894)? stat_mem_o[6] : 
                                   (N896)? stat_mem_o[7] : 1'b0;

  bsg_decode_00000008
  tag_mem_way_decode
  (
    .i(tag_mem_pkt_i[28:26]),
    .o(tag_mem_way_one_hot)
  );

  assign N902 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N903 = tag_mem_pkt_i[1] | N901;
  assign N904 = N902 | N903;
  assign N907 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N908 = N906 | tag_mem_pkt_i[0];
  assign N909 = N907 | N908;
  assign N913 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N914 = N911 | N912;
  assign N915 = N913 | N914;
  assign N917 = N1529 & tag_mem_pkt_i[2];
  assign N920 = N1529 & N918;
  assign N921 = N920 & N919;
  assign N924 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N925 = tag_mem_pkt_i[1] | N923;
  assign N926 = N924 | N925;
  assign N929 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N930 = N928 | tag_mem_pkt_i[0];
  assign N931 = N929 | N930;
  assign N935 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N936 = N933 | N934;
  assign N937 = N935 | N936;
  assign N939 = N1529 & tag_mem_pkt_i[2];
  assign N942 = N1529 & N940;
  assign N943 = N942 & N941;
  assign N946 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N947 = tag_mem_pkt_i[1] | N945;
  assign N948 = N946 | N947;
  assign N951 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N952 = N950 | tag_mem_pkt_i[0];
  assign N953 = N951 | N952;
  assign N957 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N958 = N955 | N956;
  assign N959 = N957 | N958;
  assign N961 = N1529 & tag_mem_pkt_i[2];
  assign N964 = N1529 & N962;
  assign N965 = N964 & N963;
  assign N968 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N969 = tag_mem_pkt_i[1] | N967;
  assign N970 = N968 | N969;
  assign N973 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N974 = N972 | tag_mem_pkt_i[0];
  assign N975 = N973 | N974;
  assign N979 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N980 = N977 | N978;
  assign N981 = N979 | N980;
  assign N983 = N1529 & tag_mem_pkt_i[2];
  assign N986 = N1529 & N984;
  assign N987 = N986 & N985;
  assign N990 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N991 = tag_mem_pkt_i[1] | N989;
  assign N992 = N990 | N991;
  assign N995 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N996 = N994 | tag_mem_pkt_i[0];
  assign N997 = N995 | N996;
  assign N1001 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1002 = N999 | N1000;
  assign N1003 = N1001 | N1002;
  assign N1005 = N1529 & tag_mem_pkt_i[2];
  assign N1008 = N1529 & N1006;
  assign N1009 = N1008 & N1007;
  assign N1012 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1013 = tag_mem_pkt_i[1] | N1011;
  assign N1014 = N1012 | N1013;
  assign N1017 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1018 = N1016 | tag_mem_pkt_i[0];
  assign N1019 = N1017 | N1018;
  assign N1023 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1024 = N1021 | N1022;
  assign N1025 = N1023 | N1024;
  assign N1027 = N1529 & tag_mem_pkt_i[2];
  assign N1030 = N1529 & N1028;
  assign N1031 = N1030 & N1029;
  assign N1034 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1035 = tag_mem_pkt_i[1] | N1033;
  assign N1036 = N1034 | N1035;
  assign N1039 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1040 = N1038 | tag_mem_pkt_i[0];
  assign N1041 = N1039 | N1040;
  assign N1045 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1046 = N1043 | N1044;
  assign N1047 = N1045 | N1046;
  assign N1049 = N1529 & tag_mem_pkt_i[2];
  assign N1052 = N1529 & N1050;
  assign N1053 = N1052 & N1051;
  assign N1056 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1057 = tag_mem_pkt_i[1] | N1055;
  assign N1058 = N1056 | N1057;
  assign N1061 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1062 = N1060 | tag_mem_pkt_i[0];
  assign N1063 = N1061 | N1062;
  assign N1067 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1068 = N1065 | N1066;
  assign N1069 = N1067 | N1068;
  assign N1071 = N1529 & tag_mem_pkt_i[2];
  assign N1074 = N1529 & N1072;
  assign N1075 = N1074 & N1073;

  bsg_dff_00000003
  tag_mem_pkt_way_reg
  (
    .clk_i(clk_i),
    .data_i(tag_mem_pkt_i[28:26]),
    .data_o(tag_mem_pkt_way_r)
  );

  assign tag_mem_o[22] = (N1084)? tag_mem_data_lo[22] : 
                         (N1086)? tag_mem_data_lo[45] : 
                         (N1088)? tag_mem_data_lo[68] : 
                         (N1090)? tag_mem_data_lo[91] : 
                         (N1085)? tag_mem_data_lo[114] : 
                         (N1087)? tag_mem_data_lo[137] : 
                         (N1089)? tag_mem_data_lo[160] : 
                         (N1091)? tag_mem_data_lo[183] : 1'b0;
  assign tag_mem_o[21] = (N1084)? tag_mem_data_lo[21] : 
                         (N1086)? tag_mem_data_lo[44] : 
                         (N1088)? tag_mem_data_lo[67] : 
                         (N1090)? tag_mem_data_lo[90] : 
                         (N1085)? tag_mem_data_lo[113] : 
                         (N1087)? tag_mem_data_lo[136] : 
                         (N1089)? tag_mem_data_lo[159] : 
                         (N1091)? tag_mem_data_lo[182] : 1'b0;
  assign tag_mem_o[20] = (N1084)? tag_mem_data_lo[20] : 
                         (N1086)? tag_mem_data_lo[43] : 
                         (N1088)? tag_mem_data_lo[66] : 
                         (N1090)? tag_mem_data_lo[89] : 
                         (N1085)? tag_mem_data_lo[112] : 
                         (N1087)? tag_mem_data_lo[135] : 
                         (N1089)? tag_mem_data_lo[158] : 
                         (N1091)? tag_mem_data_lo[181] : 1'b0;
  assign tag_mem_o[19] = (N1084)? tag_mem_data_lo[19] : 
                         (N1086)? tag_mem_data_lo[42] : 
                         (N1088)? tag_mem_data_lo[65] : 
                         (N1090)? tag_mem_data_lo[88] : 
                         (N1085)? tag_mem_data_lo[111] : 
                         (N1087)? tag_mem_data_lo[134] : 
                         (N1089)? tag_mem_data_lo[157] : 
                         (N1091)? tag_mem_data_lo[180] : 1'b0;
  assign tag_mem_o[18] = (N1084)? tag_mem_data_lo[18] : 
                         (N1086)? tag_mem_data_lo[41] : 
                         (N1088)? tag_mem_data_lo[64] : 
                         (N1090)? tag_mem_data_lo[87] : 
                         (N1085)? tag_mem_data_lo[110] : 
                         (N1087)? tag_mem_data_lo[133] : 
                         (N1089)? tag_mem_data_lo[156] : 
                         (N1091)? tag_mem_data_lo[179] : 1'b0;
  assign tag_mem_o[17] = (N1084)? tag_mem_data_lo[17] : 
                         (N1086)? tag_mem_data_lo[40] : 
                         (N1088)? tag_mem_data_lo[63] : 
                         (N1090)? tag_mem_data_lo[86] : 
                         (N1085)? tag_mem_data_lo[109] : 
                         (N1087)? tag_mem_data_lo[132] : 
                         (N1089)? tag_mem_data_lo[155] : 
                         (N1091)? tag_mem_data_lo[178] : 1'b0;
  assign tag_mem_o[16] = (N1084)? tag_mem_data_lo[16] : 
                         (N1086)? tag_mem_data_lo[39] : 
                         (N1088)? tag_mem_data_lo[62] : 
                         (N1090)? tag_mem_data_lo[85] : 
                         (N1085)? tag_mem_data_lo[108] : 
                         (N1087)? tag_mem_data_lo[131] : 
                         (N1089)? tag_mem_data_lo[154] : 
                         (N1091)? tag_mem_data_lo[177] : 1'b0;
  assign tag_mem_o[15] = (N1084)? tag_mem_data_lo[15] : 
                         (N1086)? tag_mem_data_lo[38] : 
                         (N1088)? tag_mem_data_lo[61] : 
                         (N1090)? tag_mem_data_lo[84] : 
                         (N1085)? tag_mem_data_lo[107] : 
                         (N1087)? tag_mem_data_lo[130] : 
                         (N1089)? tag_mem_data_lo[153] : 
                         (N1091)? tag_mem_data_lo[176] : 1'b0;
  assign tag_mem_o[14] = (N1084)? tag_mem_data_lo[14] : 
                         (N1086)? tag_mem_data_lo[37] : 
                         (N1088)? tag_mem_data_lo[60] : 
                         (N1090)? tag_mem_data_lo[83] : 
                         (N1085)? tag_mem_data_lo[106] : 
                         (N1087)? tag_mem_data_lo[129] : 
                         (N1089)? tag_mem_data_lo[152] : 
                         (N1091)? tag_mem_data_lo[175] : 1'b0;
  assign tag_mem_o[13] = (N1084)? tag_mem_data_lo[13] : 
                         (N1086)? tag_mem_data_lo[36] : 
                         (N1088)? tag_mem_data_lo[59] : 
                         (N1090)? tag_mem_data_lo[82] : 
                         (N1085)? tag_mem_data_lo[105] : 
                         (N1087)? tag_mem_data_lo[128] : 
                         (N1089)? tag_mem_data_lo[151] : 
                         (N1091)? tag_mem_data_lo[174] : 1'b0;
  assign tag_mem_o[12] = (N1084)? tag_mem_data_lo[12] : 
                         (N1086)? tag_mem_data_lo[35] : 
                         (N1088)? tag_mem_data_lo[58] : 
                         (N1090)? tag_mem_data_lo[81] : 
                         (N1085)? tag_mem_data_lo[104] : 
                         (N1087)? tag_mem_data_lo[127] : 
                         (N1089)? tag_mem_data_lo[150] : 
                         (N1091)? tag_mem_data_lo[173] : 1'b0;
  assign tag_mem_o[11] = (N1084)? tag_mem_data_lo[11] : 
                         (N1086)? tag_mem_data_lo[34] : 
                         (N1088)? tag_mem_data_lo[57] : 
                         (N1090)? tag_mem_data_lo[80] : 
                         (N1085)? tag_mem_data_lo[103] : 
                         (N1087)? tag_mem_data_lo[126] : 
                         (N1089)? tag_mem_data_lo[149] : 
                         (N1091)? tag_mem_data_lo[172] : 1'b0;
  assign tag_mem_o[10] = (N1084)? tag_mem_data_lo[10] : 
                         (N1086)? tag_mem_data_lo[33] : 
                         (N1088)? tag_mem_data_lo[56] : 
                         (N1090)? tag_mem_data_lo[79] : 
                         (N1085)? tag_mem_data_lo[102] : 
                         (N1087)? tag_mem_data_lo[125] : 
                         (N1089)? tag_mem_data_lo[148] : 
                         (N1091)? tag_mem_data_lo[171] : 1'b0;
  assign tag_mem_o[9] = (N1084)? tag_mem_data_lo[9] : 
                        (N1086)? tag_mem_data_lo[32] : 
                        (N1088)? tag_mem_data_lo[55] : 
                        (N1090)? tag_mem_data_lo[78] : 
                        (N1085)? tag_mem_data_lo[101] : 
                        (N1087)? tag_mem_data_lo[124] : 
                        (N1089)? tag_mem_data_lo[147] : 
                        (N1091)? tag_mem_data_lo[170] : 1'b0;
  assign tag_mem_o[8] = (N1084)? tag_mem_data_lo[8] : 
                        (N1086)? tag_mem_data_lo[31] : 
                        (N1088)? tag_mem_data_lo[54] : 
                        (N1090)? tag_mem_data_lo[77] : 
                        (N1085)? tag_mem_data_lo[100] : 
                        (N1087)? tag_mem_data_lo[123] : 
                        (N1089)? tag_mem_data_lo[146] : 
                        (N1091)? tag_mem_data_lo[169] : 1'b0;
  assign tag_mem_o[7] = (N1084)? tag_mem_data_lo[7] : 
                        (N1086)? tag_mem_data_lo[30] : 
                        (N1088)? tag_mem_data_lo[53] : 
                        (N1090)? tag_mem_data_lo[76] : 
                        (N1085)? tag_mem_data_lo[99] : 
                        (N1087)? tag_mem_data_lo[122] : 
                        (N1089)? tag_mem_data_lo[145] : 
                        (N1091)? tag_mem_data_lo[168] : 1'b0;
  assign tag_mem_o[6] = (N1084)? tag_mem_data_lo[6] : 
                        (N1086)? tag_mem_data_lo[29] : 
                        (N1088)? tag_mem_data_lo[52] : 
                        (N1090)? tag_mem_data_lo[75] : 
                        (N1085)? tag_mem_data_lo[98] : 
                        (N1087)? tag_mem_data_lo[121] : 
                        (N1089)? tag_mem_data_lo[144] : 
                        (N1091)? tag_mem_data_lo[167] : 1'b0;
  assign tag_mem_o[5] = (N1084)? tag_mem_data_lo[5] : 
                        (N1086)? tag_mem_data_lo[28] : 
                        (N1088)? tag_mem_data_lo[51] : 
                        (N1090)? tag_mem_data_lo[74] : 
                        (N1085)? tag_mem_data_lo[97] : 
                        (N1087)? tag_mem_data_lo[120] : 
                        (N1089)? tag_mem_data_lo[143] : 
                        (N1091)? tag_mem_data_lo[166] : 1'b0;
  assign tag_mem_o[4] = (N1084)? tag_mem_data_lo[4] : 
                        (N1086)? tag_mem_data_lo[27] : 
                        (N1088)? tag_mem_data_lo[50] : 
                        (N1090)? tag_mem_data_lo[73] : 
                        (N1085)? tag_mem_data_lo[96] : 
                        (N1087)? tag_mem_data_lo[119] : 
                        (N1089)? tag_mem_data_lo[142] : 
                        (N1091)? tag_mem_data_lo[165] : 1'b0;
  assign tag_mem_o[3] = (N1084)? tag_mem_data_lo[3] : 
                        (N1086)? tag_mem_data_lo[26] : 
                        (N1088)? tag_mem_data_lo[49] : 
                        (N1090)? tag_mem_data_lo[72] : 
                        (N1085)? tag_mem_data_lo[95] : 
                        (N1087)? tag_mem_data_lo[118] : 
                        (N1089)? tag_mem_data_lo[141] : 
                        (N1091)? tag_mem_data_lo[164] : 1'b0;
  assign tag_mem_o[2] = (N1084)? tag_mem_data_lo[2] : 
                        (N1086)? tag_mem_data_lo[25] : 
                        (N1088)? tag_mem_data_lo[48] : 
                        (N1090)? tag_mem_data_lo[71] : 
                        (N1085)? tag_mem_data_lo[94] : 
                        (N1087)? tag_mem_data_lo[117] : 
                        (N1089)? tag_mem_data_lo[140] : 
                        (N1091)? tag_mem_data_lo[163] : 1'b0;
  assign tag_mem_o[1] = (N1084)? tag_mem_data_lo[1] : 
                        (N1086)? tag_mem_data_lo[24] : 
                        (N1088)? tag_mem_data_lo[47] : 
                        (N1090)? tag_mem_data_lo[70] : 
                        (N1085)? tag_mem_data_lo[93] : 
                        (N1087)? tag_mem_data_lo[116] : 
                        (N1089)? tag_mem_data_lo[139] : 
                        (N1091)? tag_mem_data_lo[162] : 1'b0;
  assign tag_mem_o[0] = (N1084)? tag_mem_data_lo[0] : 
                        (N1086)? tag_mem_data_lo[23] : 
                        (N1088)? tag_mem_data_lo[46] : 
                        (N1090)? tag_mem_data_lo[69] : 
                        (N1085)? tag_mem_data_lo[92] : 
                        (N1087)? tag_mem_data_lo[115] : 
                        (N1089)? tag_mem_data_lo[138] : 
                        (N1091)? tag_mem_data_lo[161] : 1'b0;

  bsg_expand_bitmask_in_width_p4_expand_p2
  fill_mask_expand
  (
    .i(data_mem_pkt_i[5:2]),
    .o(data_mem_pkt_fill_mask_expanded)
  );


  bsg_rotate_left_00000008
  write_mask_rotate
  (
    .data_i(data_mem_pkt_fill_mask_expanded),
    .rot_i(data_mem_pkt_i[136:134]),
    .o(data_mem_write_bank_mask)
  );


  bsg_rotate_left_00000080
  write_data_rotate
  (
    .data_i(data_mem_pkt_i[133:6]),
    .rot_i({ data_mem_pkt_i[134:134], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .o(data_mem_pkt_fill_data_li)
  );


  bsg_dff_00000003
  data_mem_pkt_way_reg
  (
    .clk_i(clk_i),
    .data_i(data_mem_pkt_i[136:134]),
    .data_o(data_mem_pkt_way_r)
  );


  bsg_rotate_right_00000200
  read_data_rotate
  (
    .data_i(data_mem_data_lo),
    .rot_i({ data_mem_pkt_way_r, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .o(data_mem_o)
  );


  bsg_lru_pseudo_tree_decode_00000008
  lru_decode
  (
    .way_id_i(lru_decode_way_li),
    .data_o(lru_decode_data_lo),
    .mask_o(lru_decode_mask_lo)
  );


  bsg_decode_with_v_00000008
  \tdm.dirty_mask_decode 
  (
    .i(\tdm.dirty_mask_way_li ),
    .v_i(\tdm.dirty_mask_v_li ),
    .o(dirty_mask_lo)
  );

  assign N1132 = N1513 & N1131;

  bsg_dff_00000003
  stat_mem_pkt_way_reg
  (
    .clk_i(clk_i),
    .data_i(stat_mem_pkt_i[4:2]),
    .data_o(stat_mem_pkt_way_r)
  );

  assign N1144 = tag_mem_pkt_i[34:29] == \l1_lrsc.load_reserved_index_r ;
  assign N1145 = tag_mem_pkt_i[22:3] == \l1_lrsc.load_reserved_tag_r ;

  bsg_dff_reset_set_clear_width_p1_clear_over_set_p1
  \l1_lrsc.load_reserved_v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .set_i(\l1_lrsc.set_reservation ),
    .clear_i(\l1_lrsc.clear_reservation ),
    .data_o(\l1_lrsc.load_reserved_v_r )
  );


  bsg_dff_en_0000001a
  \l1_lrsc.load_reserved_addr 
  (
    .clk_i(clk_i),
    .data_i(cache_req_o[39:14]),
    .en_i(\l1_lrsc.set_reservation ),
    .data_o({ \l1_lrsc.load_reserved_tag_r , \l1_lrsc.load_reserved_index_r  })
  );

  assign N1146 = \l1_lrsc.load_reserved_index_r  == cache_req_o[19:14];
  assign N1147 = \l1_lrsc.load_reserved_tag_r  == cache_req_o[39:20];

  bsg_counter_clear_up_max_val_p15_init_val_p0_disable_overflow_warning_p1
  \l1_lrsc.lrsc_lock_counter 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(sc_success_tv),
    .up_i(\l1_lrsc.lrsc_lock_up ),
    .count_o(\l1_lrsc.lrsc_lock_cnt )
  );


  bsg_dff_en_0000008a
  mshr_reg
  (
    .clk_i(clk_i),
    .data_i({ uncached_tv_r, amo64_reg_in, amo32_reg_in, cache_req_o[47:8], tag_o, decode_tv_r_load_op_, ret_o, decode_tv_r_store_op_, decode_tv_r_signed_op_, float_o, int_o, ptw_o, decode_tv_r_cache_op_, decode_tv_r_block_op_, decode_tv_r_double_op_, decode_tv_r_word_op_, decode_tv_r_half_op_, decode_tv_r_byte_op_, decode_tv_r_uncached_op_, decode_tv_r_lr_op_, decode_tv_r_sc_op_, decode_tv_r_amo_op_, decode_tv_r_clean_op_, decode_tv_r_inval_op_, decode_tv_r_bclean_op_, decode_tv_r_binval_op_, decode_tv_r_bzero_op_, decode_tv_r_amo_subop__3_, decode_tv_r_amo_subop__2_, decode_tv_r_amo_subop__1_, decode_tv_r_amo_subop__0_, rd_addr_o }),
    .en_i(blocking_sent),
    .data_o({ snoop_uncached, snoop_st_data, snoop_paddr, \hum.fill_index , snoop_paddr_5, snoop_paddr_4, snoop_paddr_3, snoop_paddr_2, snoop_paddr_1, snoop_paddr_0, snoop_decode })
  );

  assign { N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << data_mem_pkt_i[136:134];

  bsg_dff_reset_en_00000010
  \hum.fill_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(_25_net_),
    .data_i({ \hum.fill_bank_mask_n , \hum.fill_hit_n  }),
    .data_o({ \hum.fill_bank_mask_r , \hum.fill_hit_r  })
  );

  assign N1178 = \hum.fill_index  == paddr_tl[11:6];
  assign { N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, data_mem_pkt_v_i } << data_mem_pkt_i[136:134];
  assign { N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tag_mem_pkt_v_i } << tag_mem_pkt_i[28:26];

  bsg_decode_00000008
  snoop_offset_decode
  (
    .i({ snoop_paddr_5, snoop_paddr_4, snoop_paddr_3 }),
    .o(snoop_bank_sel_one_hot)
  );

  assign N1195 = tag_mem_data_lo[182] | tag_mem_data_lo[183];
  assign N1196 = tag_mem_data_lo[181] | N1195;
  assign N1197 = tag_mem_data_lo[159] | tag_mem_data_lo[160];
  assign N1198 = tag_mem_data_lo[158] | N1197;
  assign N1199 = tag_mem_data_lo[136] | tag_mem_data_lo[137];
  assign N1200 = tag_mem_data_lo[135] | N1199;
  assign N1201 = tag_mem_data_lo[113] | tag_mem_data_lo[114];
  assign N1202 = tag_mem_data_lo[112] | N1201;
  assign N1203 = tag_mem_data_lo[90] | tag_mem_data_lo[91];
  assign N1204 = tag_mem_data_lo[89] | N1203;
  assign N1205 = tag_mem_data_lo[67] | tag_mem_data_lo[68];
  assign N1206 = tag_mem_data_lo[66] | N1205;
  assign N1207 = tag_mem_data_lo[44] | tag_mem_data_lo[45];
  assign N1208 = tag_mem_data_lo[43] | N1207;
  assign N1209 = tag_mem_data_lo[21] | tag_mem_data_lo[22];
  assign N1210 = tag_mem_data_lo[20] | N1209;
  assign N1211 = load_hit_way_tv[1] & load_hit_way_tv[2];
  assign N1212 = load_hit_way_tv[0] & N1211;
  assign N1213 = ~load_hit_way_tv[2];
  assign N1214 = ~load_hit_way_tv[1];
  assign N1215 = N1214 | N1213;
  assign N1216 = load_hit_way_tv[0] | N1215;
  assign N1217 = ~N1216;
  assign N1218 = ~load_hit_way_tv[2];
  assign N1219 = ~load_hit_way_tv[0];
  assign N1220 = load_hit_way_tv[1] | N1218;
  assign N1221 = N1219 | N1220;
  assign N1222 = ~N1221;
  assign N1223 = ~load_hit_way_tv[2];
  assign N1224 = load_hit_way_tv[1] | N1223;
  assign N1225 = load_hit_way_tv[0] | N1224;
  assign N1226 = ~N1225;
  assign N1227 = ~load_hit_way_tv[1];
  assign N1228 = ~load_hit_way_tv[0];
  assign N1229 = N1227 | load_hit_way_tv[2];
  assign N1230 = N1228 | N1229;
  assign N1231 = ~N1230;
  assign N1232 = ~load_hit_way_tv[1];
  assign N1233 = N1232 | load_hit_way_tv[2];
  assign N1234 = load_hit_way_tv[0] | N1233;
  assign N1235 = ~N1234;
  assign N1236 = ~load_hit_way_tv[0];
  assign N1237 = load_hit_way_tv[1] | load_hit_way_tv[2];
  assign N1238 = N1236 | N1237;
  assign N1239 = ~N1238;
  assign N1240 = load_hit_way_tv[1] | load_hit_way_tv[2];
  assign N1241 = load_hit_way_tv[0] | N1240;
  assign N1242 = ~N1241;
  assign N1243 = ~tag_mem_pkt_i[2];
  assign N1244 = tag_mem_pkt_i[1] | N1243;
  assign N1245 = tag_mem_pkt_i[0] | N1244;
  assign N1246 = ~N1245;
  assign N1247 = ~tag_mem_pkt_i[2];
  assign N1248 = tag_mem_pkt_i[1] | N1247;
  assign N1249 = tag_mem_pkt_i[0] | N1248;
  assign N1250 = ~data_mem_pkt_i[0];
  assign N1251 = N1250 | data_mem_pkt_i[1];
  assign N1252 = ~N1251;
  assign N1253 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1254 = ~N1253;
  assign N1255 = ~data_mem_pkt_i[0];
  assign N1256 = N1255 | data_mem_pkt_i[1];
  assign N1257 = ~N1256;
  assign N1258 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1259 = ~N1258;
  assign N1260 = ~data_mem_pkt_i[0];
  assign N1261 = N1260 | data_mem_pkt_i[1];
  assign N1262 = ~N1261;
  assign N1263 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1264 = ~N1263;
  assign N1265 = ~data_mem_pkt_i[0];
  assign N1266 = N1265 | data_mem_pkt_i[1];
  assign N1267 = ~N1266;
  assign N1268 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1269 = ~N1268;
  assign N1270 = ~data_mem_pkt_i[0];
  assign N1271 = N1270 | data_mem_pkt_i[1];
  assign N1272 = ~N1271;
  assign N1273 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1274 = ~N1273;
  assign N1275 = ~data_mem_pkt_i[0];
  assign N1276 = N1275 | data_mem_pkt_i[1];
  assign N1277 = ~N1276;
  assign N1278 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1279 = ~N1278;
  assign N1280 = ~data_mem_pkt_i[0];
  assign N1281 = N1280 | data_mem_pkt_i[1];
  assign N1282 = ~N1281;
  assign N1283 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1284 = ~N1283;
  assign N1285 = ~data_mem_pkt_i[0];
  assign N1286 = N1285 | data_mem_pkt_i[1];
  assign N1287 = ~N1286;
  assign N1288 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1289 = ~N1288;
  assign N1290 = ~stat_mem_pkt_i[0];
  assign N1291 = N1290 | stat_mem_pkt_i[1];
  assign N1292 = ~N1291;
  assign N1293 = ~stat_mem_pkt_i[0];
  assign N1294 = N1293 | stat_mem_pkt_i[1];
  assign N1295 = tag_mem_data_lo[182] | tag_mem_data_lo[183];
  assign N1296 = tag_mem_data_lo[181] | N1295;
  assign N1297 = tag_mem_data_lo[159] | tag_mem_data_lo[160];
  assign N1298 = tag_mem_data_lo[158] | N1297;
  assign N1299 = tag_mem_data_lo[136] | tag_mem_data_lo[137];
  assign N1300 = tag_mem_data_lo[135] | N1299;
  assign N1301 = tag_mem_data_lo[113] | tag_mem_data_lo[114];
  assign N1302 = tag_mem_data_lo[112] | N1301;
  assign N1303 = tag_mem_data_lo[90] | tag_mem_data_lo[91];
  assign N1304 = tag_mem_data_lo[89] | N1303;
  assign N1305 = tag_mem_data_lo[67] | tag_mem_data_lo[68];
  assign N1306 = tag_mem_data_lo[66] | N1305;
  assign N1307 = tag_mem_data_lo[44] | tag_mem_data_lo[45];
  assign N1308 = tag_mem_data_lo[43] | N1307;
  assign N1309 = tag_mem_data_lo[21] | tag_mem_data_lo[22];
  assign N1310 = tag_mem_data_lo[20] | N1309;
  assign N1311 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1312 = ~N1311;
  assign N1313 = ~stat_mem_pkt_i[0];
  assign N1314 = N1313 | stat_mem_pkt_i[1];
  assign N1315 = ~N1314;
  assign N1316 = \l1_lrsc.lrsc_lock_cnt [2] | \l1_lrsc.lrsc_lock_cnt [3];
  assign N1317 = \l1_lrsc.lrsc_lock_cnt [1] | N1316;
  assign N1318 = \l1_lrsc.lrsc_lock_cnt [0] | N1317;
  assign N1319 = ~data_mem_pkt_i[0];
  assign N1320 = N1319 | data_mem_pkt_i[1];
  assign N1321 = ~N1320;
  assign N1322 = ~data_mem_pkt_i[0];
  assign N1323 = N1322 | data_mem_pkt_i[1];
  assign N1324 = ~N1323;
  assign N1325 = state_r[0] | state_r[1];
  assign N1326 = ~N1325;
  assign N1327 = ~state_r[0];
  assign N1328 = N1327 | state_r[1];
  assign N1329 = ~N1328;
  assign \data_mem_lines_0_.data_mem_pkt_offset  = 1'b0 - data_mem_pkt_i[136:134];
  assign \data_mem_lines_1_.data_mem_pkt_offset  = 1'b1 - data_mem_pkt_i[136:134];
  assign \data_mem_lines_2_.data_mem_pkt_offset  = { 1'b1, 1'b0 } - data_mem_pkt_i[136:134];
  assign \data_mem_lines_3_.data_mem_pkt_offset  = { 1'b1, 1'b1 } - data_mem_pkt_i[136:134];
  assign \data_mem_lines_4_.data_mem_pkt_offset  = { 1'b1, 1'b0, 1'b0 } - data_mem_pkt_i[136:134];
  assign \data_mem_lines_5_.data_mem_pkt_offset  = { 1'b1, 1'b0, 1'b1 } - data_mem_pkt_i[136:134];
  assign \data_mem_lines_6_.data_mem_pkt_offset  = { 1'b1, 1'b1, 1'b0 } - data_mem_pkt_i[136:134];
  assign \data_mem_lines_7_.data_mem_pkt_offset  = { 1'b1, 1'b1, 1'b1 } - data_mem_pkt_i[136:134];
  assign { N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374 } = atomic_reg_data + atomic_mem_data;
  assign data_o = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                  (N173)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                  (N171)? final_data_tv : 1'b0;
  assign N0 = N169;
  assign atomic_reg_data = (N1)? { amo64_reg_in, amo32_reg_in } : 
                           (N175)? { amo32_reg_in, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = N174;
  assign atomic_mem_data = (N2)? final_data_tv : 
                           (N177)? { final_data_tv[31:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2 = N176;
  assign { N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440 } = (N3)? atomic_reg_data : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N439)? atomic_mem_data : 1'b0;
  assign N3 = N438;
  assign { N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506 } = (N4)? atomic_reg_data : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N505)? atomic_mem_data : 1'b0;
  assign N4 = N504;
  assign { N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572 } = (N5)? atomic_reg_data : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N571)? atomic_mem_data : 1'b0;
  assign N5 = N570;
  assign { N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638 } = (N6)? atomic_reg_data : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N637)? atomic_mem_data : 1'b0;
  assign N6 = N636;
  assign { N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702 } = (N7)? { N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N8)? { N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N9)? { N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N10)? { N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N11)? { N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N12)? { N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N13)? { N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N14)? { N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N15)? atomic_reg_data : 1'b0;
  assign N7 = N803;
  assign N8 = N805;
  assign N9 = N801;
  assign N10 = N799;
  assign N11 = N809;
  assign N12 = N811;
  assign N13 = N813;
  assign N14 = N815;
  assign N15 = N181;
  assign atomic_alu_result = (N16)? { N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702 } : 
                             (N17)? atomic_reg_data : 1'b0;
  assign N16 = N178;
  assign N17 = N179;
  assign atomic_result = (N18)? atomic_alu_result : 
                         (N845)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, atomic_alu_result[63:32] } : 1'b0;
  assign N18 = N771;
  assign \wbuf_in_2_.slice_data  = (N19)? atomic_result[31:0] : 
                                   (N767)? amo32_reg_in : 1'b0;
  assign N19 = N766;
  assign \wbuf_in_3_.slice_data  = (N20)? atomic_result : 
                                   (N768)? { amo64_reg_in, amo32_reg_in } : 1'b0;
  assign N20 = N782;
  assign cache_req_o[114:51] = (N21)? { wbuf_entry_in_data__63_, wbuf_entry_in_data__62_, wbuf_entry_in_data__61_, wbuf_entry_in_data__60_, wbuf_entry_in_data__59_, wbuf_entry_in_data__58_, wbuf_entry_in_data__57_, wbuf_entry_in_data__56_, wbuf_entry_in_data__55_, wbuf_entry_in_data__54_, wbuf_entry_in_data__53_, wbuf_entry_in_data__52_, wbuf_entry_in_data__51_, wbuf_entry_in_data__50_, wbuf_entry_in_data__49_, wbuf_entry_in_data__48_, wbuf_entry_in_data__47_, wbuf_entry_in_data__46_, wbuf_entry_in_data__45_, wbuf_entry_in_data__44_, wbuf_entry_in_data__43_, wbuf_entry_in_data__42_, wbuf_entry_in_data__41_, wbuf_entry_in_data__40_, wbuf_entry_in_data__39_, wbuf_entry_in_data__38_, wbuf_entry_in_data__37_, wbuf_entry_in_data__36_, wbuf_entry_in_data__35_, wbuf_entry_in_data__34_, wbuf_entry_in_data__33_, wbuf_entry_in_data__32_, wbuf_entry_in_data__31_, wbuf_entry_in_data__30_, wbuf_entry_in_data__29_, wbuf_entry_in_data__28_, wbuf_entry_in_data__27_, wbuf_entry_in_data__26_, wbuf_entry_in_data__25_, wbuf_entry_in_data__24_, wbuf_entry_in_data__23_, wbuf_entry_in_data__22_, wbuf_entry_in_data__21_, wbuf_entry_in_data__20_, wbuf_entry_in_data__19_, wbuf_entry_in_data__18_, wbuf_entry_in_data__17_, wbuf_entry_in_data__16_, wbuf_entry_in_data__15_, wbuf_entry_in_data__14_, wbuf_entry_in_data__13_, wbuf_entry_in_data__12_, wbuf_entry_in_data__11_, wbuf_entry_in_data__10_, wbuf_entry_in_data__9_, wbuf_entry_in_data__8_, wbuf_entry_in_data__7_, wbuf_entry_in_data__6_, wbuf_entry_in_data__5_, wbuf_entry_in_data__4_, wbuf_entry_in_data__3_, wbuf_entry_in_data__2_, wbuf_entry_in_data__1_, wbuf_entry_in_data__0_ } : 
                               (N22)? { amo64_reg_in, amo32_reg_in } : 1'b0;
  assign N21 = nonblocking_req;
  assign N22 = N1439;
  assign cache_req_o[48] = (N23)? 1'b0 : 
                           (N841)? 1'b0 : 
                           (N844)? 1'b1 : 
                           (N847)? 1'b0 : 
                           (N850)? 1'b1 : 
                           (N778)? 1'b0 : 
                           (N24)? 1'b0 : 1'b0;
  assign N23 = N769;
  assign N24 = 1'b0;
  assign cache_req_o[49] = (N23)? 1'b1 : 
                           (N841)? 1'b1 : 
                           (N844)? 1'b1 : 
                           (N847)? 1'b1 : 
                           (N779)? 1'b0 : 
                           (N24)? 1'b0 : 
                           (N24)? 1'b0 : 1'b0;
  assign cache_req_o[50] = (N23)? 1'b1 : 
                           (N841)? 1'b1 : 
                           (N780)? 1'b0 : 
                           (N24)? 1'b0 : 
                           (N24)? 1'b0 : 
                           (N24)? 1'b0 : 
                           (N24)? 1'b0 : 1'b0;
  assign { N824, N823, N822, N821 } = (N25)? { 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                      (N26)? { 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                      (N27)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                      (N10)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                      (N9)? { 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                      (N7)? { 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                      (N8)? { 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                      (N11)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                      (N12)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                                      (N13)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                                      (N14)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                      (N28)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N25 = N787;
  assign N26 = N791;
  assign N27 = N794;
  assign N28 = N820;
  assign cache_req_o[3:0] = (N20)? { N824, N823, N822, N821 } : 
                            (N29)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N29 = N781;
  assign cache_req_o[5:4] = (N30)? { 1'b0, 1'b1 } : 
                            (N852)? { 1'b1, 1'b1 } : 
                            (N855)? { 1'b0, 1'b0 } : 
                            (N858)? { 1'b1, 1'b1 } : 
                            (N861)? { 1'b1, 1'b0 } : 
                            (N864)? { 1'b0, 1'b0 } : 
                            (N867)? { 1'b0, 1'b1 } : 
                            (N870)? { 1'b0, 1'b0 } : 
                            (N873)? { 1'b0, 1'b1 } : 
                            (N876)? { 1'b0, 1'b0 } : 
                            (N879)? { 1'b1, 1'b1 } : 
                            (N837)? { 1'b1, 1'b0 } : 1'b0;
  assign N30 = N825;
  assign cache_req_o[6] = (N30)? 1'b1 : 
                          (N852)? 1'b0 : 
                          (N855)? 1'b1 : 
                          (N858)? 1'b1 : 
                          (N861)? 1'b1 : 
                          (N864)? 1'b0 : 
                          (N867)? 1'b0 : 
                          (N870)? 1'b0 : 
                          (N873)? 1'b1 : 
                          (N876)? 1'b1 : 
                          (N838)? 1'b0 : 
                          (N24)? 1'b0 : 1'b0;
  assign cache_req_o[7] = (N30)? 1'b1 : 
                          (N852)? 1'b1 : 
                          (N855)? 1'b1 : 
                          (N858)? 1'b0 : 
                          (N861)? 1'b0 : 
                          (N864)? 1'b1 : 
                          (N839)? 1'b0 : 
                          (N24)? 1'b0 : 
                          (N24)? 1'b0 : 
                          (N24)? 1'b0 : 
                          (N24)? 1'b0 : 
                          (N24)? 1'b0 : 1'b0;
  assign lru_way_li = (N31)? metadata_invalid_way : 
                      (N32)? lru_encode : 1'b0;
  assign N31 = metadata_invalid_exist;
  assign N32 = N880;
  assign cache_req_metadata_o[3:1] = (N33)? metadata_hit_index_r : 
                                     (N34)? lru_way_li : 1'b0;
  assign N33 = metadata_hit_r;
  assign N34 = N881;
  assign tag_mem_addr_li = (N35)? cache_req_o[19:14] : 
                           (N900)? dcache_pkt_i[11:6] : 
                           (N898)? tag_mem_pkt_i[34:29] : 1'b0;
  assign N35 = tag_mem_fast_write;
  assign tag_mem_data_li[22:0] = (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N36)? tag_mem_pkt_i[25:3] : 
                                 (N37)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N38)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N39)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N36 = N905;
  assign N37 = N910;
  assign N38 = N916;
  assign N39 = N922;
  assign tag_mem_mask_li[22:0] = (N35)? { N1242, N1242, N1242, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N36)? { tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0] } : 
                                 (N37)? { tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N38)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N39)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[45:23] = (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N40)? tag_mem_pkt_i[25:3] : 
                                  (N41)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N42)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N43)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N40 = N927;
  assign N41 = N932;
  assign N42 = N938;
  assign N43 = N944;
  assign tag_mem_mask_li[45:23] = (N35)? { N1239, N1239, N1239, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N40)? { tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1] } : 
                                  (N41)? { tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N42)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N43)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[68:46] = (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N44)? tag_mem_pkt_i[25:3] : 
                                  (N45)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N46)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N47)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N44 = N949;
  assign N45 = N954;
  assign N46 = N960;
  assign N47 = N966;
  assign tag_mem_mask_li[68:46] = (N35)? { N1235, N1235, N1235, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N44)? { tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2] } : 
                                  (N45)? { tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N46)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N47)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[91:69] = (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N48)? tag_mem_pkt_i[25:3] : 
                                  (N49)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N50)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N51)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N48 = N971;
  assign N49 = N976;
  assign N50 = N982;
  assign N51 = N988;
  assign tag_mem_mask_li[91:69] = (N35)? { N1231, N1231, N1231, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N48)? { tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3] } : 
                                  (N49)? { tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N50)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N51)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[114:92] = (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N52)? tag_mem_pkt_i[25:3] : 
                                   (N53)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N54)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N55)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N52 = N993;
  assign N53 = N998;
  assign N54 = N1004;
  assign N55 = N1010;
  assign tag_mem_mask_li[114:92] = (N35)? { N1226, N1226, N1226, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N52)? { tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4] } : 
                                   (N53)? { tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N54)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N55)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[137:115] = (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N56)? tag_mem_pkt_i[25:3] : 
                                    (N57)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N58)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N59)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N56 = N1015;
  assign N57 = N1020;
  assign N58 = N1026;
  assign N59 = N1032;
  assign tag_mem_mask_li[137:115] = (N35)? { N1222, N1222, N1222, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N56)? { tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5] } : 
                                    (N57)? { tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N58)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N59)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[160:138] = (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N60)? tag_mem_pkt_i[25:3] : 
                                    (N61)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N62)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N63)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N60 = N1037;
  assign N61 = N1042;
  assign N62 = N1048;
  assign N63 = N1054;
  assign tag_mem_mask_li[160:138] = (N35)? { N1217, N1217, N1217, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N60)? { tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6] } : 
                                    (N61)? { tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N62)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N63)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[183:161] = (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N64)? tag_mem_pkt_i[25:3] : 
                                    (N65)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N66)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N67)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N64 = N1059;
  assign N65 = N1064;
  assign N66 = N1070;
  assign N67 = N1076;
  assign tag_mem_mask_li[183:161] = (N35)? { N1212, N1212, N1212, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N64)? { tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7] } : 
                                    (N65)? { tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N66)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N67)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign data_mem_mask_li[7:0] = (N68)? wbuf_data_mem_mask : 
                                 (N1092)? { data_mem_write_bank_mask[0:0], data_mem_write_bank_mask[0:0], data_mem_write_bank_mask[0:0], data_mem_write_bank_mask[0:0], data_mem_write_bank_mask[0:0], data_mem_write_bank_mask[0:0], data_mem_write_bank_mask[0:0], data_mem_write_bank_mask[0:0] } : 1'b0;
  assign N68 = data_mem_fast_write[0];
  assign data_mem_addr_li[8:0] = (N68)? { wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_ } : 
                                 (N1095)? dcache_pkt_i[11:3] : 
                                 (N1094)? { data_mem_pkt_i[142:137], \data_mem_lines_0_.data_mem_pkt_offset  } : 1'b0;
  assign data_mem_data_li[63:0] = (N68)? { wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_ } : 
                                  (N1092)? data_mem_pkt_fill_data_li[63:0] : 1'b0;
  assign data_mem_mask_li[15:8] = (N69)? wbuf_data_mem_mask : 
                                  (N1096)? { data_mem_write_bank_mask[1:1], data_mem_write_bank_mask[1:1], data_mem_write_bank_mask[1:1], data_mem_write_bank_mask[1:1], data_mem_write_bank_mask[1:1], data_mem_write_bank_mask[1:1], data_mem_write_bank_mask[1:1], data_mem_write_bank_mask[1:1] } : 1'b0;
  assign N69 = data_mem_fast_write[1];
  assign data_mem_addr_li[17:9] = (N69)? { wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_ } : 
                                  (N1099)? dcache_pkt_i[11:3] : 
                                  (N1098)? { data_mem_pkt_i[142:137], \data_mem_lines_1_.data_mem_pkt_offset  } : 1'b0;
  assign data_mem_data_li[127:64] = (N69)? { wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_ } : 
                                    (N1096)? data_mem_pkt_fill_data_li[127:64] : 1'b0;
  assign data_mem_mask_li[23:16] = (N70)? wbuf_data_mem_mask : 
                                   (N1100)? { data_mem_write_bank_mask[2:2], data_mem_write_bank_mask[2:2], data_mem_write_bank_mask[2:2], data_mem_write_bank_mask[2:2], data_mem_write_bank_mask[2:2], data_mem_write_bank_mask[2:2], data_mem_write_bank_mask[2:2], data_mem_write_bank_mask[2:2] } : 1'b0;
  assign N70 = data_mem_fast_write[2];
  assign data_mem_addr_li[26:18] = (N70)? { wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_ } : 
                                   (N1103)? dcache_pkt_i[11:3] : 
                                   (N1102)? { data_mem_pkt_i[142:137], \data_mem_lines_2_.data_mem_pkt_offset  } : 1'b0;
  assign data_mem_data_li[191:128] = (N70)? { wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_ } : 
                                     (N1100)? data_mem_pkt_fill_data_li[63:0] : 1'b0;
  assign data_mem_mask_li[31:24] = (N71)? wbuf_data_mem_mask : 
                                   (N1104)? { data_mem_write_bank_mask[3:3], data_mem_write_bank_mask[3:3], data_mem_write_bank_mask[3:3], data_mem_write_bank_mask[3:3], data_mem_write_bank_mask[3:3], data_mem_write_bank_mask[3:3], data_mem_write_bank_mask[3:3], data_mem_write_bank_mask[3:3] } : 1'b0;
  assign N71 = data_mem_fast_write[3];
  assign data_mem_addr_li[35:27] = (N71)? { wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_ } : 
                                   (N1107)? dcache_pkt_i[11:3] : 
                                   (N1106)? { data_mem_pkt_i[142:137], \data_mem_lines_3_.data_mem_pkt_offset  } : 1'b0;
  assign data_mem_data_li[255:192] = (N71)? { wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_ } : 
                                     (N1104)? data_mem_pkt_fill_data_li[127:64] : 1'b0;
  assign data_mem_mask_li[39:32] = (N72)? wbuf_data_mem_mask : 
                                   (N1108)? { data_mem_write_bank_mask[4:4], data_mem_write_bank_mask[4:4], data_mem_write_bank_mask[4:4], data_mem_write_bank_mask[4:4], data_mem_write_bank_mask[4:4], data_mem_write_bank_mask[4:4], data_mem_write_bank_mask[4:4], data_mem_write_bank_mask[4:4] } : 1'b0;
  assign N72 = data_mem_fast_write[4];
  assign data_mem_addr_li[44:36] = (N72)? { wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_ } : 
                                   (N1111)? dcache_pkt_i[11:3] : 
                                   (N1110)? { data_mem_pkt_i[142:137], \data_mem_lines_4_.data_mem_pkt_offset  } : 1'b0;
  assign data_mem_data_li[319:256] = (N72)? { wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_ } : 
                                     (N1108)? data_mem_pkt_fill_data_li[63:0] : 1'b0;
  assign data_mem_mask_li[47:40] = (N73)? wbuf_data_mem_mask : 
                                   (N1112)? { data_mem_write_bank_mask[5:5], data_mem_write_bank_mask[5:5], data_mem_write_bank_mask[5:5], data_mem_write_bank_mask[5:5], data_mem_write_bank_mask[5:5], data_mem_write_bank_mask[5:5], data_mem_write_bank_mask[5:5], data_mem_write_bank_mask[5:5] } : 1'b0;
  assign N73 = data_mem_fast_write[5];
  assign data_mem_addr_li[53:45] = (N73)? { wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_ } : 
                                   (N1115)? dcache_pkt_i[11:3] : 
                                   (N1114)? { data_mem_pkt_i[142:137], \data_mem_lines_5_.data_mem_pkt_offset  } : 1'b0;
  assign data_mem_data_li[383:320] = (N73)? { wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_ } : 
                                     (N1112)? data_mem_pkt_fill_data_li[127:64] : 1'b0;
  assign data_mem_mask_li[55:48] = (N74)? wbuf_data_mem_mask : 
                                   (N1116)? { data_mem_write_bank_mask[6:6], data_mem_write_bank_mask[6:6], data_mem_write_bank_mask[6:6], data_mem_write_bank_mask[6:6], data_mem_write_bank_mask[6:6], data_mem_write_bank_mask[6:6], data_mem_write_bank_mask[6:6], data_mem_write_bank_mask[6:6] } : 1'b0;
  assign N74 = data_mem_fast_write[6];
  assign data_mem_addr_li[62:54] = (N74)? { wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_ } : 
                                   (N1119)? dcache_pkt_i[11:3] : 
                                   (N1118)? { data_mem_pkt_i[142:137], \data_mem_lines_6_.data_mem_pkt_offset  } : 1'b0;
  assign data_mem_data_li[447:384] = (N74)? { wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_ } : 
                                     (N1116)? data_mem_pkt_fill_data_li[63:0] : 1'b0;
  assign data_mem_mask_li[63:56] = (N75)? wbuf_data_mem_mask : 
                                   (N1120)? { data_mem_write_bank_mask[7:7], data_mem_write_bank_mask[7:7], data_mem_write_bank_mask[7:7], data_mem_write_bank_mask[7:7], data_mem_write_bank_mask[7:7], data_mem_write_bank_mask[7:7], data_mem_write_bank_mask[7:7], data_mem_write_bank_mask[7:7] } : 1'b0;
  assign N75 = data_mem_fast_write[7];
  assign data_mem_addr_li[71:63] = (N75)? { wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_ } : 
                                   (N1123)? dcache_pkt_i[11:3] : 
                                   (N1122)? { data_mem_pkt_i[142:137], \data_mem_lines_7_.data_mem_pkt_offset  } : 1'b0;
  assign data_mem_data_li[511:448] = (N75)? { wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_ } : 
                                     (N1120)? data_mem_pkt_fill_data_li[127:64] : 1'b0;
  assign stat_mem_addr_li = (N76)? cache_req_o[19:14] : 
                            (N1125)? stat_mem_pkt_i[10:5] : 1'b0;
  assign N76 = N1124;
  assign { N1130, N1129, N1128 } = (N77)? store_hit_way_tv : 
                                   (N1127)? load_hit_way_tv : 1'b0;
  assign N77 = N1126;
  assign lru_decode_way_li = (N78)? { N1130, N1129, N1128 } : 
                             (N79)? stat_mem_pkt_i[4:2] : 1'b0;
  assign N78 = v_tv_r;
  assign N79 = N1513;
  assign \tdm.dirty_mask_way_li  = (N78)? store_hit_way_tv : 
                                   (N79)? stat_mem_pkt_i[4:2] : 1'b0;
  assign { N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136 } = (N80)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                      (N81)? dirty_mask_lo : 1'b0;
  assign N80 = N1134;
  assign N81 = N1135;
  assign stat_mem_data_li[0] = ~N1132;
  assign stat_mem_data_li[1] = ~N1132;
  assign stat_mem_data_li[2] = ~N1132;
  assign stat_mem_data_li[3] = ~N1132;
  assign stat_mem_data_li[4] = ~N1132;
  assign stat_mem_data_li[5] = ~N1132;
  assign stat_mem_data_li[6] = ~N1132;
  assign stat_mem_data_li[7] = ~N1132;
  assign stat_mem_data_li[14:8] = (N82)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N1133)? lru_decode_data_lo : 1'b0;
  assign N82 = N1132;
  assign stat_mem_mask_li = (N82)? { N1134, N1134, N1134, N1134, N1134, N1134, N1134, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136 } : 
                            (N1133)? { lru_decode_mask_lo, dirty_mask_lo } : 1'b0;
  assign N1154 = ~N1155;
  assign state_n = (N83)? { 1'b0, 1'b0 } : 
                   (N1157)? { N1155, N1154 } : 
                   (N1160)? { 1'b1, 1'b0 } : 
                   (N1153)? state_r : 1'b0;
  assign N83 = N1148;
  assign \hum.fill_bank_mask_n  = (N84)? { N1162, N1163, N1164, N1165, N1166, N1167, N1168, N1169 } : 
                                  (N85)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N84 = \hum.fill_v ;
  assign N85 = N1161;
  assign \hum.fill_hit_n  = (N84)? { N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170 } : 
                            (N85)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N1330 = N86 & decode_tv_r_amo_subop__0_;
  assign N86 = ~decode_tv_r_amo_subop__1_;
  assign N1331 = N1330 | decode_tv_r_amo_subop__1_;
  assign N1332 = N87 & N1331;
  assign N87 = ~decode_tv_r_amo_subop__2_;
  assign N1333 = N1332 | decode_tv_r_amo_subop__2_;
  assign N1334 = ~decode_tv_r_amo_subop__2_;
  assign N1335 = N88 & N1333;
  assign N88 = ~decode_tv_r_amo_subop__3_;
  assign N1336 = decode_tv_r_amo_subop__3_ & N1334;
  assign N178 = N1335 | N1336;
  assign flush_tv = N1339 | fill_hazard;
  assign N1339 = N1338 | nonblocking_hazard;
  assign N1338 = N1337 | blocking_hazard;
  assign N1337 = flush_i | tag_mem_fast_write;
  assign flush_tl = flush_tv | data_mem_write_hazard;
  assign critical_recv = N1345 & N1347;
  assign N1345 = N1342 & N1344;
  assign N1342 = cache_req_critical_i & N1341;
  assign N1341 = N1340 | stat_mem_pkt_yumi_o;
  assign N1340 = ~stat_mem_pkt_v_i;
  assign N1344 = N1343 | tag_mem_pkt_yumi_o;
  assign N1343 = ~tag_mem_pkt_v_i;
  assign N1347 = N1346 | data_mem_pkt_yumi_o;
  assign N1346 = ~data_mem_pkt_v_i;
  assign complete_recv = N1353 & N1355;
  assign N1353 = N1350 & N1352;
  assign N1350 = cache_req_last_i & N1349;
  assign N1349 = N1348 | stat_mem_pkt_yumi_o;
  assign N1348 = ~stat_mem_pkt_v_i;
  assign N1352 = N1351 | tag_mem_pkt_yumi_o;
  assign N1351 = ~tag_mem_pkt_v_i;
  assign N1355 = N1354 | data_mem_pkt_yumi_o;
  assign N1354 = ~data_mem_pkt_v_i;
  assign safe_tl_we = v_i & N1356;
  assign N1356 = ~busy_o;
  assign tl_we = safe_tl_we & N1357;
  assign N1357 = ~flush_tl;
  assign \tag_comp_tl_0_.tag_match_tl  = N1366 & N89;
  assign N1366 = ptag_v_i & N1365;
  assign N1365 = ~N1364;
  assign N1364 = N1363 | ptag_i[20];
  assign N1363 = N1362 | ptag_i[21];
  assign N1362 = N1361 | ptag_i[22];
  assign N1361 = N1360 | ptag_i[23];
  assign N1360 = N1359 | ptag_i[24];
  assign N1359 = N1358 | ptag_i[25];
  assign N1358 = ptag_i[27] | ptag_i[26];
  assign load_hit_tl[0] = \tag_comp_tl_0_.tag_match_tl  & N1310;
  assign store_hit_tl[0] = \tag_comp_tl_0_.tag_match_tl  & N98;
  assign \tag_comp_tl_1_.tag_match_tl  = N1375 & N99;
  assign N1375 = ptag_v_i & N1374;
  assign N1374 = ~N1373;
  assign N1373 = N1372 | ptag_i[20];
  assign N1372 = N1371 | ptag_i[21];
  assign N1371 = N1370 | ptag_i[22];
  assign N1370 = N1369 | ptag_i[23];
  assign N1369 = N1368 | ptag_i[24];
  assign N1368 = N1367 | ptag_i[25];
  assign N1367 = ptag_i[27] | ptag_i[26];
  assign load_hit_tl[1] = \tag_comp_tl_1_.tag_match_tl  & N1308;
  assign store_hit_tl[1] = \tag_comp_tl_1_.tag_match_tl  & N108;
  assign \tag_comp_tl_2_.tag_match_tl  = N1384 & N109;
  assign N1384 = ptag_v_i & N1383;
  assign N1383 = ~N1382;
  assign N1382 = N1381 | ptag_i[20];
  assign N1381 = N1380 | ptag_i[21];
  assign N1380 = N1379 | ptag_i[22];
  assign N1379 = N1378 | ptag_i[23];
  assign N1378 = N1377 | ptag_i[24];
  assign N1377 = N1376 | ptag_i[25];
  assign N1376 = ptag_i[27] | ptag_i[26];
  assign load_hit_tl[2] = \tag_comp_tl_2_.tag_match_tl  & N1306;
  assign store_hit_tl[2] = \tag_comp_tl_2_.tag_match_tl  & N118;
  assign \tag_comp_tl_3_.tag_match_tl  = N1393 & N119;
  assign N1393 = ptag_v_i & N1392;
  assign N1392 = ~N1391;
  assign N1391 = N1390 | ptag_i[20];
  assign N1390 = N1389 | ptag_i[21];
  assign N1389 = N1388 | ptag_i[22];
  assign N1388 = N1387 | ptag_i[23];
  assign N1387 = N1386 | ptag_i[24];
  assign N1386 = N1385 | ptag_i[25];
  assign N1385 = ptag_i[27] | ptag_i[26];
  assign load_hit_tl[3] = \tag_comp_tl_3_.tag_match_tl  & N1304;
  assign store_hit_tl[3] = \tag_comp_tl_3_.tag_match_tl  & N128;
  assign \tag_comp_tl_4_.tag_match_tl  = N1402 & N129;
  assign N1402 = ptag_v_i & N1401;
  assign N1401 = ~N1400;
  assign N1400 = N1399 | ptag_i[20];
  assign N1399 = N1398 | ptag_i[21];
  assign N1398 = N1397 | ptag_i[22];
  assign N1397 = N1396 | ptag_i[23];
  assign N1396 = N1395 | ptag_i[24];
  assign N1395 = N1394 | ptag_i[25];
  assign N1394 = ptag_i[27] | ptag_i[26];
  assign load_hit_tl[4] = \tag_comp_tl_4_.tag_match_tl  & N1302;
  assign store_hit_tl[4] = \tag_comp_tl_4_.tag_match_tl  & N138;
  assign \tag_comp_tl_5_.tag_match_tl  = N1411 & N139;
  assign N1411 = ptag_v_i & N1410;
  assign N1410 = ~N1409;
  assign N1409 = N1408 | ptag_i[20];
  assign N1408 = N1407 | ptag_i[21];
  assign N1407 = N1406 | ptag_i[22];
  assign N1406 = N1405 | ptag_i[23];
  assign N1405 = N1404 | ptag_i[24];
  assign N1404 = N1403 | ptag_i[25];
  assign N1403 = ptag_i[27] | ptag_i[26];
  assign load_hit_tl[5] = \tag_comp_tl_5_.tag_match_tl  & N1300;
  assign store_hit_tl[5] = \tag_comp_tl_5_.tag_match_tl  & N148;
  assign \tag_comp_tl_6_.tag_match_tl  = N1420 & N149;
  assign N1420 = ptag_v_i & N1419;
  assign N1419 = ~N1418;
  assign N1418 = N1417 | ptag_i[20];
  assign N1417 = N1416 | ptag_i[21];
  assign N1416 = N1415 | ptag_i[22];
  assign N1415 = N1414 | ptag_i[23];
  assign N1414 = N1413 | ptag_i[24];
  assign N1413 = N1412 | ptag_i[25];
  assign N1412 = ptag_i[27] | ptag_i[26];
  assign load_hit_tl[6] = \tag_comp_tl_6_.tag_match_tl  & N1298;
  assign store_hit_tl[6] = \tag_comp_tl_6_.tag_match_tl  & N158;
  assign \tag_comp_tl_7_.tag_match_tl  = N1429 & N159;
  assign N1429 = ptag_v_i & N1428;
  assign N1428 = ~N1427;
  assign N1427 = N1426 | ptag_i[20];
  assign N1426 = N1425 | ptag_i[21];
  assign N1425 = N1424 | ptag_i[22];
  assign N1424 = N1423 | ptag_i[23];
  assign N1423 = N1422 | ptag_i[24];
  assign N1422 = N1421 | ptag_i[25];
  assign N1421 = ptag_i[27] | ptag_i[26];
  assign load_hit_tl[7] = \tag_comp_tl_7_.tag_match_tl  & N1296;
  assign store_hit_tl[7] = \tag_comp_tl_7_.tag_match_tl  & N168;
  assign uncached_tl = N1430 & N1431;
  assign N1430 = ~decode_tl_r[23];
  assign N1431 = decode_tl_r[17] | ptag_uncached_i;
  assign safe_tv_we = v_tl_r & N1432;
  assign N1432 = ptag_v_i | decode_tl_r[23];
  assign tv_we = safe_tv_we & N1433;
  assign N1433 = ~flush_tv;
  assign _2_net_ = tv_we | critical_recv;
  assign store_miss_tv = N1438 & N1439;
  assign N1438 = N1436 & N1437;
  assign N1436 = N1434 & N1435;
  assign N1434 = decode_tv_r_store_op_ | decode_tv_r_lr_op_;
  assign N1435 = ~store_hit_tv;
  assign N1437 = ~sc_fail_tv;
  assign N1439 = ~nonblocking_req;
  assign load_miss_tv = N1442 & N1439;
  assign N1442 = N1441 & N1437;
  assign N1441 = decode_tv_r_load_op_ & N1440;
  assign N1440 = ~cache_req_o[115];
  assign nonblocking_miss_tv = nonblocking_req & N1443;
  assign N1443 = ~cache_req_yumi_i;
  assign engine_miss_tv = cache_req_v_o & N1444;
  assign N1444 = ~cache_req_yumi_i;
  assign any_miss_tv = N1445 | engine_miss_tv;
  assign N1445 = blocking_miss_tv | nonblocking_miss_tv;
  assign v_o = v_tv_r & N1446;
  assign N1446 = ~any_miss_tv;
  assign N169 = sc_success_tv;
  assign N170 = sc_fail_tv | N169;
  assign N171 = ~N170;
  assign N172 = ~N169;
  assign N173 = sc_fail_tv & N172;
  assign unsigned_o = ~decode_tv_r_signed_op_;
  assign wbuf_v_li = N1451 & N1446;
  assign N1451 = N1449 & N1450;
  assign N1449 = N1448 & N1437;
  assign N1448 = N1447 & store_hit_tv;
  assign N1447 = v_tv_r & decode_tv_r_store_op_;
  assign N1450 = ~uncached_tv_r;
  assign N174 = decode_tv_r_double_op_;
  assign N175 = ~N174;
  assign N176 = decode_tv_r_double_op_;
  assign N177 = ~N176;
  assign N179 = ~N178;
  assign N180 = N178;
  assign N181 = N816 | N817;
  assign N182 = atomic_reg_data[63] & atomic_mem_data[63];
  assign N183 = atomic_reg_data[62] & atomic_mem_data[62];
  assign N184 = atomic_reg_data[61] & atomic_mem_data[61];
  assign N185 = atomic_reg_data[60] & atomic_mem_data[60];
  assign N186 = atomic_reg_data[59] & atomic_mem_data[59];
  assign N187 = atomic_reg_data[58] & atomic_mem_data[58];
  assign N188 = atomic_reg_data[57] & atomic_mem_data[57];
  assign N189 = atomic_reg_data[56] & atomic_mem_data[56];
  assign N190 = atomic_reg_data[55] & atomic_mem_data[55];
  assign N191 = atomic_reg_data[54] & atomic_mem_data[54];
  assign N192 = atomic_reg_data[53] & atomic_mem_data[53];
  assign N193 = atomic_reg_data[52] & atomic_mem_data[52];
  assign N194 = atomic_reg_data[51] & atomic_mem_data[51];
  assign N195 = atomic_reg_data[50] & atomic_mem_data[50];
  assign N196 = atomic_reg_data[49] & atomic_mem_data[49];
  assign N197 = atomic_reg_data[48] & atomic_mem_data[48];
  assign N198 = atomic_reg_data[47] & atomic_mem_data[47];
  assign N199 = atomic_reg_data[46] & atomic_mem_data[46];
  assign N200 = atomic_reg_data[45] & atomic_mem_data[45];
  assign N201 = atomic_reg_data[44] & atomic_mem_data[44];
  assign N202 = atomic_reg_data[43] & atomic_mem_data[43];
  assign N203 = atomic_reg_data[42] & atomic_mem_data[42];
  assign N204 = atomic_reg_data[41] & atomic_mem_data[41];
  assign N205 = atomic_reg_data[40] & atomic_mem_data[40];
  assign N206 = atomic_reg_data[39] & atomic_mem_data[39];
  assign N207 = atomic_reg_data[38] & atomic_mem_data[38];
  assign N208 = atomic_reg_data[37] & atomic_mem_data[37];
  assign N209 = atomic_reg_data[36] & atomic_mem_data[36];
  assign N210 = atomic_reg_data[35] & atomic_mem_data[35];
  assign N211 = atomic_reg_data[34] & atomic_mem_data[34];
  assign N212 = atomic_reg_data[33] & atomic_mem_data[33];
  assign N213 = atomic_reg_data[32] & atomic_mem_data[32];
  assign N214 = atomic_reg_data[31] & atomic_mem_data[31];
  assign N215 = atomic_reg_data[30] & atomic_mem_data[30];
  assign N216 = atomic_reg_data[29] & atomic_mem_data[29];
  assign N217 = atomic_reg_data[28] & atomic_mem_data[28];
  assign N218 = atomic_reg_data[27] & atomic_mem_data[27];
  assign N219 = atomic_reg_data[26] & atomic_mem_data[26];
  assign N220 = atomic_reg_data[25] & atomic_mem_data[25];
  assign N221 = atomic_reg_data[24] & atomic_mem_data[24];
  assign N222 = atomic_reg_data[23] & atomic_mem_data[23];
  assign N223 = atomic_reg_data[22] & atomic_mem_data[22];
  assign N224 = atomic_reg_data[21] & atomic_mem_data[21];
  assign N225 = atomic_reg_data[20] & atomic_mem_data[20];
  assign N226 = atomic_reg_data[19] & atomic_mem_data[19];
  assign N227 = atomic_reg_data[18] & atomic_mem_data[18];
  assign N228 = atomic_reg_data[17] & atomic_mem_data[17];
  assign N229 = atomic_reg_data[16] & atomic_mem_data[16];
  assign N230 = atomic_reg_data[15] & atomic_mem_data[15];
  assign N231 = atomic_reg_data[14] & atomic_mem_data[14];
  assign N232 = atomic_reg_data[13] & atomic_mem_data[13];
  assign N233 = atomic_reg_data[12] & atomic_mem_data[12];
  assign N234 = atomic_reg_data[11] & atomic_mem_data[11];
  assign N235 = atomic_reg_data[10] & atomic_mem_data[10];
  assign N236 = atomic_reg_data[9] & atomic_mem_data[9];
  assign N237 = atomic_reg_data[8] & atomic_mem_data[8];
  assign N238 = atomic_reg_data[7] & atomic_mem_data[7];
  assign N239 = atomic_reg_data[6] & atomic_mem_data[6];
  assign N240 = atomic_reg_data[5] & atomic_mem_data[5];
  assign N241 = atomic_reg_data[4] & atomic_mem_data[4];
  assign N242 = atomic_reg_data[3] & atomic_mem_data[3];
  assign N243 = atomic_reg_data[2] & atomic_mem_data[2];
  assign N244 = atomic_reg_data[1] & atomic_mem_data[1];
  assign N245 = atomic_reg_data[0] & atomic_mem_data[0];
  assign N246 = atomic_reg_data[63] | atomic_mem_data[63];
  assign N247 = atomic_reg_data[62] | atomic_mem_data[62];
  assign N248 = atomic_reg_data[61] | atomic_mem_data[61];
  assign N249 = atomic_reg_data[60] | atomic_mem_data[60];
  assign N250 = atomic_reg_data[59] | atomic_mem_data[59];
  assign N251 = atomic_reg_data[58] | atomic_mem_data[58];
  assign N252 = atomic_reg_data[57] | atomic_mem_data[57];
  assign N253 = atomic_reg_data[56] | atomic_mem_data[56];
  assign N254 = atomic_reg_data[55] | atomic_mem_data[55];
  assign N255 = atomic_reg_data[54] | atomic_mem_data[54];
  assign N256 = atomic_reg_data[53] | atomic_mem_data[53];
  assign N257 = atomic_reg_data[52] | atomic_mem_data[52];
  assign N258 = atomic_reg_data[51] | atomic_mem_data[51];
  assign N259 = atomic_reg_data[50] | atomic_mem_data[50];
  assign N260 = atomic_reg_data[49] | atomic_mem_data[49];
  assign N261 = atomic_reg_data[48] | atomic_mem_data[48];
  assign N262 = atomic_reg_data[47] | atomic_mem_data[47];
  assign N263 = atomic_reg_data[46] | atomic_mem_data[46];
  assign N264 = atomic_reg_data[45] | atomic_mem_data[45];
  assign N265 = atomic_reg_data[44] | atomic_mem_data[44];
  assign N266 = atomic_reg_data[43] | atomic_mem_data[43];
  assign N267 = atomic_reg_data[42] | atomic_mem_data[42];
  assign N268 = atomic_reg_data[41] | atomic_mem_data[41];
  assign N269 = atomic_reg_data[40] | atomic_mem_data[40];
  assign N270 = atomic_reg_data[39] | atomic_mem_data[39];
  assign N271 = atomic_reg_data[38] | atomic_mem_data[38];
  assign N272 = atomic_reg_data[37] | atomic_mem_data[37];
  assign N273 = atomic_reg_data[36] | atomic_mem_data[36];
  assign N274 = atomic_reg_data[35] | atomic_mem_data[35];
  assign N275 = atomic_reg_data[34] | atomic_mem_data[34];
  assign N276 = atomic_reg_data[33] | atomic_mem_data[33];
  assign N277 = atomic_reg_data[32] | atomic_mem_data[32];
  assign N278 = atomic_reg_data[31] | atomic_mem_data[31];
  assign N279 = atomic_reg_data[30] | atomic_mem_data[30];
  assign N280 = atomic_reg_data[29] | atomic_mem_data[29];
  assign N281 = atomic_reg_data[28] | atomic_mem_data[28];
  assign N282 = atomic_reg_data[27] | atomic_mem_data[27];
  assign N283 = atomic_reg_data[26] | atomic_mem_data[26];
  assign N284 = atomic_reg_data[25] | atomic_mem_data[25];
  assign N285 = atomic_reg_data[24] | atomic_mem_data[24];
  assign N286 = atomic_reg_data[23] | atomic_mem_data[23];
  assign N287 = atomic_reg_data[22] | atomic_mem_data[22];
  assign N288 = atomic_reg_data[21] | atomic_mem_data[21];
  assign N289 = atomic_reg_data[20] | atomic_mem_data[20];
  assign N290 = atomic_reg_data[19] | atomic_mem_data[19];
  assign N291 = atomic_reg_data[18] | atomic_mem_data[18];
  assign N292 = atomic_reg_data[17] | atomic_mem_data[17];
  assign N293 = atomic_reg_data[16] | atomic_mem_data[16];
  assign N294 = atomic_reg_data[15] | atomic_mem_data[15];
  assign N295 = atomic_reg_data[14] | atomic_mem_data[14];
  assign N296 = atomic_reg_data[13] | atomic_mem_data[13];
  assign N297 = atomic_reg_data[12] | atomic_mem_data[12];
  assign N298 = atomic_reg_data[11] | atomic_mem_data[11];
  assign N299 = atomic_reg_data[10] | atomic_mem_data[10];
  assign N300 = atomic_reg_data[9] | atomic_mem_data[9];
  assign N301 = atomic_reg_data[8] | atomic_mem_data[8];
  assign N302 = atomic_reg_data[7] | atomic_mem_data[7];
  assign N303 = atomic_reg_data[6] | atomic_mem_data[6];
  assign N304 = atomic_reg_data[5] | atomic_mem_data[5];
  assign N305 = atomic_reg_data[4] | atomic_mem_data[4];
  assign N306 = atomic_reg_data[3] | atomic_mem_data[3];
  assign N307 = atomic_reg_data[2] | atomic_mem_data[2];
  assign N308 = atomic_reg_data[1] | atomic_mem_data[1];
  assign N309 = atomic_reg_data[0] | atomic_mem_data[0];
  assign N310 = atomic_reg_data[63] ^ atomic_mem_data[63];
  assign N311 = atomic_reg_data[62] ^ atomic_mem_data[62];
  assign N312 = atomic_reg_data[61] ^ atomic_mem_data[61];
  assign N313 = atomic_reg_data[60] ^ atomic_mem_data[60];
  assign N314 = atomic_reg_data[59] ^ atomic_mem_data[59];
  assign N315 = atomic_reg_data[58] ^ atomic_mem_data[58];
  assign N316 = atomic_reg_data[57] ^ atomic_mem_data[57];
  assign N317 = atomic_reg_data[56] ^ atomic_mem_data[56];
  assign N318 = atomic_reg_data[55] ^ atomic_mem_data[55];
  assign N319 = atomic_reg_data[54] ^ atomic_mem_data[54];
  assign N320 = atomic_reg_data[53] ^ atomic_mem_data[53];
  assign N321 = atomic_reg_data[52] ^ atomic_mem_data[52];
  assign N322 = atomic_reg_data[51] ^ atomic_mem_data[51];
  assign N323 = atomic_reg_data[50] ^ atomic_mem_data[50];
  assign N324 = atomic_reg_data[49] ^ atomic_mem_data[49];
  assign N325 = atomic_reg_data[48] ^ atomic_mem_data[48];
  assign N326 = atomic_reg_data[47] ^ atomic_mem_data[47];
  assign N327 = atomic_reg_data[46] ^ atomic_mem_data[46];
  assign N328 = atomic_reg_data[45] ^ atomic_mem_data[45];
  assign N329 = atomic_reg_data[44] ^ atomic_mem_data[44];
  assign N330 = atomic_reg_data[43] ^ atomic_mem_data[43];
  assign N331 = atomic_reg_data[42] ^ atomic_mem_data[42];
  assign N332 = atomic_reg_data[41] ^ atomic_mem_data[41];
  assign N333 = atomic_reg_data[40] ^ atomic_mem_data[40];
  assign N334 = atomic_reg_data[39] ^ atomic_mem_data[39];
  assign N335 = atomic_reg_data[38] ^ atomic_mem_data[38];
  assign N336 = atomic_reg_data[37] ^ atomic_mem_data[37];
  assign N337 = atomic_reg_data[36] ^ atomic_mem_data[36];
  assign N338 = atomic_reg_data[35] ^ atomic_mem_data[35];
  assign N339 = atomic_reg_data[34] ^ atomic_mem_data[34];
  assign N340 = atomic_reg_data[33] ^ atomic_mem_data[33];
  assign N341 = atomic_reg_data[32] ^ atomic_mem_data[32];
  assign N342 = atomic_reg_data[31] ^ atomic_mem_data[31];
  assign N343 = atomic_reg_data[30] ^ atomic_mem_data[30];
  assign N344 = atomic_reg_data[29] ^ atomic_mem_data[29];
  assign N345 = atomic_reg_data[28] ^ atomic_mem_data[28];
  assign N346 = atomic_reg_data[27] ^ atomic_mem_data[27];
  assign N347 = atomic_reg_data[26] ^ atomic_mem_data[26];
  assign N348 = atomic_reg_data[25] ^ atomic_mem_data[25];
  assign N349 = atomic_reg_data[24] ^ atomic_mem_data[24];
  assign N350 = atomic_reg_data[23] ^ atomic_mem_data[23];
  assign N351 = atomic_reg_data[22] ^ atomic_mem_data[22];
  assign N352 = atomic_reg_data[21] ^ atomic_mem_data[21];
  assign N353 = atomic_reg_data[20] ^ atomic_mem_data[20];
  assign N354 = atomic_reg_data[19] ^ atomic_mem_data[19];
  assign N355 = atomic_reg_data[18] ^ atomic_mem_data[18];
  assign N356 = atomic_reg_data[17] ^ atomic_mem_data[17];
  assign N357 = atomic_reg_data[16] ^ atomic_mem_data[16];
  assign N358 = atomic_reg_data[15] ^ atomic_mem_data[15];
  assign N359 = atomic_reg_data[14] ^ atomic_mem_data[14];
  assign N360 = atomic_reg_data[13] ^ atomic_mem_data[13];
  assign N361 = atomic_reg_data[12] ^ atomic_mem_data[12];
  assign N362 = atomic_reg_data[11] ^ atomic_mem_data[11];
  assign N363 = atomic_reg_data[10] ^ atomic_mem_data[10];
  assign N364 = atomic_reg_data[9] ^ atomic_mem_data[9];
  assign N365 = atomic_reg_data[8] ^ atomic_mem_data[8];
  assign N366 = atomic_reg_data[7] ^ atomic_mem_data[7];
  assign N367 = atomic_reg_data[6] ^ atomic_mem_data[6];
  assign N368 = atomic_reg_data[5] ^ atomic_mem_data[5];
  assign N369 = atomic_reg_data[4] ^ atomic_mem_data[4];
  assign N370 = atomic_reg_data[3] ^ atomic_mem_data[3];
  assign N371 = atomic_reg_data[2] ^ atomic_mem_data[2];
  assign N372 = atomic_reg_data[1] ^ atomic_mem_data[1];
  assign N373 = atomic_reg_data[0] ^ atomic_mem_data[0];
  assign N439 = ~N438;
  assign N505 = ~N504;
  assign N571 = ~N570;
  assign N637 = ~N636;
  assign N766 = decode_tv_r_amo_op_;
  assign N767 = ~N766;
  assign N768 = ~N782;
  assign wbuf_entry_in_bank_sel__7_ = ld_data_way_select_tv[7] | decode_tv_r_block_op_;
  assign wbuf_entry_in_bank_sel__6_ = ld_data_way_select_tv[6] | decode_tv_r_block_op_;
  assign wbuf_entry_in_bank_sel__5_ = ld_data_way_select_tv[5] | decode_tv_r_block_op_;
  assign wbuf_entry_in_bank_sel__4_ = ld_data_way_select_tv[4] | decode_tv_r_block_op_;
  assign wbuf_entry_in_bank_sel__3_ = ld_data_way_select_tv[3] | decode_tv_r_block_op_;
  assign wbuf_entry_in_bank_sel__2_ = ld_data_way_select_tv[2] | decode_tv_r_block_op_;
  assign wbuf_entry_in_bank_sel__1_ = ld_data_way_select_tv[1] | decode_tv_r_block_op_;
  assign wbuf_entry_in_bank_sel__0_ = ld_data_way_select_tv[0] | decode_tv_r_block_op_;
  assign load_req = N1454 & N1455;
  assign N1454 = N1453 & load_miss_tv;
  assign N1453 = v_tv_r & N1452;
  assign N1452 = ~uncached_tv_r;
  assign N1455 = ~late_o;
  assign store_req = N1458 & N1459;
  assign N1458 = N1457 & store_miss_tv;
  assign N1457 = v_tv_r & N1456;
  assign N1456 = ~uncached_tv_r;
  assign N1459 = ~late_o;
  assign uncached_amo_req = N1462 & N1463;
  assign N1462 = N1461 & ret_o;
  assign N1461 = N1460 & decode_tv_r_amo_op_;
  assign N1460 = v_tv_r & uncached_tv_r;
  assign N1463 = ~late_o;
  assign uncached_load_req = N1467 & N1468;
  assign N1467 = N1466 & decode_tv_r_load_op_;
  assign N1466 = N1464 & N1465;
  assign N1464 = v_tv_r & uncached_tv_r;
  assign N1465 = ~decode_tv_r_amo_op_;
  assign N1468 = ~late_o;
  assign uncached_store_req = N1472 & N1473;
  assign N1472 = N1470 & N1471;
  assign N1470 = N1469 & decode_tv_r_store_op_;
  assign N1469 = v_tv_r & uncached_tv_r;
  assign N1471 = ~ret_o;
  assign N1473 = ~late_o;
  assign bclean_req = N1477 & N1478;
  assign N1477 = N1476 & store_hit_tv;
  assign N1476 = N1475 & decode_tv_r_bclean_op_;
  assign N1475 = v_tv_r & N1474;
  assign N1474 = ~uncached_tv_r;
  assign N1478 = ~late_o;
  assign inval_req = N1483 & N1484;
  assign N1483 = N1481 & N1482;
  assign N1481 = N1480 & decode_tv_r_inval_op_;
  assign N1480 = v_tv_r & N1479;
  assign N1479 = ~uncached_tv_r;
  assign N1482 = ~decode_tv_r_clean_op_;
  assign N1484 = ~late_o;
  assign clean_req = N1489 & N1490;
  assign N1489 = N1487 & N1488;
  assign N1487 = N1486 & decode_tv_r_clean_op_;
  assign N1486 = v_tv_r & N1485;
  assign N1485 = ~uncached_tv_r;
  assign N1488 = ~decode_tv_r_inval_op_;
  assign N1490 = ~late_o;
  assign flush_req = N1494 & N1495;
  assign N1494 = N1493 & decode_tv_r_clean_op_;
  assign N1493 = N1492 & decode_tv_r_inval_op_;
  assign N1492 = v_tv_r & N1491;
  assign N1491 = ~uncached_tv_r;
  assign N1495 = ~late_o;
  assign nonblocking_req = N1496 | N1498;
  assign N1496 = uncached_store_req | 1'b0;
  assign N1498 = N1497 | 1'b0;
  assign N1497 = 1'b0 | bclean_req;
  assign blocking_miss_tv = N1501 | N1503;
  assign N1501 = N1500 | uncached_load_req;
  assign N1500 = N1499 | uncached_amo_req;
  assign N1499 = load_req | store_req;
  assign N1503 = N1502 | flush_req;
  assign N1502 = inval_req | clean_req;
  assign blocking_sent = blocking_miss_tv & cache_req_yumi_i;
  assign cache_req_v_o = N1326 & N1504;
  assign N1504 = blocking_miss_tv | nonblocking_req;
  assign blocking_hazard = cache_req_v_o & blocking_miss_tv;
  assign nonblocking_hazard = nonblocking_req & N1505;
  assign N1505 = ~cache_req_yumi_i;
  assign N769 = N1509 | clean_req;
  assign N1509 = N1508 | inval_req;
  assign N1508 = N1507 | 1'b0;
  assign N1507 = N1506 | bclean_req;
  assign N1506 = load_req | store_req;
  assign N770 = decode_tv_r_block_op_;
  assign N771 = decode_tv_r_double_op_;
  assign N772 = decode_tv_r_word_op_;
  assign N773 = decode_tv_r_half_op_;
  assign N774 = N770 | N769;
  assign N775 = N771 | N774;
  assign N776 = N772 | N775;
  assign N777 = N773 | N776;
  assign N778 = ~N777;
  assign N779 = ~N776;
  assign N780 = ~N774;
  assign N781 = ~decode_tv_r_amo_op_;
  assign N782 = decode_tv_r_amo_op_;
  assign N783 = ~decode_tv_r_amo_subop__0_;
  assign N787 = ~N786;
  assign N788 = ~decode_tv_r_amo_subop__1_;
  assign N791 = ~N790;
  assign N794 = ~N793;
  assign N795 = ~decode_tv_r_amo_subop__2_;
  assign N799 = ~N798;
  assign N801 = ~N800;
  assign N803 = ~N802;
  assign N805 = ~N804;
  assign N806 = ~decode_tv_r_amo_subop__3_;
  assign N809 = ~N808;
  assign N811 = ~N810;
  assign N813 = ~N812;
  assign N815 = ~N814;
  assign N820 = N816 | N819;
  assign N825 = 1'b0;
  assign N826 = 1'b0;
  assign N827 = bclean_req | N825;
  assign N828 = N826 | N827;
  assign N829 = inval_req | N828;
  assign N830 = clean_req | N829;
  assign N831 = flush_req | N830;
  assign N832 = store_req | N831;
  assign N833 = load_req | N832;
  assign N834 = uncached_amo_req | N833;
  assign N835 = uncached_store_req | N834;
  assign N836 = uncached_load_req | N835;
  assign N837 = ~N836;
  assign N838 = ~N835;
  assign N839 = ~N831;
  assign N840 = ~N769;
  assign N841 = N770 & N840;
  assign N842 = ~N770;
  assign N843 = N840 & N842;
  assign N844 = N771 & N843;
  assign N845 = ~N771;
  assign N846 = N843 & N845;
  assign N847 = N772 & N846;
  assign N848 = ~N772;
  assign N849 = N846 & N848;
  assign N850 = N773 & N849;
  assign N851 = ~N825;
  assign N852 = bclean_req & N851;
  assign N853 = ~bclean_req;
  assign N854 = N851 & N853;
  assign N855 = N826 & N854;
  assign N856 = ~N826;
  assign N857 = N854 & N856;
  assign N858 = inval_req & N857;
  assign N859 = ~inval_req;
  assign N860 = N857 & N859;
  assign N861 = clean_req & N860;
  assign N862 = ~clean_req;
  assign N863 = N860 & N862;
  assign N864 = flush_req & N863;
  assign N865 = ~flush_req;
  assign N866 = N863 & N865;
  assign N867 = store_req & N866;
  assign N868 = ~store_req;
  assign N869 = N866 & N868;
  assign N870 = load_req & N869;
  assign N871 = ~load_req;
  assign N872 = N869 & N871;
  assign N873 = uncached_amo_req & N872;
  assign N874 = ~uncached_amo_req;
  assign N875 = N872 & N874;
  assign N876 = uncached_store_req & N875;
  assign N877 = ~uncached_store_req;
  assign N878 = N875 & N877;
  assign N879 = uncached_load_req & N878;
  assign _14_net__7_ = ~metadata_way_v_r[7];
  assign _14_net__6_ = ~metadata_way_v_r[6];
  assign _14_net__5_ = ~metadata_way_v_r[5];
  assign _14_net__4_ = ~metadata_way_v_r[4];
  assign _14_net__3_ = ~metadata_way_v_r[3];
  assign _14_net__2_ = ~metadata_way_v_r[2];
  assign _14_net__1_ = ~metadata_way_v_r[1];
  assign _14_net__0_ = ~metadata_way_v_r[0];
  assign N880 = ~metadata_invalid_exist;
  assign N881 = ~metadata_hit_r;
  assign N882 = ~cache_req_metadata_o[1];
  assign N883 = ~cache_req_metadata_o[2];
  assign N884 = N882 & N883;
  assign N885 = N882 & cache_req_metadata_o[2];
  assign N886 = cache_req_metadata_o[1] & N883;
  assign N887 = cache_req_metadata_o[1] & cache_req_metadata_o[2];
  assign N888 = ~cache_req_metadata_o[3];
  assign N889 = N884 & N888;
  assign N890 = N884 & cache_req_metadata_o[3];
  assign N891 = N886 & N888;
  assign N892 = N886 & cache_req_metadata_o[3];
  assign N893 = N885 & N888;
  assign N894 = N885 & cache_req_metadata_o[3];
  assign N895 = N887 & N888;
  assign N896 = N887 & cache_req_metadata_o[3];
  assign busy_o = cache_req_lock_i | N1511;
  assign N1511 = ~N1510;
  assign N1510 = N1326 | N1329;
  assign ordered_o = N1514 & cache_req_credits_empty_i;
  assign N1514 = N1512 & N1513;
  assign N1512 = ~v_tl_r;
  assign N1513 = ~v_tv_r;
  assign tag_mem_fast_read = safe_tl_we & N1515;
  assign N1515 = ~decode_lo[23];
  assign tag_mem_slow_read = tag_mem_pkt_yumi_o & N1246;
  assign tag_mem_slow_write = tag_mem_pkt_yumi_o & N1249;
  assign tag_mem_fast_write = N1519 | N1522;
  assign N1519 = N1517 & N1518;
  assign N1517 = N1516 & cache_req_o[115];
  assign N1516 = v_tv_r & uncached_tv_r;
  assign N1518 = ~late_o;
  assign N1522 = N1521 & N1518;
  assign N1521 = N1520 & cache_req_o[115];
  assign N1520 = v_tv_r & decode_tv_r_binval_op_;
  assign tag_mem_v_li = N1524 | tag_mem_fast_write;
  assign N1524 = N1523 | tag_mem_slow_write;
  assign N1523 = tag_mem_fast_read | tag_mem_slow_read;
  assign tag_mem_w_li = tag_mem_slow_write | tag_mem_fast_write;
  assign N897 = tag_mem_fast_read | tag_mem_fast_write;
  assign N898 = ~N897;
  assign N899 = ~tag_mem_fast_write;
  assign N900 = tag_mem_fast_read & N899;
  assign tag_mem_pkt_yumi_o = N1530 & N1531;
  assign N1530 = N1528 & N1529;
  assign N1528 = N1526 & N1527;
  assign N1526 = tag_mem_pkt_v_i & N1525;
  assign N1525 = ~N1318;
  assign N1527 = ~tag_mem_fast_read;
  assign N1529 = ~tag_mem_fast_write;
  assign N1531 = ~wbuf_snoop_match_lo;
  assign N901 = ~tag_mem_pkt_i[0];
  assign N905 = ~N904;
  assign N906 = ~tag_mem_pkt_i[1];
  assign N910 = ~N909;
  assign N911 = ~tag_mem_pkt_i[1];
  assign N912 = ~tag_mem_pkt_i[0];
  assign N916 = ~N915;
  assign N918 = ~tag_mem_pkt_i[1];
  assign N919 = ~tag_mem_pkt_i[0];
  assign N922 = N917 | N921;
  assign N923 = ~tag_mem_pkt_i[0];
  assign N927 = ~N926;
  assign N928 = ~tag_mem_pkt_i[1];
  assign N932 = ~N931;
  assign N933 = ~tag_mem_pkt_i[1];
  assign N934 = ~tag_mem_pkt_i[0];
  assign N938 = ~N937;
  assign N940 = ~tag_mem_pkt_i[1];
  assign N941 = ~tag_mem_pkt_i[0];
  assign N944 = N939 | N943;
  assign N945 = ~tag_mem_pkt_i[0];
  assign N949 = ~N948;
  assign N950 = ~tag_mem_pkt_i[1];
  assign N954 = ~N953;
  assign N955 = ~tag_mem_pkt_i[1];
  assign N956 = ~tag_mem_pkt_i[0];
  assign N960 = ~N959;
  assign N962 = ~tag_mem_pkt_i[1];
  assign N963 = ~tag_mem_pkt_i[0];
  assign N966 = N961 | N965;
  assign N967 = ~tag_mem_pkt_i[0];
  assign N971 = ~N970;
  assign N972 = ~tag_mem_pkt_i[1];
  assign N976 = ~N975;
  assign N977 = ~tag_mem_pkt_i[1];
  assign N978 = ~tag_mem_pkt_i[0];
  assign N982 = ~N981;
  assign N984 = ~tag_mem_pkt_i[1];
  assign N985 = ~tag_mem_pkt_i[0];
  assign N988 = N983 | N987;
  assign N989 = ~tag_mem_pkt_i[0];
  assign N993 = ~N992;
  assign N994 = ~tag_mem_pkt_i[1];
  assign N998 = ~N997;
  assign N999 = ~tag_mem_pkt_i[1];
  assign N1000 = ~tag_mem_pkt_i[0];
  assign N1004 = ~N1003;
  assign N1006 = ~tag_mem_pkt_i[1];
  assign N1007 = ~tag_mem_pkt_i[0];
  assign N1010 = N1005 | N1009;
  assign N1011 = ~tag_mem_pkt_i[0];
  assign N1015 = ~N1014;
  assign N1016 = ~tag_mem_pkt_i[1];
  assign N1020 = ~N1019;
  assign N1021 = ~tag_mem_pkt_i[1];
  assign N1022 = ~tag_mem_pkt_i[0];
  assign N1026 = ~N1025;
  assign N1028 = ~tag_mem_pkt_i[1];
  assign N1029 = ~tag_mem_pkt_i[0];
  assign N1032 = N1027 | N1031;
  assign N1033 = ~tag_mem_pkt_i[0];
  assign N1037 = ~N1036;
  assign N1038 = ~tag_mem_pkt_i[1];
  assign N1042 = ~N1041;
  assign N1043 = ~tag_mem_pkt_i[1];
  assign N1044 = ~tag_mem_pkt_i[0];
  assign N1048 = ~N1047;
  assign N1050 = ~tag_mem_pkt_i[1];
  assign N1051 = ~tag_mem_pkt_i[0];
  assign N1054 = N1049 | N1053;
  assign N1055 = ~tag_mem_pkt_i[0];
  assign N1059 = ~N1058;
  assign N1060 = ~tag_mem_pkt_i[1];
  assign N1064 = ~N1063;
  assign N1065 = ~tag_mem_pkt_i[1];
  assign N1066 = ~tag_mem_pkt_i[0];
  assign N1070 = ~N1069;
  assign N1072 = ~tag_mem_pkt_i[1];
  assign N1073 = ~tag_mem_pkt_i[0];
  assign N1076 = N1071 | N1075;
  assign N1077 = ~tag_mem_pkt_way_r[0];
  assign N1078 = ~tag_mem_pkt_way_r[1];
  assign N1079 = N1077 & N1078;
  assign N1080 = N1077 & tag_mem_pkt_way_r[1];
  assign N1081 = tag_mem_pkt_way_r[0] & N1078;
  assign N1082 = tag_mem_pkt_way_r[0] & tag_mem_pkt_way_r[1];
  assign N1083 = ~tag_mem_pkt_way_r[2];
  assign N1084 = N1079 & N1083;
  assign N1085 = N1079 & tag_mem_pkt_way_r[2];
  assign N1086 = N1081 & N1083;
  assign N1087 = N1081 & tag_mem_pkt_way_r[2];
  assign N1088 = N1080 & N1083;
  assign N1089 = N1080 & tag_mem_pkt_way_r[2];
  assign N1090 = N1082 & N1083;
  assign N1091 = N1082 & tag_mem_pkt_way_r[2];
  assign data_mem_fast_read[0] = safe_tl_we & decode_lo[30];
  assign data_mem_force_write[0] = N1532 & wbuf_entry_out_bank_sel__0_;
  assign N1532 = wbuf_v_lo & wbuf_force_lo;
  assign data_mem_slow_write[0] = N1533 & data_mem_write_bank_mask[0];
  assign N1533 = data_mem_pkt_yumi_o & N1254;
  assign data_mem_slow_read[0] = data_mem_pkt_yumi_o & N1252;
  assign data_mem_fast_write[0] = wbuf_yumi_li & wbuf_entry_out_bank_sel__0_;
  assign data_mem_v_li[0] = N1535 | data_mem_slow_write[0];
  assign N1535 = N1534 | data_mem_slow_read[0];
  assign N1534 = data_mem_fast_read[0] | data_mem_fast_write[0];
  assign data_mem_w_li[0] = data_mem_fast_write[0] | data_mem_slow_write[0];
  assign N1092 = ~data_mem_fast_write[0];
  assign N1093 = data_mem_fast_read[0] | data_mem_fast_write[0];
  assign N1094 = ~N1093;
  assign N1095 = data_mem_fast_read[0] & N1092;
  assign data_mem_force_write[1] = N1536 & wbuf_entry_out_bank_sel__1_;
  assign N1536 = wbuf_v_lo & wbuf_force_lo;
  assign data_mem_slow_write[1] = N1537 & data_mem_write_bank_mask[1];
  assign N1537 = data_mem_pkt_yumi_o & N1259;
  assign data_mem_slow_read[1] = data_mem_pkt_yumi_o & N1257;
  assign data_mem_fast_write[1] = wbuf_yumi_li & wbuf_entry_out_bank_sel__1_;
  assign data_mem_v_li[1] = N1539 | data_mem_slow_write[1];
  assign N1539 = N1538 | data_mem_slow_read[1];
  assign N1538 = data_mem_fast_read[0] | data_mem_fast_write[1];
  assign data_mem_w_li[1] = data_mem_fast_write[1] | data_mem_slow_write[1];
  assign N1096 = ~data_mem_fast_write[1];
  assign N1097 = data_mem_fast_read[0] | data_mem_fast_write[1];
  assign N1098 = ~N1097;
  assign N1099 = data_mem_fast_read[0] & N1096;
  assign data_mem_force_write[2] = N1540 & wbuf_entry_out_bank_sel__2_;
  assign N1540 = wbuf_v_lo & wbuf_force_lo;
  assign data_mem_slow_write[2] = N1541 & data_mem_write_bank_mask[2];
  assign N1541 = data_mem_pkt_yumi_o & N1264;
  assign data_mem_slow_read[2] = data_mem_pkt_yumi_o & N1262;
  assign data_mem_fast_write[2] = wbuf_yumi_li & wbuf_entry_out_bank_sel__2_;
  assign data_mem_v_li[2] = N1543 | data_mem_slow_write[2];
  assign N1543 = N1542 | data_mem_slow_read[2];
  assign N1542 = data_mem_fast_read[0] | data_mem_fast_write[2];
  assign data_mem_w_li[2] = data_mem_fast_write[2] | data_mem_slow_write[2];
  assign N1100 = ~data_mem_fast_write[2];
  assign N1101 = data_mem_fast_read[0] | data_mem_fast_write[2];
  assign N1102 = ~N1101;
  assign N1103 = data_mem_fast_read[0] & N1100;
  assign data_mem_force_write[3] = N1544 & wbuf_entry_out_bank_sel__3_;
  assign N1544 = wbuf_v_lo & wbuf_force_lo;
  assign data_mem_slow_write[3] = N1545 & data_mem_write_bank_mask[3];
  assign N1545 = data_mem_pkt_yumi_o & N1269;
  assign data_mem_slow_read[3] = data_mem_pkt_yumi_o & N1267;
  assign data_mem_fast_write[3] = wbuf_yumi_li & wbuf_entry_out_bank_sel__3_;
  assign data_mem_v_li[3] = N1547 | data_mem_slow_write[3];
  assign N1547 = N1546 | data_mem_slow_read[3];
  assign N1546 = data_mem_fast_read[0] | data_mem_fast_write[3];
  assign data_mem_w_li[3] = data_mem_fast_write[3] | data_mem_slow_write[3];
  assign N1104 = ~data_mem_fast_write[3];
  assign N1105 = data_mem_fast_read[0] | data_mem_fast_write[3];
  assign N1106 = ~N1105;
  assign N1107 = data_mem_fast_read[0] & N1104;
  assign data_mem_force_write[4] = N1548 & wbuf_entry_out_bank_sel__4_;
  assign N1548 = wbuf_v_lo & wbuf_force_lo;
  assign data_mem_slow_write[4] = N1549 & data_mem_write_bank_mask[4];
  assign N1549 = data_mem_pkt_yumi_o & N1274;
  assign data_mem_slow_read[4] = data_mem_pkt_yumi_o & N1272;
  assign data_mem_fast_write[4] = wbuf_yumi_li & wbuf_entry_out_bank_sel__4_;
  assign data_mem_v_li[4] = N1551 | data_mem_slow_write[4];
  assign N1551 = N1550 | data_mem_slow_read[4];
  assign N1550 = data_mem_fast_read[0] | data_mem_fast_write[4];
  assign data_mem_w_li[4] = data_mem_fast_write[4] | data_mem_slow_write[4];
  assign N1108 = ~data_mem_fast_write[4];
  assign N1109 = data_mem_fast_read[0] | data_mem_fast_write[4];
  assign N1110 = ~N1109;
  assign N1111 = data_mem_fast_read[0] & N1108;
  assign data_mem_force_write[5] = N1552 & wbuf_entry_out_bank_sel__5_;
  assign N1552 = wbuf_v_lo & wbuf_force_lo;
  assign data_mem_slow_write[5] = N1553 & data_mem_write_bank_mask[5];
  assign N1553 = data_mem_pkt_yumi_o & N1279;
  assign data_mem_slow_read[5] = data_mem_pkt_yumi_o & N1277;
  assign data_mem_fast_write[5] = wbuf_yumi_li & wbuf_entry_out_bank_sel__5_;
  assign data_mem_v_li[5] = N1555 | data_mem_slow_write[5];
  assign N1555 = N1554 | data_mem_slow_read[5];
  assign N1554 = data_mem_fast_read[0] | data_mem_fast_write[5];
  assign data_mem_w_li[5] = data_mem_fast_write[5] | data_mem_slow_write[5];
  assign N1112 = ~data_mem_fast_write[5];
  assign N1113 = data_mem_fast_read[0] | data_mem_fast_write[5];
  assign N1114 = ~N1113;
  assign N1115 = data_mem_fast_read[0] & N1112;
  assign data_mem_force_write[6] = N1556 & wbuf_entry_out_bank_sel__6_;
  assign N1556 = wbuf_v_lo & wbuf_force_lo;
  assign data_mem_slow_write[6] = N1557 & data_mem_write_bank_mask[6];
  assign N1557 = data_mem_pkt_yumi_o & N1284;
  assign data_mem_slow_read[6] = data_mem_pkt_yumi_o & N1282;
  assign data_mem_fast_write[6] = wbuf_yumi_li & wbuf_entry_out_bank_sel__6_;
  assign data_mem_v_li[6] = N1559 | data_mem_slow_write[6];
  assign N1559 = N1558 | data_mem_slow_read[6];
  assign N1558 = data_mem_fast_read[0] | data_mem_fast_write[6];
  assign data_mem_w_li[6] = data_mem_fast_write[6] | data_mem_slow_write[6];
  assign N1116 = ~data_mem_fast_write[6];
  assign N1117 = data_mem_fast_read[0] | data_mem_fast_write[6];
  assign N1118 = ~N1117;
  assign N1119 = data_mem_fast_read[0] & N1116;
  assign data_mem_force_write[7] = N1560 & wbuf_entry_out_bank_sel__7_;
  assign N1560 = wbuf_v_lo & wbuf_force_lo;
  assign data_mem_slow_write[7] = N1561 & data_mem_write_bank_mask[7];
  assign N1561 = data_mem_pkt_yumi_o & N1289;
  assign data_mem_slow_read[7] = data_mem_pkt_yumi_o & N1287;
  assign data_mem_fast_write[7] = wbuf_yumi_li & wbuf_entry_out_bank_sel__7_;
  assign data_mem_v_li[7] = N1563 | data_mem_slow_write[7];
  assign N1563 = N1562 | data_mem_slow_read[7];
  assign N1562 = data_mem_fast_read[0] | data_mem_fast_write[7];
  assign data_mem_w_li[7] = data_mem_fast_write[7] | data_mem_slow_write[7];
  assign N1120 = ~data_mem_fast_write[7];
  assign N1121 = data_mem_fast_read[0] | data_mem_fast_write[7];
  assign N1122 = ~N1121;
  assign N1123 = data_mem_fast_read[0] & N1120;
  assign wbuf_yumi_li = wbuf_v_lo & N1580;
  assign N1580 = N1579 | wbuf_force_lo;
  assign N1579 = ~N1578;
  assign N1578 = N1576 | N1577;
  assign N1576 = N1574 | N1575;
  assign N1574 = N1572 | N1573;
  assign N1572 = N1570 | N1571;
  assign N1570 = N1568 | N1569;
  assign N1568 = N1566 | N1567;
  assign N1566 = N1564 | N1565;
  assign N1564 = data_mem_fast_read[0] & wbuf_entry_out_bank_sel__7_;
  assign N1565 = data_mem_fast_read[0] & wbuf_entry_out_bank_sel__6_;
  assign N1567 = data_mem_fast_read[0] & wbuf_entry_out_bank_sel__5_;
  assign N1569 = data_mem_fast_read[0] & wbuf_entry_out_bank_sel__4_;
  assign N1571 = data_mem_fast_read[0] & wbuf_entry_out_bank_sel__3_;
  assign N1573 = data_mem_fast_read[0] & wbuf_entry_out_bank_sel__2_;
  assign N1575 = data_mem_fast_read[0] & wbuf_entry_out_bank_sel__1_;
  assign N1577 = data_mem_fast_read[0] & wbuf_entry_out_bank_sel__0_;
  assign data_mem_write_hazard = N1593 | N1594;
  assign N1593 = N1591 | N1592;
  assign N1591 = N1589 | N1590;
  assign N1589 = N1587 | N1588;
  assign N1587 = N1585 | N1586;
  assign N1585 = N1583 | N1584;
  assign N1583 = N1581 | N1582;
  assign N1581 = data_mem_fast_read[0] & data_mem_force_write[7];
  assign N1582 = data_mem_fast_read[0] & data_mem_force_write[6];
  assign N1584 = data_mem_fast_read[0] & data_mem_force_write[5];
  assign N1586 = data_mem_fast_read[0] & data_mem_force_write[4];
  assign N1588 = data_mem_fast_read[0] & data_mem_force_write[3];
  assign N1590 = data_mem_fast_read[0] & data_mem_force_write[2];
  assign N1592 = data_mem_fast_read[0] & data_mem_force_write[1];
  assign N1594 = data_mem_fast_read[0] & data_mem_force_write[0];
  assign data_mem_pkt_yumi_o = N1652 & N1531;
  assign N1652 = N1649 & N1651;
  assign N1649 = N1632 & N1648;
  assign N1632 = N1615 & N1631;
  assign N1615 = N1605 & N1614;
  assign N1605 = N1595 & N1604;
  assign N1595 = data_mem_pkt_v_i & N1525;
  assign N1604 = ~N1603;
  assign N1603 = N1602 & N1321;
  assign N1602 = N1601 | data_mem_fast_read[0];
  assign N1601 = N1600 | data_mem_fast_read[0];
  assign N1600 = N1599 | data_mem_fast_read[0];
  assign N1599 = N1598 | data_mem_fast_read[0];
  assign N1598 = N1597 | data_mem_fast_read[0];
  assign N1597 = N1596 | data_mem_fast_read[0];
  assign N1596 = data_mem_fast_read[0] | data_mem_fast_read[0];
  assign N1614 = ~N1613;
  assign N1613 = N1612 & N1324;
  assign N1612 = N1611 | data_mem_fast_write[0];
  assign N1611 = N1610 | data_mem_fast_write[1];
  assign N1610 = N1609 | data_mem_fast_write[2];
  assign N1609 = N1608 | data_mem_fast_write[3];
  assign N1608 = N1607 | data_mem_fast_write[4];
  assign N1607 = N1606 | data_mem_fast_write[5];
  assign N1606 = data_mem_fast_write[7] | data_mem_fast_write[6];
  assign N1631 = ~N1630;
  assign N1630 = N1628 | N1629;
  assign N1628 = N1626 | N1627;
  assign N1626 = N1624 | N1625;
  assign N1624 = N1622 | N1623;
  assign N1622 = N1620 | N1621;
  assign N1620 = N1618 | N1619;
  assign N1618 = N1616 | N1617;
  assign N1616 = data_mem_fast_read[0] & data_mem_write_bank_mask[7];
  assign N1617 = data_mem_fast_read[0] & data_mem_write_bank_mask[6];
  assign N1619 = data_mem_fast_read[0] & data_mem_write_bank_mask[5];
  assign N1621 = data_mem_fast_read[0] & data_mem_write_bank_mask[4];
  assign N1623 = data_mem_fast_read[0] & data_mem_write_bank_mask[3];
  assign N1625 = data_mem_fast_read[0] & data_mem_write_bank_mask[2];
  assign N1627 = data_mem_fast_read[0] & data_mem_write_bank_mask[1];
  assign N1629 = data_mem_fast_read[0] & data_mem_write_bank_mask[0];
  assign N1648 = ~N1647;
  assign N1647 = N1645 | N1646;
  assign N1645 = N1643 | N1644;
  assign N1643 = N1641 | N1642;
  assign N1641 = N1639 | N1640;
  assign N1639 = N1637 | N1638;
  assign N1637 = N1635 | N1636;
  assign N1635 = N1633 | N1634;
  assign N1633 = data_mem_fast_write[7] & data_mem_write_bank_mask[7];
  assign N1634 = data_mem_fast_write[6] & data_mem_write_bank_mask[6];
  assign N1636 = data_mem_fast_write[5] & data_mem_write_bank_mask[5];
  assign N1638 = data_mem_fast_write[4] & data_mem_write_bank_mask[4];
  assign N1640 = data_mem_fast_write[3] & data_mem_write_bank_mask[3];
  assign N1642 = data_mem_fast_write[2] & data_mem_write_bank_mask[2];
  assign N1644 = data_mem_fast_write[1] & data_mem_write_bank_mask[1];
  assign N1646 = data_mem_fast_write[0] & data_mem_write_bank_mask[0];
  assign N1651 = ~N1650;
  assign N1650 = v_tl_r & cache_req_critical_i;
  assign stat_mem_fast_read = N1653 & N1654;
  assign N1653 = v_tv_r & cache_req_yumi_i;
  assign N1654 = ~decode_tv_r_cache_op_;
  assign stat_mem_fast_write = N1659 & N1660;
  assign N1659 = N1657 & N1658;
  assign N1657 = N1655 & N1656;
  assign N1655 = v_tv_r & cache_req_o[115];
  assign N1656 = ~decode_tv_r_cache_op_;
  assign N1658 = ~uncached_tv_r;
  assign N1660 = ~cache_req_yumi_i;
  assign stat_mem_slow_write = stat_mem_pkt_yumi_o & N1294;
  assign stat_mem_slow_read = stat_mem_pkt_yumi_o & N1292;
  assign stat_mem_v_li = N1661 | N1662;
  assign N1661 = stat_mem_fast_read | stat_mem_fast_write;
  assign N1662 = stat_mem_slow_write | stat_mem_slow_read;
  assign stat_mem_w_li = stat_mem_fast_write | stat_mem_slow_write;
  assign N1124 = stat_mem_fast_write | stat_mem_fast_read;
  assign N1125 = ~N1124;
  assign stat_mem_pkt_yumi_o = N1667 & N1669;
  assign N1667 = N1665 & N1666;
  assign N1665 = N1663 & N1664;
  assign N1663 = stat_mem_pkt_v_i & N1525;
  assign N1664 = ~stat_mem_fast_read;
  assign N1666 = ~stat_mem_fast_write;
  assign N1669 = ~N1668;
  assign N1668 = wbuf_snoop_match_lo & N1315;
  assign N1126 = decode_tv_r_store_op_;
  assign N1127 = ~N1126;
  assign \tdm.dirty_mask_v_li  = stat_mem_slow_write | N1670;
  assign N1670 = v_tv_r & decode_tv_r_store_op_;
  assign N1131 = ~stat_mem_pkt_i[0];
  assign N1133 = ~N1132;
  assign N1134 = ~stat_mem_pkt_i[1];
  assign N1135 = stat_mem_pkt_i[1];
  assign \l1_lrsc.set_reservation  = N1671 & store_hit_tv;
  assign N1671 = v_tv_r & decode_tv_r_lr_op_;
  assign \l1_lrsc.clear_reservation  = N1672 | N1675;
  assign N1672 = v_tv_r & decode_tv_r_sc_op_;
  assign N1675 = N1674 & N1145;
  assign N1674 = N1673 & N1144;
  assign N1673 = tag_mem_pkt_yumi_o & \l1_lrsc.load_reserved_v_r ;
  assign \l1_lrsc.load_reservation_match_tv  = N1676 & N1147;
  assign N1676 = \l1_lrsc.load_reserved_v_r  & N1146;
  assign sc_success_tv = N1678 & \l1_lrsc.load_reservation_match_tv ;
  assign N1678 = N1677 & store_hit_tv;
  assign N1677 = v_tv_r & decode_tv_r_sc_op_;
  assign sc_fail_tv = N1679 & N1680;
  assign N1679 = v_tv_r & decode_tv_r_sc_op_;
  assign N1680 = ~sc_success_tv;
  assign \l1_lrsc.lrsc_lock_up  = sc_fail_tv | N1318;
  assign N1148 = N1325 & complete_recv;
  assign N1149 = N1326 & blocking_sent;
  assign N1150 = N1681 & any_miss_tv;
  assign N1681 = N1329 & v_tv_r;
  assign N1151 = N1149 | N1148;
  assign N1152 = N1150 | N1151;
  assign N1153 = ~N1152;
  assign N1155 = decode_tv_r_cache_op_;
  assign N1156 = ~N1148;
  assign N1157 = N1149 & N1156;
  assign N1158 = ~N1149;
  assign N1159 = N1156 & N1158;
  assign N1160 = N1150 & N1159;
  assign \hum.fill_v  = data_mem_pkt_v_i & N1312;
  assign \hum.fill_recv  = N1687 & N1689;
  assign N1687 = N1684 & N1686;
  assign N1684 = \hum.fill_v  & N1683;
  assign N1683 = N1682 | stat_mem_pkt_yumi_o;
  assign N1682 = ~stat_mem_pkt_v_i;
  assign N1686 = N1685 | tag_mem_pkt_yumi_o;
  assign N1685 = ~tag_mem_pkt_v_i;
  assign N1689 = N1688 | data_mem_pkt_yumi_o;
  assign N1688 = ~data_mem_pkt_v_i;
  assign N1161 = ~\hum.fill_v ;
  assign N1162 = \hum.fill_bank_mask_r [7] & N1690;
  assign N1690 = ~data_mem_pkt_fill_mask_expanded[7];
  assign N1163 = \hum.fill_bank_mask_r [6] & N1691;
  assign N1691 = ~data_mem_pkt_fill_mask_expanded[6];
  assign N1164 = \hum.fill_bank_mask_r [5] & N1692;
  assign N1692 = ~data_mem_pkt_fill_mask_expanded[5];
  assign N1165 = \hum.fill_bank_mask_r [4] & N1693;
  assign N1693 = ~data_mem_pkt_fill_mask_expanded[4];
  assign N1166 = \hum.fill_bank_mask_r [3] & N1694;
  assign N1694 = ~data_mem_pkt_fill_mask_expanded[3];
  assign N1167 = \hum.fill_bank_mask_r [2] & N1695;
  assign N1695 = ~data_mem_pkt_fill_mask_expanded[2];
  assign N1168 = \hum.fill_bank_mask_r [1] & N1696;
  assign N1696 = ~data_mem_pkt_fill_mask_expanded[1];
  assign N1169 = \hum.fill_bank_mask_r [0] & N1697;
  assign N1697 = ~data_mem_pkt_fill_mask_expanded[0];
  assign _25_net_ = \hum.fill_recv  | blocking_sent;
  assign fill_hazard = N1715 & N1730;
  assign N1715 = N1699 & N1714;
  assign N1699 = N1698 & N1178;
  assign N1698 = N1325 & v_tl_r;
  assign N1714 = N1712 | N1713;
  assign N1712 = N1710 | N1711;
  assign N1710 = N1708 | N1709;
  assign N1708 = N1706 | N1707;
  assign N1706 = N1704 | N1705;
  assign N1704 = N1702 | N1703;
  assign N1702 = N1700 | N1701;
  assign N1700 = \hum.fill_hit_r [7] & load_hit_tl[7];
  assign N1701 = \hum.fill_hit_r [6] & load_hit_tl[6];
  assign N1703 = \hum.fill_hit_r [5] & load_hit_tl[5];
  assign N1705 = \hum.fill_hit_r [4] & load_hit_tl[4];
  assign N1707 = \hum.fill_hit_r [3] & load_hit_tl[3];
  assign N1709 = \hum.fill_hit_r [2] & load_hit_tl[2];
  assign N1711 = \hum.fill_hit_r [1] & load_hit_tl[1];
  assign N1713 = \hum.fill_hit_r [0] & load_hit_tl[0];
  assign N1730 = N1728 | N1729;
  assign N1728 = N1726 | N1727;
  assign N1726 = N1724 | N1725;
  assign N1724 = N1722 | N1723;
  assign N1722 = N1720 | N1721;
  assign N1720 = N1718 | N1719;
  assign N1718 = N1716 | N1717;
  assign N1716 = \hum.fill_bank_mask_r [7] & bank_sel_one_hot_tl[7];
  assign N1717 = \hum.fill_bank_mask_r [6] & bank_sel_one_hot_tl[6];
  assign N1719 = \hum.fill_bank_mask_r [5] & bank_sel_one_hot_tl[5];
  assign N1721 = \hum.fill_bank_mask_r [4] & bank_sel_one_hot_tl[4];
  assign N1723 = \hum.fill_bank_mask_r [3] & bank_sel_one_hot_tl[3];
  assign N1725 = \hum.fill_bank_mask_r [2] & bank_sel_one_hot_tl[2];
  assign N1727 = \hum.fill_bank_mask_r [1] & bank_sel_one_hot_tl[1];
  assign N1729 = \hum.fill_bank_mask_r [0] & bank_sel_one_hot_tl[0];
  assign pseudo_hit[7] = N1186 | N1194;
  assign pseudo_hit[6] = N1185 | N1193;
  assign pseudo_hit[5] = N1184 | N1192;
  assign pseudo_hit[4] = N1183 | N1191;
  assign pseudo_hit[3] = N1182 | N1190;
  assign pseudo_hit[2] = N1181 | N1189;
  assign pseudo_hit[1] = N1180 | N1188;
  assign pseudo_hit[0] = N1179 | N1187;

  always @(posedge clk_i) begin
    if(reset_i) begin
      state_r_1_sv2v_reg <= 1'b0;
      state_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      state_r_1_sv2v_reg <= state_n[1];
      state_r_0_sv2v_reg <= state_n[0];
    end 
  end


endmodule

