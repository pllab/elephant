

module bsg_dff_reset_en_00000027_0_0
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [38:0] data_i;
  output [38:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [38:0] data_o;
  wire N0,N1,N2;
  reg data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,
  data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,
  data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,
  data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,
  data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,
  data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_en_bypass_00000027
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [38:0] data_i;
  output [38:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [38:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_reset_en_00000027_0_0
  dff
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(en_i),
    .data_i(data_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_dff_reset_set_clear_width_p2_clear_over_set_p1
(
  clk_i,
  reset_i,
  set_i,
  clear_i,
  data_o
);

  input [1:0] set_i;
  input [1:0] clear_i;
  output [1:0] data_o;
  input clk_i;
  input reset_i;
  wire [1:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  reg data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N0 = N2 & N3;
  assign N2 = data_o[1] | set_i[1];
  assign N3 = ~clear_i[1];
  assign N1 = N4 & N5;
  assign N4 = data_o[0] | set_i[0];
  assign N5 = ~clear_i[0];

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_1_sv2v_reg <= N0;
      data_o_0_sv2v_reg <= N1;
    end 
  end


endmodule



module bsg_circular_ptr_00000004_1
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [0:0] add_i;
  output [1:0] o;
  output [1:0] n_o;
  input clk;
  input reset_i;
  wire [1:0] o,n_o,\genblk1.genblk1.ptr_r_p1 ;
  wire N0,N1,N2;
  reg o_1_sv2v_reg,o_0_sv2v_reg;
  assign o[1] = o_1_sv2v_reg;
  assign o[0] = o_0_sv2v_reg;
  assign \genblk1.genblk1.ptr_r_p1  = o + 1'b1;
  assign n_o = (N0)? \genblk1.genblk1.ptr_r_p1  : 
               (N1)? o : 1'b0;
  assign N0 = add_i[0];
  assign N1 = N2;
  assign N2 = ~add_i[0];

  always @(posedge clk) begin
    if(reset_i) begin
      o_1_sv2v_reg <= 1'b0;
      o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      o_1_sv2v_reg <= n_o[1];
      o_0_sv2v_reg <= n_o[0];
    end 
  end


endmodule



module bsg_fifo_tracker_00000004
(
  clk_i,
  reset_i,
  enq_i,
  deq_i,
  wptr_r_o,
  rptr_r_o,
  rptr_n_o,
  full_o,
  empty_o
);

  output [1:0] wptr_r_o;
  output [1:0] rptr_r_o;
  output [1:0] rptr_n_o;
  input clk_i;
  input reset_i;
  input enq_i;
  input deq_i;
  output full_o;
  output empty_o;
  wire [1:0] wptr_r_o,rptr_r_o,rptr_n_o;
  wire full_o,empty_o,enq_r,deq_r,N0,equal_ptrs,sv2v_dc_1,sv2v_dc_2;
  reg deq_r_sv2v_reg,enq_r_sv2v_reg;
  assign deq_r = deq_r_sv2v_reg;
  assign enq_r = enq_r_sv2v_reg;

  bsg_circular_ptr_00000004_1
  rptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(deq_i),
    .o(rptr_r_o),
    .n_o(rptr_n_o)
  );


  bsg_circular_ptr_00000004_1
  wptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(enq_i),
    .o(wptr_r_o),
    .n_o({ sv2v_dc_1, sv2v_dc_2 })
  );

  assign equal_ptrs = rptr_r_o == wptr_r_o;
  assign N0 = enq_i | deq_i;
  assign empty_o = equal_ptrs & deq_r;
  assign full_o = equal_ptrs & enq_r;

  always @(posedge clk_i) begin
    if(reset_i) begin
      deq_r_sv2v_reg <= 1'b1;
      enq_r_sv2v_reg <= 1'b0;
    end else if(N0) begin
      deq_r_sv2v_reg <= deq_i;
      enq_r_sv2v_reg <= enq_i;
    end 
  end


endmodule



module bsg_mem_1r1w_synth_114_00000004_0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [1:0] w_addr_i;
  input [113:0] w_data_i;
  input [1:0] r_addr_i;
  output [113:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [113:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24;
  wire [455:0] \nz.mem ;
  reg \nz.mem_455_sv2v_reg ,\nz.mem_454_sv2v_reg ,\nz.mem_453_sv2v_reg ,
  \nz.mem_452_sv2v_reg ,\nz.mem_451_sv2v_reg ,\nz.mem_450_sv2v_reg ,\nz.mem_449_sv2v_reg ,
  \nz.mem_448_sv2v_reg ,\nz.mem_447_sv2v_reg ,\nz.mem_446_sv2v_reg ,
  \nz.mem_445_sv2v_reg ,\nz.mem_444_sv2v_reg ,\nz.mem_443_sv2v_reg ,\nz.mem_442_sv2v_reg ,
  \nz.mem_441_sv2v_reg ,\nz.mem_440_sv2v_reg ,\nz.mem_439_sv2v_reg ,\nz.mem_438_sv2v_reg ,
  \nz.mem_437_sv2v_reg ,\nz.mem_436_sv2v_reg ,\nz.mem_435_sv2v_reg ,
  \nz.mem_434_sv2v_reg ,\nz.mem_433_sv2v_reg ,\nz.mem_432_sv2v_reg ,\nz.mem_431_sv2v_reg ,
  \nz.mem_430_sv2v_reg ,\nz.mem_429_sv2v_reg ,\nz.mem_428_sv2v_reg ,\nz.mem_427_sv2v_reg ,
  \nz.mem_426_sv2v_reg ,\nz.mem_425_sv2v_reg ,\nz.mem_424_sv2v_reg ,
  \nz.mem_423_sv2v_reg ,\nz.mem_422_sv2v_reg ,\nz.mem_421_sv2v_reg ,\nz.mem_420_sv2v_reg ,
  \nz.mem_419_sv2v_reg ,\nz.mem_418_sv2v_reg ,\nz.mem_417_sv2v_reg ,\nz.mem_416_sv2v_reg ,
  \nz.mem_415_sv2v_reg ,\nz.mem_414_sv2v_reg ,\nz.mem_413_sv2v_reg ,
  \nz.mem_412_sv2v_reg ,\nz.mem_411_sv2v_reg ,\nz.mem_410_sv2v_reg ,\nz.mem_409_sv2v_reg ,
  \nz.mem_408_sv2v_reg ,\nz.mem_407_sv2v_reg ,\nz.mem_406_sv2v_reg ,
  \nz.mem_405_sv2v_reg ,\nz.mem_404_sv2v_reg ,\nz.mem_403_sv2v_reg ,\nz.mem_402_sv2v_reg ,
  \nz.mem_401_sv2v_reg ,\nz.mem_400_sv2v_reg ,\nz.mem_399_sv2v_reg ,\nz.mem_398_sv2v_reg ,
  \nz.mem_397_sv2v_reg ,\nz.mem_396_sv2v_reg ,\nz.mem_395_sv2v_reg ,
  \nz.mem_394_sv2v_reg ,\nz.mem_393_sv2v_reg ,\nz.mem_392_sv2v_reg ,\nz.mem_391_sv2v_reg ,
  \nz.mem_390_sv2v_reg ,\nz.mem_389_sv2v_reg ,\nz.mem_388_sv2v_reg ,\nz.mem_387_sv2v_reg ,
  \nz.mem_386_sv2v_reg ,\nz.mem_385_sv2v_reg ,\nz.mem_384_sv2v_reg ,
  \nz.mem_383_sv2v_reg ,\nz.mem_382_sv2v_reg ,\nz.mem_381_sv2v_reg ,\nz.mem_380_sv2v_reg ,
  \nz.mem_379_sv2v_reg ,\nz.mem_378_sv2v_reg ,\nz.mem_377_sv2v_reg ,\nz.mem_376_sv2v_reg ,
  \nz.mem_375_sv2v_reg ,\nz.mem_374_sv2v_reg ,\nz.mem_373_sv2v_reg ,
  \nz.mem_372_sv2v_reg ,\nz.mem_371_sv2v_reg ,\nz.mem_370_sv2v_reg ,\nz.mem_369_sv2v_reg ,
  \nz.mem_368_sv2v_reg ,\nz.mem_367_sv2v_reg ,\nz.mem_366_sv2v_reg ,
  \nz.mem_365_sv2v_reg ,\nz.mem_364_sv2v_reg ,\nz.mem_363_sv2v_reg ,\nz.mem_362_sv2v_reg ,
  \nz.mem_361_sv2v_reg ,\nz.mem_360_sv2v_reg ,\nz.mem_359_sv2v_reg ,\nz.mem_358_sv2v_reg ,
  \nz.mem_357_sv2v_reg ,\nz.mem_356_sv2v_reg ,\nz.mem_355_sv2v_reg ,
  \nz.mem_354_sv2v_reg ,\nz.mem_353_sv2v_reg ,\nz.mem_352_sv2v_reg ,\nz.mem_351_sv2v_reg ,
  \nz.mem_350_sv2v_reg ,\nz.mem_349_sv2v_reg ,\nz.mem_348_sv2v_reg ,\nz.mem_347_sv2v_reg ,
  \nz.mem_346_sv2v_reg ,\nz.mem_345_sv2v_reg ,\nz.mem_344_sv2v_reg ,
  \nz.mem_343_sv2v_reg ,\nz.mem_342_sv2v_reg ,\nz.mem_341_sv2v_reg ,\nz.mem_340_sv2v_reg ,
  \nz.mem_339_sv2v_reg ,\nz.mem_338_sv2v_reg ,\nz.mem_337_sv2v_reg ,\nz.mem_336_sv2v_reg ,
  \nz.mem_335_sv2v_reg ,\nz.mem_334_sv2v_reg ,\nz.mem_333_sv2v_reg ,
  \nz.mem_332_sv2v_reg ,\nz.mem_331_sv2v_reg ,\nz.mem_330_sv2v_reg ,\nz.mem_329_sv2v_reg ,
  \nz.mem_328_sv2v_reg ,\nz.mem_327_sv2v_reg ,\nz.mem_326_sv2v_reg ,
  \nz.mem_325_sv2v_reg ,\nz.mem_324_sv2v_reg ,\nz.mem_323_sv2v_reg ,\nz.mem_322_sv2v_reg ,
  \nz.mem_321_sv2v_reg ,\nz.mem_320_sv2v_reg ,\nz.mem_319_sv2v_reg ,\nz.mem_318_sv2v_reg ,
  \nz.mem_317_sv2v_reg ,\nz.mem_316_sv2v_reg ,\nz.mem_315_sv2v_reg ,
  \nz.mem_314_sv2v_reg ,\nz.mem_313_sv2v_reg ,\nz.mem_312_sv2v_reg ,\nz.mem_311_sv2v_reg ,
  \nz.mem_310_sv2v_reg ,\nz.mem_309_sv2v_reg ,\nz.mem_308_sv2v_reg ,\nz.mem_307_sv2v_reg ,
  \nz.mem_306_sv2v_reg ,\nz.mem_305_sv2v_reg ,\nz.mem_304_sv2v_reg ,
  \nz.mem_303_sv2v_reg ,\nz.mem_302_sv2v_reg ,\nz.mem_301_sv2v_reg ,\nz.mem_300_sv2v_reg ,
  \nz.mem_299_sv2v_reg ,\nz.mem_298_sv2v_reg ,\nz.mem_297_sv2v_reg ,\nz.mem_296_sv2v_reg ,
  \nz.mem_295_sv2v_reg ,\nz.mem_294_sv2v_reg ,\nz.mem_293_sv2v_reg ,
  \nz.mem_292_sv2v_reg ,\nz.mem_291_sv2v_reg ,\nz.mem_290_sv2v_reg ,\nz.mem_289_sv2v_reg ,
  \nz.mem_288_sv2v_reg ,\nz.mem_287_sv2v_reg ,\nz.mem_286_sv2v_reg ,
  \nz.mem_285_sv2v_reg ,\nz.mem_284_sv2v_reg ,\nz.mem_283_sv2v_reg ,\nz.mem_282_sv2v_reg ,
  \nz.mem_281_sv2v_reg ,\nz.mem_280_sv2v_reg ,\nz.mem_279_sv2v_reg ,\nz.mem_278_sv2v_reg ,
  \nz.mem_277_sv2v_reg ,\nz.mem_276_sv2v_reg ,\nz.mem_275_sv2v_reg ,
  \nz.mem_274_sv2v_reg ,\nz.mem_273_sv2v_reg ,\nz.mem_272_sv2v_reg ,\nz.mem_271_sv2v_reg ,
  \nz.mem_270_sv2v_reg ,\nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,\nz.mem_267_sv2v_reg ,
  \nz.mem_266_sv2v_reg ,\nz.mem_265_sv2v_reg ,\nz.mem_264_sv2v_reg ,
  \nz.mem_263_sv2v_reg ,\nz.mem_262_sv2v_reg ,\nz.mem_261_sv2v_reg ,\nz.mem_260_sv2v_reg ,
  \nz.mem_259_sv2v_reg ,\nz.mem_258_sv2v_reg ,\nz.mem_257_sv2v_reg ,\nz.mem_256_sv2v_reg ,
  \nz.mem_255_sv2v_reg ,\nz.mem_254_sv2v_reg ,\nz.mem_253_sv2v_reg ,
  \nz.mem_252_sv2v_reg ,\nz.mem_251_sv2v_reg ,\nz.mem_250_sv2v_reg ,\nz.mem_249_sv2v_reg ,
  \nz.mem_248_sv2v_reg ,\nz.mem_247_sv2v_reg ,\nz.mem_246_sv2v_reg ,
  \nz.mem_245_sv2v_reg ,\nz.mem_244_sv2v_reg ,\nz.mem_243_sv2v_reg ,\nz.mem_242_sv2v_reg ,
  \nz.mem_241_sv2v_reg ,\nz.mem_240_sv2v_reg ,\nz.mem_239_sv2v_reg ,\nz.mem_238_sv2v_reg ,
  \nz.mem_237_sv2v_reg ,\nz.mem_236_sv2v_reg ,\nz.mem_235_sv2v_reg ,
  \nz.mem_234_sv2v_reg ,\nz.mem_233_sv2v_reg ,\nz.mem_232_sv2v_reg ,\nz.mem_231_sv2v_reg ,
  \nz.mem_230_sv2v_reg ,\nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,\nz.mem_227_sv2v_reg ,
  \nz.mem_226_sv2v_reg ,\nz.mem_225_sv2v_reg ,\nz.mem_224_sv2v_reg ,
  \nz.mem_223_sv2v_reg ,\nz.mem_222_sv2v_reg ,\nz.mem_221_sv2v_reg ,\nz.mem_220_sv2v_reg ,
  \nz.mem_219_sv2v_reg ,\nz.mem_218_sv2v_reg ,\nz.mem_217_sv2v_reg ,\nz.mem_216_sv2v_reg ,
  \nz.mem_215_sv2v_reg ,\nz.mem_214_sv2v_reg ,\nz.mem_213_sv2v_reg ,
  \nz.mem_212_sv2v_reg ,\nz.mem_211_sv2v_reg ,\nz.mem_210_sv2v_reg ,\nz.mem_209_sv2v_reg ,
  \nz.mem_208_sv2v_reg ,\nz.mem_207_sv2v_reg ,\nz.mem_206_sv2v_reg ,
  \nz.mem_205_sv2v_reg ,\nz.mem_204_sv2v_reg ,\nz.mem_203_sv2v_reg ,\nz.mem_202_sv2v_reg ,
  \nz.mem_201_sv2v_reg ,\nz.mem_200_sv2v_reg ,\nz.mem_199_sv2v_reg ,\nz.mem_198_sv2v_reg ,
  \nz.mem_197_sv2v_reg ,\nz.mem_196_sv2v_reg ,\nz.mem_195_sv2v_reg ,
  \nz.mem_194_sv2v_reg ,\nz.mem_193_sv2v_reg ,\nz.mem_192_sv2v_reg ,\nz.mem_191_sv2v_reg ,
  \nz.mem_190_sv2v_reg ,\nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,\nz.mem_187_sv2v_reg ,
  \nz.mem_186_sv2v_reg ,\nz.mem_185_sv2v_reg ,\nz.mem_184_sv2v_reg ,
  \nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,\nz.mem_181_sv2v_reg ,\nz.mem_180_sv2v_reg ,
  \nz.mem_179_sv2v_reg ,\nz.mem_178_sv2v_reg ,\nz.mem_177_sv2v_reg ,\nz.mem_176_sv2v_reg ,
  \nz.mem_175_sv2v_reg ,\nz.mem_174_sv2v_reg ,\nz.mem_173_sv2v_reg ,
  \nz.mem_172_sv2v_reg ,\nz.mem_171_sv2v_reg ,\nz.mem_170_sv2v_reg ,\nz.mem_169_sv2v_reg ,
  \nz.mem_168_sv2v_reg ,\nz.mem_167_sv2v_reg ,\nz.mem_166_sv2v_reg ,
  \nz.mem_165_sv2v_reg ,\nz.mem_164_sv2v_reg ,\nz.mem_163_sv2v_reg ,\nz.mem_162_sv2v_reg ,
  \nz.mem_161_sv2v_reg ,\nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,\nz.mem_158_sv2v_reg ,
  \nz.mem_157_sv2v_reg ,\nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,
  \nz.mem_154_sv2v_reg ,\nz.mem_153_sv2v_reg ,\nz.mem_152_sv2v_reg ,\nz.mem_151_sv2v_reg ,
  \nz.mem_150_sv2v_reg ,\nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,\nz.mem_147_sv2v_reg ,
  \nz.mem_146_sv2v_reg ,\nz.mem_145_sv2v_reg ,\nz.mem_144_sv2v_reg ,
  \nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,\nz.mem_141_sv2v_reg ,\nz.mem_140_sv2v_reg ,
  \nz.mem_139_sv2v_reg ,\nz.mem_138_sv2v_reg ,\nz.mem_137_sv2v_reg ,\nz.mem_136_sv2v_reg ,
  \nz.mem_135_sv2v_reg ,\nz.mem_134_sv2v_reg ,\nz.mem_133_sv2v_reg ,
  \nz.mem_132_sv2v_reg ,\nz.mem_131_sv2v_reg ,\nz.mem_130_sv2v_reg ,\nz.mem_129_sv2v_reg ,
  \nz.mem_128_sv2v_reg ,\nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,
  \nz.mem_125_sv2v_reg ,\nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,\nz.mem_122_sv2v_reg ,
  \nz.mem_121_sv2v_reg ,\nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,\nz.mem_118_sv2v_reg ,
  \nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,
  \nz.mem_114_sv2v_reg ,\nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,\nz.mem_111_sv2v_reg ,
  \nz.mem_110_sv2v_reg ,\nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,\nz.mem_107_sv2v_reg ,
  \nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,
  \nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,\nz.mem_100_sv2v_reg ,
  \nz.mem_99_sv2v_reg ,\nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,\nz.mem_96_sv2v_reg ,
  \nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,\nz.mem_92_sv2v_reg ,
  \nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,
  \nz.mem_88_sv2v_reg ,\nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,
  \nz.mem_84_sv2v_reg ,\nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,\nz.mem_81_sv2v_reg ,
  \nz.mem_80_sv2v_reg ,\nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,\nz.mem_77_sv2v_reg ,
  \nz.mem_76_sv2v_reg ,\nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,\nz.mem_73_sv2v_reg ,
  \nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,
  \nz.mem_69_sv2v_reg ,\nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,
  \nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,
  \nz.mem_61_sv2v_reg ,\nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,
  \nz.mem_57_sv2v_reg ,\nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,
  \nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,
  \nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,
  \nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,
  \nz.mem_42_sv2v_reg ,\nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,
  \nz.mem_38_sv2v_reg ,\nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,
  \nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,
  \nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,
  \nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,
  \nz.mem_23_sv2v_reg ,\nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,
  \nz.mem_19_sv2v_reg ,\nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,
  \nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,
  \nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,
  \nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,
  \nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,
  \nz.mem_0_sv2v_reg ;
  assign \nz.mem [455] = \nz.mem_455_sv2v_reg ;
  assign \nz.mem [454] = \nz.mem_454_sv2v_reg ;
  assign \nz.mem [453] = \nz.mem_453_sv2v_reg ;
  assign \nz.mem [452] = \nz.mem_452_sv2v_reg ;
  assign \nz.mem [451] = \nz.mem_451_sv2v_reg ;
  assign \nz.mem [450] = \nz.mem_450_sv2v_reg ;
  assign \nz.mem [449] = \nz.mem_449_sv2v_reg ;
  assign \nz.mem [448] = \nz.mem_448_sv2v_reg ;
  assign \nz.mem [447] = \nz.mem_447_sv2v_reg ;
  assign \nz.mem [446] = \nz.mem_446_sv2v_reg ;
  assign \nz.mem [445] = \nz.mem_445_sv2v_reg ;
  assign \nz.mem [444] = \nz.mem_444_sv2v_reg ;
  assign \nz.mem [443] = \nz.mem_443_sv2v_reg ;
  assign \nz.mem [442] = \nz.mem_442_sv2v_reg ;
  assign \nz.mem [441] = \nz.mem_441_sv2v_reg ;
  assign \nz.mem [440] = \nz.mem_440_sv2v_reg ;
  assign \nz.mem [439] = \nz.mem_439_sv2v_reg ;
  assign \nz.mem [438] = \nz.mem_438_sv2v_reg ;
  assign \nz.mem [437] = \nz.mem_437_sv2v_reg ;
  assign \nz.mem [436] = \nz.mem_436_sv2v_reg ;
  assign \nz.mem [435] = \nz.mem_435_sv2v_reg ;
  assign \nz.mem [434] = \nz.mem_434_sv2v_reg ;
  assign \nz.mem [433] = \nz.mem_433_sv2v_reg ;
  assign \nz.mem [432] = \nz.mem_432_sv2v_reg ;
  assign \nz.mem [431] = \nz.mem_431_sv2v_reg ;
  assign \nz.mem [430] = \nz.mem_430_sv2v_reg ;
  assign \nz.mem [429] = \nz.mem_429_sv2v_reg ;
  assign \nz.mem [428] = \nz.mem_428_sv2v_reg ;
  assign \nz.mem [427] = \nz.mem_427_sv2v_reg ;
  assign \nz.mem [426] = \nz.mem_426_sv2v_reg ;
  assign \nz.mem [425] = \nz.mem_425_sv2v_reg ;
  assign \nz.mem [424] = \nz.mem_424_sv2v_reg ;
  assign \nz.mem [423] = \nz.mem_423_sv2v_reg ;
  assign \nz.mem [422] = \nz.mem_422_sv2v_reg ;
  assign \nz.mem [421] = \nz.mem_421_sv2v_reg ;
  assign \nz.mem [420] = \nz.mem_420_sv2v_reg ;
  assign \nz.mem [419] = \nz.mem_419_sv2v_reg ;
  assign \nz.mem [418] = \nz.mem_418_sv2v_reg ;
  assign \nz.mem [417] = \nz.mem_417_sv2v_reg ;
  assign \nz.mem [416] = \nz.mem_416_sv2v_reg ;
  assign \nz.mem [415] = \nz.mem_415_sv2v_reg ;
  assign \nz.mem [414] = \nz.mem_414_sv2v_reg ;
  assign \nz.mem [413] = \nz.mem_413_sv2v_reg ;
  assign \nz.mem [412] = \nz.mem_412_sv2v_reg ;
  assign \nz.mem [411] = \nz.mem_411_sv2v_reg ;
  assign \nz.mem [410] = \nz.mem_410_sv2v_reg ;
  assign \nz.mem [409] = \nz.mem_409_sv2v_reg ;
  assign \nz.mem [408] = \nz.mem_408_sv2v_reg ;
  assign \nz.mem [407] = \nz.mem_407_sv2v_reg ;
  assign \nz.mem [406] = \nz.mem_406_sv2v_reg ;
  assign \nz.mem [405] = \nz.mem_405_sv2v_reg ;
  assign \nz.mem [404] = \nz.mem_404_sv2v_reg ;
  assign \nz.mem [403] = \nz.mem_403_sv2v_reg ;
  assign \nz.mem [402] = \nz.mem_402_sv2v_reg ;
  assign \nz.mem [401] = \nz.mem_401_sv2v_reg ;
  assign \nz.mem [400] = \nz.mem_400_sv2v_reg ;
  assign \nz.mem [399] = \nz.mem_399_sv2v_reg ;
  assign \nz.mem [398] = \nz.mem_398_sv2v_reg ;
  assign \nz.mem [397] = \nz.mem_397_sv2v_reg ;
  assign \nz.mem [396] = \nz.mem_396_sv2v_reg ;
  assign \nz.mem [395] = \nz.mem_395_sv2v_reg ;
  assign \nz.mem [394] = \nz.mem_394_sv2v_reg ;
  assign \nz.mem [393] = \nz.mem_393_sv2v_reg ;
  assign \nz.mem [392] = \nz.mem_392_sv2v_reg ;
  assign \nz.mem [391] = \nz.mem_391_sv2v_reg ;
  assign \nz.mem [390] = \nz.mem_390_sv2v_reg ;
  assign \nz.mem [389] = \nz.mem_389_sv2v_reg ;
  assign \nz.mem [388] = \nz.mem_388_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[113] = (N8)? \nz.mem [113] : 
                         (N10)? \nz.mem [227] : 
                         (N9)? \nz.mem [341] : 
                         (N11)? \nz.mem [455] : 1'b0;
  assign r_data_o[112] = (N8)? \nz.mem [112] : 
                         (N10)? \nz.mem [226] : 
                         (N9)? \nz.mem [340] : 
                         (N11)? \nz.mem [454] : 1'b0;
  assign r_data_o[111] = (N8)? \nz.mem [111] : 
                         (N10)? \nz.mem [225] : 
                         (N9)? \nz.mem [339] : 
                         (N11)? \nz.mem [453] : 1'b0;
  assign r_data_o[110] = (N8)? \nz.mem [110] : 
                         (N10)? \nz.mem [224] : 
                         (N9)? \nz.mem [338] : 
                         (N11)? \nz.mem [452] : 1'b0;
  assign r_data_o[109] = (N8)? \nz.mem [109] : 
                         (N10)? \nz.mem [223] : 
                         (N9)? \nz.mem [337] : 
                         (N11)? \nz.mem [451] : 1'b0;
  assign r_data_o[108] = (N8)? \nz.mem [108] : 
                         (N10)? \nz.mem [222] : 
                         (N9)? \nz.mem [336] : 
                         (N11)? \nz.mem [450] : 1'b0;
  assign r_data_o[107] = (N8)? \nz.mem [107] : 
                         (N10)? \nz.mem [221] : 
                         (N9)? \nz.mem [335] : 
                         (N11)? \nz.mem [449] : 1'b0;
  assign r_data_o[106] = (N8)? \nz.mem [106] : 
                         (N10)? \nz.mem [220] : 
                         (N9)? \nz.mem [334] : 
                         (N11)? \nz.mem [448] : 1'b0;
  assign r_data_o[105] = (N8)? \nz.mem [105] : 
                         (N10)? \nz.mem [219] : 
                         (N9)? \nz.mem [333] : 
                         (N11)? \nz.mem [447] : 1'b0;
  assign r_data_o[104] = (N8)? \nz.mem [104] : 
                         (N10)? \nz.mem [218] : 
                         (N9)? \nz.mem [332] : 
                         (N11)? \nz.mem [446] : 1'b0;
  assign r_data_o[103] = (N8)? \nz.mem [103] : 
                         (N10)? \nz.mem [217] : 
                         (N9)? \nz.mem [331] : 
                         (N11)? \nz.mem [445] : 1'b0;
  assign r_data_o[102] = (N8)? \nz.mem [102] : 
                         (N10)? \nz.mem [216] : 
                         (N9)? \nz.mem [330] : 
                         (N11)? \nz.mem [444] : 1'b0;
  assign r_data_o[101] = (N8)? \nz.mem [101] : 
                         (N10)? \nz.mem [215] : 
                         (N9)? \nz.mem [329] : 
                         (N11)? \nz.mem [443] : 1'b0;
  assign r_data_o[100] = (N8)? \nz.mem [100] : 
                         (N10)? \nz.mem [214] : 
                         (N9)? \nz.mem [328] : 
                         (N11)? \nz.mem [442] : 1'b0;
  assign r_data_o[99] = (N8)? \nz.mem [99] : 
                        (N10)? \nz.mem [213] : 
                        (N9)? \nz.mem [327] : 
                        (N11)? \nz.mem [441] : 1'b0;
  assign r_data_o[98] = (N8)? \nz.mem [98] : 
                        (N10)? \nz.mem [212] : 
                        (N9)? \nz.mem [326] : 
                        (N11)? \nz.mem [440] : 1'b0;
  assign r_data_o[97] = (N8)? \nz.mem [97] : 
                        (N10)? \nz.mem [211] : 
                        (N9)? \nz.mem [325] : 
                        (N11)? \nz.mem [439] : 1'b0;
  assign r_data_o[96] = (N8)? \nz.mem [96] : 
                        (N10)? \nz.mem [210] : 
                        (N9)? \nz.mem [324] : 
                        (N11)? \nz.mem [438] : 1'b0;
  assign r_data_o[95] = (N8)? \nz.mem [95] : 
                        (N10)? \nz.mem [209] : 
                        (N9)? \nz.mem [323] : 
                        (N11)? \nz.mem [437] : 1'b0;
  assign r_data_o[94] = (N8)? \nz.mem [94] : 
                        (N10)? \nz.mem [208] : 
                        (N9)? \nz.mem [322] : 
                        (N11)? \nz.mem [436] : 1'b0;
  assign r_data_o[93] = (N8)? \nz.mem [93] : 
                        (N10)? \nz.mem [207] : 
                        (N9)? \nz.mem [321] : 
                        (N11)? \nz.mem [435] : 1'b0;
  assign r_data_o[92] = (N8)? \nz.mem [92] : 
                        (N10)? \nz.mem [206] : 
                        (N9)? \nz.mem [320] : 
                        (N11)? \nz.mem [434] : 1'b0;
  assign r_data_o[91] = (N8)? \nz.mem [91] : 
                        (N10)? \nz.mem [205] : 
                        (N9)? \nz.mem [319] : 
                        (N11)? \nz.mem [433] : 1'b0;
  assign r_data_o[90] = (N8)? \nz.mem [90] : 
                        (N10)? \nz.mem [204] : 
                        (N9)? \nz.mem [318] : 
                        (N11)? \nz.mem [432] : 1'b0;
  assign r_data_o[89] = (N8)? \nz.mem [89] : 
                        (N10)? \nz.mem [203] : 
                        (N9)? \nz.mem [317] : 
                        (N11)? \nz.mem [431] : 1'b0;
  assign r_data_o[88] = (N8)? \nz.mem [88] : 
                        (N10)? \nz.mem [202] : 
                        (N9)? \nz.mem [316] : 
                        (N11)? \nz.mem [430] : 1'b0;
  assign r_data_o[87] = (N8)? \nz.mem [87] : 
                        (N10)? \nz.mem [201] : 
                        (N9)? \nz.mem [315] : 
                        (N11)? \nz.mem [429] : 1'b0;
  assign r_data_o[86] = (N8)? \nz.mem [86] : 
                        (N10)? \nz.mem [200] : 
                        (N9)? \nz.mem [314] : 
                        (N11)? \nz.mem [428] : 1'b0;
  assign r_data_o[85] = (N8)? \nz.mem [85] : 
                        (N10)? \nz.mem [199] : 
                        (N9)? \nz.mem [313] : 
                        (N11)? \nz.mem [427] : 1'b0;
  assign r_data_o[84] = (N8)? \nz.mem [84] : 
                        (N10)? \nz.mem [198] : 
                        (N9)? \nz.mem [312] : 
                        (N11)? \nz.mem [426] : 1'b0;
  assign r_data_o[83] = (N8)? \nz.mem [83] : 
                        (N10)? \nz.mem [197] : 
                        (N9)? \nz.mem [311] : 
                        (N11)? \nz.mem [425] : 1'b0;
  assign r_data_o[82] = (N8)? \nz.mem [82] : 
                        (N10)? \nz.mem [196] : 
                        (N9)? \nz.mem [310] : 
                        (N11)? \nz.mem [424] : 1'b0;
  assign r_data_o[81] = (N8)? \nz.mem [81] : 
                        (N10)? \nz.mem [195] : 
                        (N9)? \nz.mem [309] : 
                        (N11)? \nz.mem [423] : 1'b0;
  assign r_data_o[80] = (N8)? \nz.mem [80] : 
                        (N10)? \nz.mem [194] : 
                        (N9)? \nz.mem [308] : 
                        (N11)? \nz.mem [422] : 1'b0;
  assign r_data_o[79] = (N8)? \nz.mem [79] : 
                        (N10)? \nz.mem [193] : 
                        (N9)? \nz.mem [307] : 
                        (N11)? \nz.mem [421] : 1'b0;
  assign r_data_o[78] = (N8)? \nz.mem [78] : 
                        (N10)? \nz.mem [192] : 
                        (N9)? \nz.mem [306] : 
                        (N11)? \nz.mem [420] : 1'b0;
  assign r_data_o[77] = (N8)? \nz.mem [77] : 
                        (N10)? \nz.mem [191] : 
                        (N9)? \nz.mem [305] : 
                        (N11)? \nz.mem [419] : 1'b0;
  assign r_data_o[76] = (N8)? \nz.mem [76] : 
                        (N10)? \nz.mem [190] : 
                        (N9)? \nz.mem [304] : 
                        (N11)? \nz.mem [418] : 1'b0;
  assign r_data_o[75] = (N8)? \nz.mem [75] : 
                        (N10)? \nz.mem [189] : 
                        (N9)? \nz.mem [303] : 
                        (N11)? \nz.mem [417] : 1'b0;
  assign r_data_o[74] = (N8)? \nz.mem [74] : 
                        (N10)? \nz.mem [188] : 
                        (N9)? \nz.mem [302] : 
                        (N11)? \nz.mem [416] : 1'b0;
  assign r_data_o[73] = (N8)? \nz.mem [73] : 
                        (N10)? \nz.mem [187] : 
                        (N9)? \nz.mem [301] : 
                        (N11)? \nz.mem [415] : 1'b0;
  assign r_data_o[72] = (N8)? \nz.mem [72] : 
                        (N10)? \nz.mem [186] : 
                        (N9)? \nz.mem [300] : 
                        (N11)? \nz.mem [414] : 1'b0;
  assign r_data_o[71] = (N8)? \nz.mem [71] : 
                        (N10)? \nz.mem [185] : 
                        (N9)? \nz.mem [299] : 
                        (N11)? \nz.mem [413] : 1'b0;
  assign r_data_o[70] = (N8)? \nz.mem [70] : 
                        (N10)? \nz.mem [184] : 
                        (N9)? \nz.mem [298] : 
                        (N11)? \nz.mem [412] : 1'b0;
  assign r_data_o[69] = (N8)? \nz.mem [69] : 
                        (N10)? \nz.mem [183] : 
                        (N9)? \nz.mem [297] : 
                        (N11)? \nz.mem [411] : 1'b0;
  assign r_data_o[68] = (N8)? \nz.mem [68] : 
                        (N10)? \nz.mem [182] : 
                        (N9)? \nz.mem [296] : 
                        (N11)? \nz.mem [410] : 1'b0;
  assign r_data_o[67] = (N8)? \nz.mem [67] : 
                        (N10)? \nz.mem [181] : 
                        (N9)? \nz.mem [295] : 
                        (N11)? \nz.mem [409] : 1'b0;
  assign r_data_o[66] = (N8)? \nz.mem [66] : 
                        (N10)? \nz.mem [180] : 
                        (N9)? \nz.mem [294] : 
                        (N11)? \nz.mem [408] : 1'b0;
  assign r_data_o[65] = (N8)? \nz.mem [65] : 
                        (N10)? \nz.mem [179] : 
                        (N9)? \nz.mem [293] : 
                        (N11)? \nz.mem [407] : 1'b0;
  assign r_data_o[64] = (N8)? \nz.mem [64] : 
                        (N10)? \nz.mem [178] : 
                        (N9)? \nz.mem [292] : 
                        (N11)? \nz.mem [406] : 1'b0;
  assign r_data_o[63] = (N8)? \nz.mem [63] : 
                        (N10)? \nz.mem [177] : 
                        (N9)? \nz.mem [291] : 
                        (N11)? \nz.mem [405] : 1'b0;
  assign r_data_o[62] = (N8)? \nz.mem [62] : 
                        (N10)? \nz.mem [176] : 
                        (N9)? \nz.mem [290] : 
                        (N11)? \nz.mem [404] : 1'b0;
  assign r_data_o[61] = (N8)? \nz.mem [61] : 
                        (N10)? \nz.mem [175] : 
                        (N9)? \nz.mem [289] : 
                        (N11)? \nz.mem [403] : 1'b0;
  assign r_data_o[60] = (N8)? \nz.mem [60] : 
                        (N10)? \nz.mem [174] : 
                        (N9)? \nz.mem [288] : 
                        (N11)? \nz.mem [402] : 1'b0;
  assign r_data_o[59] = (N8)? \nz.mem [59] : 
                        (N10)? \nz.mem [173] : 
                        (N9)? \nz.mem [287] : 
                        (N11)? \nz.mem [401] : 1'b0;
  assign r_data_o[58] = (N8)? \nz.mem [58] : 
                        (N10)? \nz.mem [172] : 
                        (N9)? \nz.mem [286] : 
                        (N11)? \nz.mem [400] : 1'b0;
  assign r_data_o[57] = (N8)? \nz.mem [57] : 
                        (N10)? \nz.mem [171] : 
                        (N9)? \nz.mem [285] : 
                        (N11)? \nz.mem [399] : 1'b0;
  assign r_data_o[56] = (N8)? \nz.mem [56] : 
                        (N10)? \nz.mem [170] : 
                        (N9)? \nz.mem [284] : 
                        (N11)? \nz.mem [398] : 1'b0;
  assign r_data_o[55] = (N8)? \nz.mem [55] : 
                        (N10)? \nz.mem [169] : 
                        (N9)? \nz.mem [283] : 
                        (N11)? \nz.mem [397] : 1'b0;
  assign r_data_o[54] = (N8)? \nz.mem [54] : 
                        (N10)? \nz.mem [168] : 
                        (N9)? \nz.mem [282] : 
                        (N11)? \nz.mem [396] : 1'b0;
  assign r_data_o[53] = (N8)? \nz.mem [53] : 
                        (N10)? \nz.mem [167] : 
                        (N9)? \nz.mem [281] : 
                        (N11)? \nz.mem [395] : 1'b0;
  assign r_data_o[52] = (N8)? \nz.mem [52] : 
                        (N10)? \nz.mem [166] : 
                        (N9)? \nz.mem [280] : 
                        (N11)? \nz.mem [394] : 1'b0;
  assign r_data_o[51] = (N8)? \nz.mem [51] : 
                        (N10)? \nz.mem [165] : 
                        (N9)? \nz.mem [279] : 
                        (N11)? \nz.mem [393] : 1'b0;
  assign r_data_o[50] = (N8)? \nz.mem [50] : 
                        (N10)? \nz.mem [164] : 
                        (N9)? \nz.mem [278] : 
                        (N11)? \nz.mem [392] : 1'b0;
  assign r_data_o[49] = (N8)? \nz.mem [49] : 
                        (N10)? \nz.mem [163] : 
                        (N9)? \nz.mem [277] : 
                        (N11)? \nz.mem [391] : 1'b0;
  assign r_data_o[48] = (N8)? \nz.mem [48] : 
                        (N10)? \nz.mem [162] : 
                        (N9)? \nz.mem [276] : 
                        (N11)? \nz.mem [390] : 1'b0;
  assign r_data_o[47] = (N8)? \nz.mem [47] : 
                        (N10)? \nz.mem [161] : 
                        (N9)? \nz.mem [275] : 
                        (N11)? \nz.mem [389] : 1'b0;
  assign r_data_o[46] = (N8)? \nz.mem [46] : 
                        (N10)? \nz.mem [160] : 
                        (N9)? \nz.mem [274] : 
                        (N11)? \nz.mem [388] : 1'b0;
  assign r_data_o[45] = (N8)? \nz.mem [45] : 
                        (N10)? \nz.mem [159] : 
                        (N9)? \nz.mem [273] : 
                        (N11)? \nz.mem [387] : 1'b0;
  assign r_data_o[44] = (N8)? \nz.mem [44] : 
                        (N10)? \nz.mem [158] : 
                        (N9)? \nz.mem [272] : 
                        (N11)? \nz.mem [386] : 1'b0;
  assign r_data_o[43] = (N8)? \nz.mem [43] : 
                        (N10)? \nz.mem [157] : 
                        (N9)? \nz.mem [271] : 
                        (N11)? \nz.mem [385] : 1'b0;
  assign r_data_o[42] = (N8)? \nz.mem [42] : 
                        (N10)? \nz.mem [156] : 
                        (N9)? \nz.mem [270] : 
                        (N11)? \nz.mem [384] : 1'b0;
  assign r_data_o[41] = (N8)? \nz.mem [41] : 
                        (N10)? \nz.mem [155] : 
                        (N9)? \nz.mem [269] : 
                        (N11)? \nz.mem [383] : 1'b0;
  assign r_data_o[40] = (N8)? \nz.mem [40] : 
                        (N10)? \nz.mem [154] : 
                        (N9)? \nz.mem [268] : 
                        (N11)? \nz.mem [382] : 1'b0;
  assign r_data_o[39] = (N8)? \nz.mem [39] : 
                        (N10)? \nz.mem [153] : 
                        (N9)? \nz.mem [267] : 
                        (N11)? \nz.mem [381] : 1'b0;
  assign r_data_o[38] = (N8)? \nz.mem [38] : 
                        (N10)? \nz.mem [152] : 
                        (N9)? \nz.mem [266] : 
                        (N11)? \nz.mem [380] : 1'b0;
  assign r_data_o[37] = (N8)? \nz.mem [37] : 
                        (N10)? \nz.mem [151] : 
                        (N9)? \nz.mem [265] : 
                        (N11)? \nz.mem [379] : 1'b0;
  assign r_data_o[36] = (N8)? \nz.mem [36] : 
                        (N10)? \nz.mem [150] : 
                        (N9)? \nz.mem [264] : 
                        (N11)? \nz.mem [378] : 1'b0;
  assign r_data_o[35] = (N8)? \nz.mem [35] : 
                        (N10)? \nz.mem [149] : 
                        (N9)? \nz.mem [263] : 
                        (N11)? \nz.mem [377] : 1'b0;
  assign r_data_o[34] = (N8)? \nz.mem [34] : 
                        (N10)? \nz.mem [148] : 
                        (N9)? \nz.mem [262] : 
                        (N11)? \nz.mem [376] : 1'b0;
  assign r_data_o[33] = (N8)? \nz.mem [33] : 
                        (N10)? \nz.mem [147] : 
                        (N9)? \nz.mem [261] : 
                        (N11)? \nz.mem [375] : 1'b0;
  assign r_data_o[32] = (N8)? \nz.mem [32] : 
                        (N10)? \nz.mem [146] : 
                        (N9)? \nz.mem [260] : 
                        (N11)? \nz.mem [374] : 1'b0;
  assign r_data_o[31] = (N8)? \nz.mem [31] : 
                        (N10)? \nz.mem [145] : 
                        (N9)? \nz.mem [259] : 
                        (N11)? \nz.mem [373] : 1'b0;
  assign r_data_o[30] = (N8)? \nz.mem [30] : 
                        (N10)? \nz.mem [144] : 
                        (N9)? \nz.mem [258] : 
                        (N11)? \nz.mem [372] : 1'b0;
  assign r_data_o[29] = (N8)? \nz.mem [29] : 
                        (N10)? \nz.mem [143] : 
                        (N9)? \nz.mem [257] : 
                        (N11)? \nz.mem [371] : 1'b0;
  assign r_data_o[28] = (N8)? \nz.mem [28] : 
                        (N10)? \nz.mem [142] : 
                        (N9)? \nz.mem [256] : 
                        (N11)? \nz.mem [370] : 1'b0;
  assign r_data_o[27] = (N8)? \nz.mem [27] : 
                        (N10)? \nz.mem [141] : 
                        (N9)? \nz.mem [255] : 
                        (N11)? \nz.mem [369] : 1'b0;
  assign r_data_o[26] = (N8)? \nz.mem [26] : 
                        (N10)? \nz.mem [140] : 
                        (N9)? \nz.mem [254] : 
                        (N11)? \nz.mem [368] : 1'b0;
  assign r_data_o[25] = (N8)? \nz.mem [25] : 
                        (N10)? \nz.mem [139] : 
                        (N9)? \nz.mem [253] : 
                        (N11)? \nz.mem [367] : 1'b0;
  assign r_data_o[24] = (N8)? \nz.mem [24] : 
                        (N10)? \nz.mem [138] : 
                        (N9)? \nz.mem [252] : 
                        (N11)? \nz.mem [366] : 1'b0;
  assign r_data_o[23] = (N8)? \nz.mem [23] : 
                        (N10)? \nz.mem [137] : 
                        (N9)? \nz.mem [251] : 
                        (N11)? \nz.mem [365] : 1'b0;
  assign r_data_o[22] = (N8)? \nz.mem [22] : 
                        (N10)? \nz.mem [136] : 
                        (N9)? \nz.mem [250] : 
                        (N11)? \nz.mem [364] : 1'b0;
  assign r_data_o[21] = (N8)? \nz.mem [21] : 
                        (N10)? \nz.mem [135] : 
                        (N9)? \nz.mem [249] : 
                        (N11)? \nz.mem [363] : 1'b0;
  assign r_data_o[20] = (N8)? \nz.mem [20] : 
                        (N10)? \nz.mem [134] : 
                        (N9)? \nz.mem [248] : 
                        (N11)? \nz.mem [362] : 1'b0;
  assign r_data_o[19] = (N8)? \nz.mem [19] : 
                        (N10)? \nz.mem [133] : 
                        (N9)? \nz.mem [247] : 
                        (N11)? \nz.mem [361] : 1'b0;
  assign r_data_o[18] = (N8)? \nz.mem [18] : 
                        (N10)? \nz.mem [132] : 
                        (N9)? \nz.mem [246] : 
                        (N11)? \nz.mem [360] : 1'b0;
  assign r_data_o[17] = (N8)? \nz.mem [17] : 
                        (N10)? \nz.mem [131] : 
                        (N9)? \nz.mem [245] : 
                        (N11)? \nz.mem [359] : 1'b0;
  assign r_data_o[16] = (N8)? \nz.mem [16] : 
                        (N10)? \nz.mem [130] : 
                        (N9)? \nz.mem [244] : 
                        (N11)? \nz.mem [358] : 1'b0;
  assign r_data_o[15] = (N8)? \nz.mem [15] : 
                        (N10)? \nz.mem [129] : 
                        (N9)? \nz.mem [243] : 
                        (N11)? \nz.mem [357] : 1'b0;
  assign r_data_o[14] = (N8)? \nz.mem [14] : 
                        (N10)? \nz.mem [128] : 
                        (N9)? \nz.mem [242] : 
                        (N11)? \nz.mem [356] : 1'b0;
  assign r_data_o[13] = (N8)? \nz.mem [13] : 
                        (N10)? \nz.mem [127] : 
                        (N9)? \nz.mem [241] : 
                        (N11)? \nz.mem [355] : 1'b0;
  assign r_data_o[12] = (N8)? \nz.mem [12] : 
                        (N10)? \nz.mem [126] : 
                        (N9)? \nz.mem [240] : 
                        (N11)? \nz.mem [354] : 1'b0;
  assign r_data_o[11] = (N8)? \nz.mem [11] : 
                        (N10)? \nz.mem [125] : 
                        (N9)? \nz.mem [239] : 
                        (N11)? \nz.mem [353] : 1'b0;
  assign r_data_o[10] = (N8)? \nz.mem [10] : 
                        (N10)? \nz.mem [124] : 
                        (N9)? \nz.mem [238] : 
                        (N11)? \nz.mem [352] : 1'b0;
  assign r_data_o[9] = (N8)? \nz.mem [9] : 
                       (N10)? \nz.mem [123] : 
                       (N9)? \nz.mem [237] : 
                       (N11)? \nz.mem [351] : 1'b0;
  assign r_data_o[8] = (N8)? \nz.mem [8] : 
                       (N10)? \nz.mem [122] : 
                       (N9)? \nz.mem [236] : 
                       (N11)? \nz.mem [350] : 1'b0;
  assign r_data_o[7] = (N8)? \nz.mem [7] : 
                       (N10)? \nz.mem [121] : 
                       (N9)? \nz.mem [235] : 
                       (N11)? \nz.mem [349] : 1'b0;
  assign r_data_o[6] = (N8)? \nz.mem [6] : 
                       (N10)? \nz.mem [120] : 
                       (N9)? \nz.mem [234] : 
                       (N11)? \nz.mem [348] : 1'b0;
  assign r_data_o[5] = (N8)? \nz.mem [5] : 
                       (N10)? \nz.mem [119] : 
                       (N9)? \nz.mem [233] : 
                       (N11)? \nz.mem [347] : 1'b0;
  assign r_data_o[4] = (N8)? \nz.mem [4] : 
                       (N10)? \nz.mem [118] : 
                       (N9)? \nz.mem [232] : 
                       (N11)? \nz.mem [346] : 1'b0;
  assign r_data_o[3] = (N8)? \nz.mem [3] : 
                       (N10)? \nz.mem [117] : 
                       (N9)? \nz.mem [231] : 
                       (N11)? \nz.mem [345] : 1'b0;
  assign r_data_o[2] = (N8)? \nz.mem [2] : 
                       (N10)? \nz.mem [116] : 
                       (N9)? \nz.mem [230] : 
                       (N11)? \nz.mem [344] : 1'b0;
  assign r_data_o[1] = (N8)? \nz.mem [1] : 
                       (N10)? \nz.mem [115] : 
                       (N9)? \nz.mem [229] : 
                       (N11)? \nz.mem [343] : 1'b0;
  assign r_data_o[0] = (N8)? \nz.mem [0] : 
                       (N10)? \nz.mem [114] : 
                       (N9)? \nz.mem [228] : 
                       (N11)? \nz.mem [342] : 1'b0;
  assign N16 = w_addr_i[0] & w_addr_i[1];
  assign N15 = N0 & w_addr_i[1];
  assign N0 = ~w_addr_i[0];
  assign N14 = w_addr_i[0] & N1;
  assign N1 = ~w_addr_i[1];
  assign N13 = N2 & N3;
  assign N2 = ~w_addr_i[0];
  assign N3 = ~w_addr_i[1];
  assign { N24, N23, N22, N21, N20, N19, N18, N17 } = (N4)? { N16, N16, N15, N15, N14, N14, N13, N13 } : 
                                                      (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N4 = w_v_i;
  assign N5 = N12;
  assign N6 = ~r_addr_i[0];
  assign N7 = ~r_addr_i[1];
  assign N8 = N6 & N7;
  assign N9 = N6 & r_addr_i[1];
  assign N10 = r_addr_i[0] & N7;
  assign N11 = r_addr_i[0] & r_addr_i[1];
  assign N12 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N23) begin
      \nz.mem_455_sv2v_reg  <= w_data_i[113];
      \nz.mem_454_sv2v_reg  <= w_data_i[112];
      \nz.mem_453_sv2v_reg  <= w_data_i[111];
      \nz.mem_452_sv2v_reg  <= w_data_i[110];
      \nz.mem_451_sv2v_reg  <= w_data_i[109];
      \nz.mem_450_sv2v_reg  <= w_data_i[108];
      \nz.mem_449_sv2v_reg  <= w_data_i[107];
      \nz.mem_448_sv2v_reg  <= w_data_i[106];
      \nz.mem_447_sv2v_reg  <= w_data_i[105];
      \nz.mem_446_sv2v_reg  <= w_data_i[104];
      \nz.mem_445_sv2v_reg  <= w_data_i[103];
      \nz.mem_444_sv2v_reg  <= w_data_i[102];
      \nz.mem_443_sv2v_reg  <= w_data_i[101];
      \nz.mem_442_sv2v_reg  <= w_data_i[100];
      \nz.mem_441_sv2v_reg  <= w_data_i[99];
      \nz.mem_440_sv2v_reg  <= w_data_i[98];
      \nz.mem_439_sv2v_reg  <= w_data_i[97];
      \nz.mem_438_sv2v_reg  <= w_data_i[96];
      \nz.mem_437_sv2v_reg  <= w_data_i[95];
      \nz.mem_436_sv2v_reg  <= w_data_i[94];
      \nz.mem_435_sv2v_reg  <= w_data_i[93];
      \nz.mem_434_sv2v_reg  <= w_data_i[92];
      \nz.mem_433_sv2v_reg  <= w_data_i[91];
      \nz.mem_432_sv2v_reg  <= w_data_i[90];
      \nz.mem_431_sv2v_reg  <= w_data_i[89];
      \nz.mem_430_sv2v_reg  <= w_data_i[88];
      \nz.mem_429_sv2v_reg  <= w_data_i[87];
      \nz.mem_428_sv2v_reg  <= w_data_i[86];
      \nz.mem_427_sv2v_reg  <= w_data_i[85];
      \nz.mem_426_sv2v_reg  <= w_data_i[84];
      \nz.mem_425_sv2v_reg  <= w_data_i[83];
      \nz.mem_424_sv2v_reg  <= w_data_i[82];
      \nz.mem_423_sv2v_reg  <= w_data_i[81];
      \nz.mem_422_sv2v_reg  <= w_data_i[80];
      \nz.mem_421_sv2v_reg  <= w_data_i[79];
      \nz.mem_420_sv2v_reg  <= w_data_i[78];
      \nz.mem_419_sv2v_reg  <= w_data_i[77];
      \nz.mem_418_sv2v_reg  <= w_data_i[76];
      \nz.mem_417_sv2v_reg  <= w_data_i[75];
      \nz.mem_416_sv2v_reg  <= w_data_i[74];
      \nz.mem_415_sv2v_reg  <= w_data_i[73];
      \nz.mem_414_sv2v_reg  <= w_data_i[72];
      \nz.mem_413_sv2v_reg  <= w_data_i[71];
      \nz.mem_412_sv2v_reg  <= w_data_i[70];
      \nz.mem_411_sv2v_reg  <= w_data_i[69];
      \nz.mem_410_sv2v_reg  <= w_data_i[68];
      \nz.mem_409_sv2v_reg  <= w_data_i[67];
      \nz.mem_408_sv2v_reg  <= w_data_i[66];
      \nz.mem_407_sv2v_reg  <= w_data_i[65];
      \nz.mem_406_sv2v_reg  <= w_data_i[64];
      \nz.mem_405_sv2v_reg  <= w_data_i[63];
      \nz.mem_404_sv2v_reg  <= w_data_i[62];
      \nz.mem_403_sv2v_reg  <= w_data_i[61];
      \nz.mem_402_sv2v_reg  <= w_data_i[60];
      \nz.mem_401_sv2v_reg  <= w_data_i[59];
      \nz.mem_400_sv2v_reg  <= w_data_i[58];
      \nz.mem_399_sv2v_reg  <= w_data_i[57];
      \nz.mem_398_sv2v_reg  <= w_data_i[56];
      \nz.mem_397_sv2v_reg  <= w_data_i[55];
      \nz.mem_396_sv2v_reg  <= w_data_i[54];
      \nz.mem_395_sv2v_reg  <= w_data_i[53];
      \nz.mem_394_sv2v_reg  <= w_data_i[52];
      \nz.mem_393_sv2v_reg  <= w_data_i[51];
      \nz.mem_392_sv2v_reg  <= w_data_i[50];
      \nz.mem_391_sv2v_reg  <= w_data_i[49];
      \nz.mem_390_sv2v_reg  <= w_data_i[48];
      \nz.mem_389_sv2v_reg  <= w_data_i[47];
      \nz.mem_388_sv2v_reg  <= w_data_i[46];
      \nz.mem_387_sv2v_reg  <= w_data_i[45];
      \nz.mem_386_sv2v_reg  <= w_data_i[44];
      \nz.mem_385_sv2v_reg  <= w_data_i[43];
      \nz.mem_384_sv2v_reg  <= w_data_i[42];
      \nz.mem_383_sv2v_reg  <= w_data_i[41];
      \nz.mem_382_sv2v_reg  <= w_data_i[40];
      \nz.mem_381_sv2v_reg  <= w_data_i[39];
      \nz.mem_380_sv2v_reg  <= w_data_i[38];
      \nz.mem_379_sv2v_reg  <= w_data_i[37];
      \nz.mem_378_sv2v_reg  <= w_data_i[36];
      \nz.mem_377_sv2v_reg  <= w_data_i[35];
      \nz.mem_376_sv2v_reg  <= w_data_i[34];
      \nz.mem_375_sv2v_reg  <= w_data_i[33];
      \nz.mem_374_sv2v_reg  <= w_data_i[32];
      \nz.mem_373_sv2v_reg  <= w_data_i[31];
      \nz.mem_372_sv2v_reg  <= w_data_i[30];
      \nz.mem_371_sv2v_reg  <= w_data_i[29];
      \nz.mem_370_sv2v_reg  <= w_data_i[28];
      \nz.mem_369_sv2v_reg  <= w_data_i[27];
      \nz.mem_368_sv2v_reg  <= w_data_i[26];
      \nz.mem_367_sv2v_reg  <= w_data_i[25];
      \nz.mem_366_sv2v_reg  <= w_data_i[24];
      \nz.mem_365_sv2v_reg  <= w_data_i[23];
      \nz.mem_364_sv2v_reg  <= w_data_i[22];
      \nz.mem_363_sv2v_reg  <= w_data_i[21];
      \nz.mem_362_sv2v_reg  <= w_data_i[20];
      \nz.mem_361_sv2v_reg  <= w_data_i[19];
      \nz.mem_360_sv2v_reg  <= w_data_i[18];
      \nz.mem_359_sv2v_reg  <= w_data_i[17];
      \nz.mem_358_sv2v_reg  <= w_data_i[16];
      \nz.mem_357_sv2v_reg  <= w_data_i[15];
      \nz.mem_342_sv2v_reg  <= w_data_i[0];
    end 
    if(N24) begin
      \nz.mem_356_sv2v_reg  <= w_data_i[14];
      \nz.mem_355_sv2v_reg  <= w_data_i[13];
      \nz.mem_354_sv2v_reg  <= w_data_i[12];
      \nz.mem_353_sv2v_reg  <= w_data_i[11];
      \nz.mem_352_sv2v_reg  <= w_data_i[10];
      \nz.mem_351_sv2v_reg  <= w_data_i[9];
      \nz.mem_350_sv2v_reg  <= w_data_i[8];
      \nz.mem_349_sv2v_reg  <= w_data_i[7];
      \nz.mem_348_sv2v_reg  <= w_data_i[6];
      \nz.mem_347_sv2v_reg  <= w_data_i[5];
      \nz.mem_346_sv2v_reg  <= w_data_i[4];
      \nz.mem_345_sv2v_reg  <= w_data_i[3];
      \nz.mem_344_sv2v_reg  <= w_data_i[2];
      \nz.mem_343_sv2v_reg  <= w_data_i[1];
    end 
    if(N21) begin
      \nz.mem_341_sv2v_reg  <= w_data_i[113];
      \nz.mem_340_sv2v_reg  <= w_data_i[112];
      \nz.mem_339_sv2v_reg  <= w_data_i[111];
      \nz.mem_338_sv2v_reg  <= w_data_i[110];
      \nz.mem_337_sv2v_reg  <= w_data_i[109];
      \nz.mem_336_sv2v_reg  <= w_data_i[108];
      \nz.mem_335_sv2v_reg  <= w_data_i[107];
      \nz.mem_334_sv2v_reg  <= w_data_i[106];
      \nz.mem_333_sv2v_reg  <= w_data_i[105];
      \nz.mem_332_sv2v_reg  <= w_data_i[104];
      \nz.mem_331_sv2v_reg  <= w_data_i[103];
      \nz.mem_330_sv2v_reg  <= w_data_i[102];
      \nz.mem_329_sv2v_reg  <= w_data_i[101];
      \nz.mem_328_sv2v_reg  <= w_data_i[100];
      \nz.mem_327_sv2v_reg  <= w_data_i[99];
      \nz.mem_326_sv2v_reg  <= w_data_i[98];
      \nz.mem_325_sv2v_reg  <= w_data_i[97];
      \nz.mem_324_sv2v_reg  <= w_data_i[96];
      \nz.mem_323_sv2v_reg  <= w_data_i[95];
      \nz.mem_322_sv2v_reg  <= w_data_i[94];
      \nz.mem_321_sv2v_reg  <= w_data_i[93];
      \nz.mem_320_sv2v_reg  <= w_data_i[92];
      \nz.mem_319_sv2v_reg  <= w_data_i[91];
      \nz.mem_318_sv2v_reg  <= w_data_i[90];
      \nz.mem_317_sv2v_reg  <= w_data_i[89];
      \nz.mem_316_sv2v_reg  <= w_data_i[88];
      \nz.mem_315_sv2v_reg  <= w_data_i[87];
      \nz.mem_314_sv2v_reg  <= w_data_i[86];
      \nz.mem_313_sv2v_reg  <= w_data_i[85];
      \nz.mem_312_sv2v_reg  <= w_data_i[84];
      \nz.mem_311_sv2v_reg  <= w_data_i[83];
      \nz.mem_310_sv2v_reg  <= w_data_i[82];
      \nz.mem_309_sv2v_reg  <= w_data_i[81];
      \nz.mem_308_sv2v_reg  <= w_data_i[80];
      \nz.mem_307_sv2v_reg  <= w_data_i[79];
      \nz.mem_306_sv2v_reg  <= w_data_i[78];
      \nz.mem_305_sv2v_reg  <= w_data_i[77];
      \nz.mem_304_sv2v_reg  <= w_data_i[76];
      \nz.mem_303_sv2v_reg  <= w_data_i[75];
      \nz.mem_302_sv2v_reg  <= w_data_i[74];
      \nz.mem_301_sv2v_reg  <= w_data_i[73];
      \nz.mem_300_sv2v_reg  <= w_data_i[72];
      \nz.mem_299_sv2v_reg  <= w_data_i[71];
      \nz.mem_298_sv2v_reg  <= w_data_i[70];
      \nz.mem_297_sv2v_reg  <= w_data_i[69];
      \nz.mem_296_sv2v_reg  <= w_data_i[68];
      \nz.mem_295_sv2v_reg  <= w_data_i[67];
      \nz.mem_294_sv2v_reg  <= w_data_i[66];
      \nz.mem_293_sv2v_reg  <= w_data_i[65];
      \nz.mem_292_sv2v_reg  <= w_data_i[64];
      \nz.mem_291_sv2v_reg  <= w_data_i[63];
      \nz.mem_290_sv2v_reg  <= w_data_i[62];
      \nz.mem_289_sv2v_reg  <= w_data_i[61];
      \nz.mem_288_sv2v_reg  <= w_data_i[60];
      \nz.mem_287_sv2v_reg  <= w_data_i[59];
      \nz.mem_286_sv2v_reg  <= w_data_i[58];
      \nz.mem_285_sv2v_reg  <= w_data_i[57];
      \nz.mem_284_sv2v_reg  <= w_data_i[56];
      \nz.mem_283_sv2v_reg  <= w_data_i[55];
      \nz.mem_282_sv2v_reg  <= w_data_i[54];
      \nz.mem_281_sv2v_reg  <= w_data_i[53];
      \nz.mem_280_sv2v_reg  <= w_data_i[52];
      \nz.mem_279_sv2v_reg  <= w_data_i[51];
      \nz.mem_278_sv2v_reg  <= w_data_i[50];
      \nz.mem_277_sv2v_reg  <= w_data_i[49];
      \nz.mem_276_sv2v_reg  <= w_data_i[48];
      \nz.mem_275_sv2v_reg  <= w_data_i[47];
      \nz.mem_274_sv2v_reg  <= w_data_i[46];
      \nz.mem_273_sv2v_reg  <= w_data_i[45];
      \nz.mem_272_sv2v_reg  <= w_data_i[44];
      \nz.mem_271_sv2v_reg  <= w_data_i[43];
      \nz.mem_270_sv2v_reg  <= w_data_i[42];
      \nz.mem_269_sv2v_reg  <= w_data_i[41];
      \nz.mem_268_sv2v_reg  <= w_data_i[40];
      \nz.mem_267_sv2v_reg  <= w_data_i[39];
      \nz.mem_266_sv2v_reg  <= w_data_i[38];
      \nz.mem_265_sv2v_reg  <= w_data_i[37];
      \nz.mem_264_sv2v_reg  <= w_data_i[36];
      \nz.mem_263_sv2v_reg  <= w_data_i[35];
      \nz.mem_262_sv2v_reg  <= w_data_i[34];
      \nz.mem_261_sv2v_reg  <= w_data_i[33];
      \nz.mem_260_sv2v_reg  <= w_data_i[32];
      \nz.mem_259_sv2v_reg  <= w_data_i[31];
      \nz.mem_258_sv2v_reg  <= w_data_i[30];
      \nz.mem_257_sv2v_reg  <= w_data_i[29];
      \nz.mem_256_sv2v_reg  <= w_data_i[28];
      \nz.mem_255_sv2v_reg  <= w_data_i[27];
      \nz.mem_254_sv2v_reg  <= w_data_i[26];
      \nz.mem_253_sv2v_reg  <= w_data_i[25];
      \nz.mem_252_sv2v_reg  <= w_data_i[24];
      \nz.mem_251_sv2v_reg  <= w_data_i[23];
      \nz.mem_250_sv2v_reg  <= w_data_i[22];
      \nz.mem_249_sv2v_reg  <= w_data_i[21];
      \nz.mem_248_sv2v_reg  <= w_data_i[20];
      \nz.mem_247_sv2v_reg  <= w_data_i[19];
      \nz.mem_246_sv2v_reg  <= w_data_i[18];
      \nz.mem_245_sv2v_reg  <= w_data_i[17];
      \nz.mem_244_sv2v_reg  <= w_data_i[16];
      \nz.mem_243_sv2v_reg  <= w_data_i[15];
      \nz.mem_228_sv2v_reg  <= w_data_i[0];
    end 
    if(N22) begin
      \nz.mem_242_sv2v_reg  <= w_data_i[14];
      \nz.mem_241_sv2v_reg  <= w_data_i[13];
      \nz.mem_240_sv2v_reg  <= w_data_i[12];
      \nz.mem_239_sv2v_reg  <= w_data_i[11];
      \nz.mem_238_sv2v_reg  <= w_data_i[10];
      \nz.mem_237_sv2v_reg  <= w_data_i[9];
      \nz.mem_236_sv2v_reg  <= w_data_i[8];
      \nz.mem_235_sv2v_reg  <= w_data_i[7];
      \nz.mem_234_sv2v_reg  <= w_data_i[6];
      \nz.mem_233_sv2v_reg  <= w_data_i[5];
      \nz.mem_232_sv2v_reg  <= w_data_i[4];
      \nz.mem_231_sv2v_reg  <= w_data_i[3];
      \nz.mem_230_sv2v_reg  <= w_data_i[2];
      \nz.mem_229_sv2v_reg  <= w_data_i[1];
    end 
    if(N19) begin
      \nz.mem_227_sv2v_reg  <= w_data_i[113];
      \nz.mem_226_sv2v_reg  <= w_data_i[112];
      \nz.mem_225_sv2v_reg  <= w_data_i[111];
      \nz.mem_224_sv2v_reg  <= w_data_i[110];
      \nz.mem_223_sv2v_reg  <= w_data_i[109];
      \nz.mem_222_sv2v_reg  <= w_data_i[108];
      \nz.mem_221_sv2v_reg  <= w_data_i[107];
      \nz.mem_220_sv2v_reg  <= w_data_i[106];
      \nz.mem_219_sv2v_reg  <= w_data_i[105];
      \nz.mem_218_sv2v_reg  <= w_data_i[104];
      \nz.mem_217_sv2v_reg  <= w_data_i[103];
      \nz.mem_216_sv2v_reg  <= w_data_i[102];
      \nz.mem_215_sv2v_reg  <= w_data_i[101];
      \nz.mem_214_sv2v_reg  <= w_data_i[100];
      \nz.mem_213_sv2v_reg  <= w_data_i[99];
      \nz.mem_212_sv2v_reg  <= w_data_i[98];
      \nz.mem_211_sv2v_reg  <= w_data_i[97];
      \nz.mem_210_sv2v_reg  <= w_data_i[96];
      \nz.mem_209_sv2v_reg  <= w_data_i[95];
      \nz.mem_208_sv2v_reg  <= w_data_i[94];
      \nz.mem_207_sv2v_reg  <= w_data_i[93];
      \nz.mem_206_sv2v_reg  <= w_data_i[92];
      \nz.mem_205_sv2v_reg  <= w_data_i[91];
      \nz.mem_204_sv2v_reg  <= w_data_i[90];
      \nz.mem_203_sv2v_reg  <= w_data_i[89];
      \nz.mem_202_sv2v_reg  <= w_data_i[88];
      \nz.mem_201_sv2v_reg  <= w_data_i[87];
      \nz.mem_200_sv2v_reg  <= w_data_i[86];
      \nz.mem_199_sv2v_reg  <= w_data_i[85];
      \nz.mem_198_sv2v_reg  <= w_data_i[84];
      \nz.mem_197_sv2v_reg  <= w_data_i[83];
      \nz.mem_196_sv2v_reg  <= w_data_i[82];
      \nz.mem_195_sv2v_reg  <= w_data_i[81];
      \nz.mem_194_sv2v_reg  <= w_data_i[80];
      \nz.mem_193_sv2v_reg  <= w_data_i[79];
      \nz.mem_192_sv2v_reg  <= w_data_i[78];
      \nz.mem_191_sv2v_reg  <= w_data_i[77];
      \nz.mem_190_sv2v_reg  <= w_data_i[76];
      \nz.mem_189_sv2v_reg  <= w_data_i[75];
      \nz.mem_188_sv2v_reg  <= w_data_i[74];
      \nz.mem_187_sv2v_reg  <= w_data_i[73];
      \nz.mem_186_sv2v_reg  <= w_data_i[72];
      \nz.mem_185_sv2v_reg  <= w_data_i[71];
      \nz.mem_184_sv2v_reg  <= w_data_i[70];
      \nz.mem_183_sv2v_reg  <= w_data_i[69];
      \nz.mem_182_sv2v_reg  <= w_data_i[68];
      \nz.mem_181_sv2v_reg  <= w_data_i[67];
      \nz.mem_180_sv2v_reg  <= w_data_i[66];
      \nz.mem_179_sv2v_reg  <= w_data_i[65];
      \nz.mem_178_sv2v_reg  <= w_data_i[64];
      \nz.mem_177_sv2v_reg  <= w_data_i[63];
      \nz.mem_176_sv2v_reg  <= w_data_i[62];
      \nz.mem_175_sv2v_reg  <= w_data_i[61];
      \nz.mem_174_sv2v_reg  <= w_data_i[60];
      \nz.mem_173_sv2v_reg  <= w_data_i[59];
      \nz.mem_172_sv2v_reg  <= w_data_i[58];
      \nz.mem_171_sv2v_reg  <= w_data_i[57];
      \nz.mem_170_sv2v_reg  <= w_data_i[56];
      \nz.mem_169_sv2v_reg  <= w_data_i[55];
      \nz.mem_168_sv2v_reg  <= w_data_i[54];
      \nz.mem_167_sv2v_reg  <= w_data_i[53];
      \nz.mem_166_sv2v_reg  <= w_data_i[52];
      \nz.mem_165_sv2v_reg  <= w_data_i[51];
      \nz.mem_164_sv2v_reg  <= w_data_i[50];
      \nz.mem_163_sv2v_reg  <= w_data_i[49];
      \nz.mem_162_sv2v_reg  <= w_data_i[48];
      \nz.mem_161_sv2v_reg  <= w_data_i[47];
      \nz.mem_160_sv2v_reg  <= w_data_i[46];
      \nz.mem_159_sv2v_reg  <= w_data_i[45];
      \nz.mem_158_sv2v_reg  <= w_data_i[44];
      \nz.mem_157_sv2v_reg  <= w_data_i[43];
      \nz.mem_156_sv2v_reg  <= w_data_i[42];
      \nz.mem_155_sv2v_reg  <= w_data_i[41];
      \nz.mem_154_sv2v_reg  <= w_data_i[40];
      \nz.mem_153_sv2v_reg  <= w_data_i[39];
      \nz.mem_152_sv2v_reg  <= w_data_i[38];
      \nz.mem_151_sv2v_reg  <= w_data_i[37];
      \nz.mem_150_sv2v_reg  <= w_data_i[36];
      \nz.mem_149_sv2v_reg  <= w_data_i[35];
      \nz.mem_148_sv2v_reg  <= w_data_i[34];
      \nz.mem_147_sv2v_reg  <= w_data_i[33];
      \nz.mem_146_sv2v_reg  <= w_data_i[32];
      \nz.mem_145_sv2v_reg  <= w_data_i[31];
      \nz.mem_144_sv2v_reg  <= w_data_i[30];
      \nz.mem_143_sv2v_reg  <= w_data_i[29];
      \nz.mem_142_sv2v_reg  <= w_data_i[28];
      \nz.mem_141_sv2v_reg  <= w_data_i[27];
      \nz.mem_140_sv2v_reg  <= w_data_i[26];
      \nz.mem_139_sv2v_reg  <= w_data_i[25];
      \nz.mem_138_sv2v_reg  <= w_data_i[24];
      \nz.mem_137_sv2v_reg  <= w_data_i[23];
      \nz.mem_136_sv2v_reg  <= w_data_i[22];
      \nz.mem_135_sv2v_reg  <= w_data_i[21];
      \nz.mem_134_sv2v_reg  <= w_data_i[20];
      \nz.mem_133_sv2v_reg  <= w_data_i[19];
      \nz.mem_132_sv2v_reg  <= w_data_i[18];
      \nz.mem_131_sv2v_reg  <= w_data_i[17];
      \nz.mem_130_sv2v_reg  <= w_data_i[16];
      \nz.mem_129_sv2v_reg  <= w_data_i[15];
      \nz.mem_114_sv2v_reg  <= w_data_i[0];
    end 
    if(N20) begin
      \nz.mem_128_sv2v_reg  <= w_data_i[14];
      \nz.mem_127_sv2v_reg  <= w_data_i[13];
      \nz.mem_126_sv2v_reg  <= w_data_i[12];
      \nz.mem_125_sv2v_reg  <= w_data_i[11];
      \nz.mem_124_sv2v_reg  <= w_data_i[10];
      \nz.mem_123_sv2v_reg  <= w_data_i[9];
      \nz.mem_122_sv2v_reg  <= w_data_i[8];
      \nz.mem_121_sv2v_reg  <= w_data_i[7];
      \nz.mem_120_sv2v_reg  <= w_data_i[6];
      \nz.mem_119_sv2v_reg  <= w_data_i[5];
      \nz.mem_118_sv2v_reg  <= w_data_i[4];
      \nz.mem_117_sv2v_reg  <= w_data_i[3];
      \nz.mem_116_sv2v_reg  <= w_data_i[2];
      \nz.mem_115_sv2v_reg  <= w_data_i[1];
    end 
    if(N17) begin
      \nz.mem_113_sv2v_reg  <= w_data_i[113];
      \nz.mem_112_sv2v_reg  <= w_data_i[112];
      \nz.mem_111_sv2v_reg  <= w_data_i[111];
      \nz.mem_110_sv2v_reg  <= w_data_i[110];
      \nz.mem_109_sv2v_reg  <= w_data_i[109];
      \nz.mem_108_sv2v_reg  <= w_data_i[108];
      \nz.mem_107_sv2v_reg  <= w_data_i[107];
      \nz.mem_106_sv2v_reg  <= w_data_i[106];
      \nz.mem_105_sv2v_reg  <= w_data_i[105];
      \nz.mem_104_sv2v_reg  <= w_data_i[104];
      \nz.mem_103_sv2v_reg  <= w_data_i[103];
      \nz.mem_102_sv2v_reg  <= w_data_i[102];
      \nz.mem_101_sv2v_reg  <= w_data_i[101];
      \nz.mem_100_sv2v_reg  <= w_data_i[100];
      \nz.mem_99_sv2v_reg  <= w_data_i[99];
      \nz.mem_98_sv2v_reg  <= w_data_i[98];
      \nz.mem_97_sv2v_reg  <= w_data_i[97];
      \nz.mem_96_sv2v_reg  <= w_data_i[96];
      \nz.mem_95_sv2v_reg  <= w_data_i[95];
      \nz.mem_94_sv2v_reg  <= w_data_i[94];
      \nz.mem_93_sv2v_reg  <= w_data_i[93];
      \nz.mem_92_sv2v_reg  <= w_data_i[92];
      \nz.mem_91_sv2v_reg  <= w_data_i[91];
      \nz.mem_90_sv2v_reg  <= w_data_i[90];
      \nz.mem_89_sv2v_reg  <= w_data_i[89];
      \nz.mem_88_sv2v_reg  <= w_data_i[88];
      \nz.mem_87_sv2v_reg  <= w_data_i[87];
      \nz.mem_86_sv2v_reg  <= w_data_i[86];
      \nz.mem_85_sv2v_reg  <= w_data_i[85];
      \nz.mem_84_sv2v_reg  <= w_data_i[84];
      \nz.mem_83_sv2v_reg  <= w_data_i[83];
      \nz.mem_82_sv2v_reg  <= w_data_i[82];
      \nz.mem_81_sv2v_reg  <= w_data_i[81];
      \nz.mem_80_sv2v_reg  <= w_data_i[80];
      \nz.mem_79_sv2v_reg  <= w_data_i[79];
      \nz.mem_78_sv2v_reg  <= w_data_i[78];
      \nz.mem_77_sv2v_reg  <= w_data_i[77];
      \nz.mem_76_sv2v_reg  <= w_data_i[76];
      \nz.mem_75_sv2v_reg  <= w_data_i[75];
      \nz.mem_74_sv2v_reg  <= w_data_i[74];
      \nz.mem_73_sv2v_reg  <= w_data_i[73];
      \nz.mem_72_sv2v_reg  <= w_data_i[72];
      \nz.mem_71_sv2v_reg  <= w_data_i[71];
      \nz.mem_70_sv2v_reg  <= w_data_i[70];
      \nz.mem_69_sv2v_reg  <= w_data_i[69];
      \nz.mem_68_sv2v_reg  <= w_data_i[68];
      \nz.mem_67_sv2v_reg  <= w_data_i[67];
      \nz.mem_66_sv2v_reg  <= w_data_i[66];
      \nz.mem_65_sv2v_reg  <= w_data_i[65];
      \nz.mem_64_sv2v_reg  <= w_data_i[64];
      \nz.mem_63_sv2v_reg  <= w_data_i[63];
      \nz.mem_62_sv2v_reg  <= w_data_i[62];
      \nz.mem_61_sv2v_reg  <= w_data_i[61];
      \nz.mem_60_sv2v_reg  <= w_data_i[60];
      \nz.mem_59_sv2v_reg  <= w_data_i[59];
      \nz.mem_58_sv2v_reg  <= w_data_i[58];
      \nz.mem_57_sv2v_reg  <= w_data_i[57];
      \nz.mem_56_sv2v_reg  <= w_data_i[56];
      \nz.mem_55_sv2v_reg  <= w_data_i[55];
      \nz.mem_54_sv2v_reg  <= w_data_i[54];
      \nz.mem_53_sv2v_reg  <= w_data_i[53];
      \nz.mem_52_sv2v_reg  <= w_data_i[52];
      \nz.mem_51_sv2v_reg  <= w_data_i[51];
      \nz.mem_50_sv2v_reg  <= w_data_i[50];
      \nz.mem_49_sv2v_reg  <= w_data_i[49];
      \nz.mem_48_sv2v_reg  <= w_data_i[48];
      \nz.mem_47_sv2v_reg  <= w_data_i[47];
      \nz.mem_46_sv2v_reg  <= w_data_i[46];
      \nz.mem_45_sv2v_reg  <= w_data_i[45];
      \nz.mem_44_sv2v_reg  <= w_data_i[44];
      \nz.mem_43_sv2v_reg  <= w_data_i[43];
      \nz.mem_42_sv2v_reg  <= w_data_i[42];
      \nz.mem_41_sv2v_reg  <= w_data_i[41];
      \nz.mem_40_sv2v_reg  <= w_data_i[40];
      \nz.mem_39_sv2v_reg  <= w_data_i[39];
      \nz.mem_38_sv2v_reg  <= w_data_i[38];
      \nz.mem_37_sv2v_reg  <= w_data_i[37];
      \nz.mem_36_sv2v_reg  <= w_data_i[36];
      \nz.mem_35_sv2v_reg  <= w_data_i[35];
      \nz.mem_34_sv2v_reg  <= w_data_i[34];
      \nz.mem_33_sv2v_reg  <= w_data_i[33];
      \nz.mem_32_sv2v_reg  <= w_data_i[32];
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
    if(N18) begin
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
    end 
  end


endmodule



module bsg_mem_1r1w_114_00000004
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [1:0] w_addr_i;
  input [113:0] w_data_i;
  input [1:0] r_addr_i;
  output [113:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [113:0] r_data_o;

  bsg_mem_1r1w_synth_114_00000004_0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bp_be_cmd_queue_00
(
  clk_i,
  reset_i,
  fe_cmd_i,
  fe_cmd_v_i,
  fe_cmd_o,
  fe_cmd_v_o,
  fe_cmd_yumi_i,
  empty_n_o,
  empty_r_o,
  full_n_o,
  full_r_o
);

  input [113:0] fe_cmd_i;
  output [113:0] fe_cmd_o;
  input clk_i;
  input reset_i;
  input fe_cmd_v_i;
  input fe_cmd_yumi_i;
  output fe_cmd_v_o;
  output empty_n_o;
  output empty_r_o;
  output full_n_o;
  output full_r_o;
  wire [113:0] fe_cmd_o;
  wire fe_cmd_v_o,empty_n_o,empty_r_o,full_n_o,full_r_o,N0,N1,almost_full,N2,N3,
  almost_empty,N4,N5,N6,N7,N8,N9;
  wire [1:0] wptr_r,rptr_r,rptr_n;

  bsg_fifo_tracker_00000004
  ft
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .enq_i(fe_cmd_v_i),
    .deq_i(fe_cmd_yumi_i),
    .wptr_r_o(wptr_r),
    .rptr_r_o(rptr_r),
    .rptr_n_o(rptr_n),
    .full_o(full_r_o),
    .empty_o(empty_r_o)
  );


  bsg_mem_1r1w_114_00000004
  fifo_mem
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(fe_cmd_v_i),
    .w_addr_i(wptr_r),
    .w_data_i(fe_cmd_i),
    .r_v_i(fe_cmd_v_o),
    .r_addr_i(rptr_r),
    .r_data_o(fe_cmd_o)
  );

  assign almost_full = rptr_r == { N1, N0 };
  assign almost_empty = rptr_r == { N3, N2 };
  assign { N1, N0 } = wptr_r + 1'b1;
  assign { N3, N2 } = wptr_r - 1'b1;
  assign fe_cmd_v_o = ~empty_r_o;
  assign empty_n_o = N5 & N6;
  assign N5 = empty_r_o | N4;
  assign N4 = almost_empty & fe_cmd_yumi_i;
  assign N6 = ~fe_cmd_v_i;
  assign full_n_o = N8 & N9;
  assign N8 = full_r_o | N7;
  assign N7 = almost_full & fe_cmd_v_i;
  assign N9 = ~fe_cmd_yumi_i;

endmodule



module bp_be_director_00
(
  clk_i,
  reset_i,
  cfg_bus_i,
  issue_pkt_i,
  expected_npc_o,
  poison_isd_o,
  clear_iss_o,
  suppress_iss_o,
  resume_o,
  irq_waiting_i,
  mem_busy_i,
  cmd_full_n_o,
  cmd_full_r_o,
  fe_cmd_o,
  fe_cmd_v_o,
  fe_cmd_yumi_i,
  br_pkt_i,
  commit_pkt_i
);

  input [60:0] cfg_bus_i;
  input [263:0] issue_pkt_i;
  output [38:0] expected_npc_o;
  output [113:0] fe_cmd_o;
  input [42:0] br_pkt_i;
  input [213:0] commit_pkt_i;
  input clk_i;
  input reset_i;
  input irq_waiting_i;
  input mem_busy_i;
  input fe_cmd_yumi_i;
  output poison_isd_o;
  output clear_iss_o;
  output suppress_iss_o;
  output resume_o;
  output cmd_full_n_o;
  output cmd_full_r_o;
  output fe_cmd_v_o;
  wire [38:0] expected_npc_o,npc_n;
  wire [113:0] fe_cmd_o;
  wire poison_isd_o,clear_iss_o,suppress_iss_o,resume_o,cmd_full_n_o,cmd_full_r_o,
  fe_cmd_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,npc_w_v,N12,N13,N14,N15,N16,N17,
  npc_match_v,btaken_pending,attaboy_pending,fe_cmd_v_li,last_instr_was_branch,
  last_instr_was_btaken,fe_cmd_li_npc__38_,fe_cmd_li_npc__37_,fe_cmd_li_npc__36_,
  fe_cmd_li_npc__35_,fe_cmd_li_npc__34_,fe_cmd_li_npc__33_,fe_cmd_li_npc__32_,
  fe_cmd_li_npc__31_,fe_cmd_li_npc__30_,fe_cmd_li_npc__29_,fe_cmd_li_npc__28_,
  fe_cmd_li_npc__27_,fe_cmd_li_npc__26_,fe_cmd_li_npc__25_,fe_cmd_li_npc__24_,fe_cmd_li_npc__23_,
  fe_cmd_li_npc__22_,fe_cmd_li_npc__21_,fe_cmd_li_npc__20_,fe_cmd_li_npc__19_,
  fe_cmd_li_npc__18_,fe_cmd_li_npc__17_,fe_cmd_li_npc__16_,fe_cmd_li_npc__15_,
  fe_cmd_li_npc__14_,fe_cmd_li_npc__13_,fe_cmd_li_npc__12_,fe_cmd_li_npc__11_,
  fe_cmd_li_npc__10_,fe_cmd_li_npc__9_,fe_cmd_li_npc__8_,fe_cmd_li_npc__7_,fe_cmd_li_npc__6_,
  fe_cmd_li_npc__5_,fe_cmd_li_npc__4_,fe_cmd_li_npc__3_,fe_cmd_li_npc__2_,
  fe_cmd_li_npc__1_,fe_cmd_li_npc__0_,fe_cmd_li_opcode__2_,fe_cmd_li_opcode__1_,
  fe_cmd_li_opcode__0_,fe_cmd_li_operands__71_,fe_cmd_li_operands__70_,
  fe_cmd_li_operands__69_,fe_cmd_li_operands__68_,fe_cmd_li_operands__67_,fe_cmd_li_operands__66_,
  fe_cmd_li_operands__65_,fe_cmd_li_operands__64_,fe_cmd_li_operands__63_,
  fe_cmd_li_operands__62_,fe_cmd_li_operands__61_,fe_cmd_li_operands__60_,
  fe_cmd_li_operands__59_,fe_cmd_li_operands__58_,fe_cmd_li_operands__57_,fe_cmd_li_operands__56_,
  fe_cmd_li_operands__55_,fe_cmd_li_operands__54_,fe_cmd_li_operands__53_,
  fe_cmd_li_operands__52_,fe_cmd_li_operands__51_,fe_cmd_li_operands__50_,
  fe_cmd_li_operands__49_,fe_cmd_li_operands__48_,fe_cmd_li_operands__47_,fe_cmd_li_operands__46_,
  fe_cmd_li_operands__45_,fe_cmd_li_operands__44_,fe_cmd_li_operands__43_,
  fe_cmd_li_operands__42_,fe_cmd_li_operands__41_,fe_cmd_li_operands__40_,
  fe_cmd_li_operands__39_,fe_cmd_li_operands__38_,fe_cmd_li_operands__37_,fe_cmd_li_operands__36_,
  fe_cmd_li_operands__35_,fe_cmd_li_operands__34_,fe_cmd_li_operands__33_,
  fe_cmd_li_operands__32_,fe_cmd_li_operands__31_,fe_cmd_li_operands__30_,
  fe_cmd_li_operands__29_,fe_cmd_li_operands__28_,fe_cmd_li_operands__27_,fe_cmd_li_operands__26_,
  fe_cmd_li_operands__25_,fe_cmd_li_operands__24_,fe_cmd_li_operands__23_,
  fe_cmd_li_operands__22_,fe_cmd_li_operands__21_,fe_cmd_li_operands__20_,
  fe_cmd_li_operands__19_,fe_cmd_li_operands__18_,fe_cmd_li_operands__17_,fe_cmd_li_operands__16_,
  fe_cmd_li_operands__15_,fe_cmd_li_operands__14_,fe_cmd_li_operands__13_,
  fe_cmd_li_operands__12_,fe_cmd_li_operands__11_,fe_cmd_li_operands__10_,fe_cmd_li_operands__9_,
  fe_cmd_li_operands__8_,fe_cmd_li_operands__7_,fe_cmd_li_operands__6_,
  fe_cmd_li_operands__5_,fe_cmd_li_operands__4_,fe_cmd_li_operands__3_,
  fe_cmd_li_operands__2_,fe_cmd_li_operands__1_,fe_cmd_nonattaboy_v,freeze_li,N18,N19,N20,N21,N22,N23,
  N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,
  N44,N45,cmd_empty_r_lo,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,cmd_empty_n_lo,N109,N110,N111,N112,
  N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,
  N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,
  N145,N146,N147;
  wire [3:0] state_r,state_n;
  reg state_r_3_sv2v_reg,state_r_2_sv2v_reg,state_r_1_sv2v_reg,state_r_0_sv2v_reg;
  assign state_r[3] = state_r_3_sv2v_reg;
  assign state_r[2] = state_r_2_sv2v_reg;
  assign state_r[1] = state_r_1_sv2v_reg;
  assign state_r[0] = state_r_0_sv2v_reg;

  bsg_dff_reset_en_bypass_00000027
  npc_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(npc_w_v),
    .data_i(npc_n),
    .data_o(expected_npc_o)
  );

  assign N16 = expected_npc_o != issue_pkt_i[244:206];
  assign N17 = expected_npc_o == issue_pkt_i[244:206];

  bsg_dff_reset_set_clear_width_p2_clear_over_set_p1
  attaboy_pending_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .set_i({ br_pkt_i[40:40], br_pkt_i[41:41] }),
    .clear_i({ fe_cmd_v_li, fe_cmd_v_li }),
    .data_o({ btaken_pending, attaboy_pending })
  );

  assign N18 = state_r[3] | state_r[2];
  assign N19 = N111 | state_r[0];
  assign N20 = N18 | N19;
  assign N23 = N22 & N120;
  assign N24 = N111 & N112;
  assign N25 = N23 & N24;
  assign N26 = state_r[3] | state_r[2];
  assign N27 = state_r[1] | N112;
  assign N28 = N26 | N27;
  assign N29 = state_r[3] | N120;
  assign N30 = state_r[1] | state_r[0];
  assign N31 = N29 | N30;
  assign N33 = state_r[2] & state_r[0];
  assign N34 = state_r[1] & state_r[0];
  assign N35 = state_r[2] & state_r[1];

  bp_be_cmd_queue_00
  fe_cmd_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .fe_cmd_i({ fe_cmd_li_npc__38_, fe_cmd_li_npc__37_, fe_cmd_li_npc__36_, fe_cmd_li_npc__35_, fe_cmd_li_npc__34_, fe_cmd_li_npc__33_, fe_cmd_li_npc__32_, fe_cmd_li_npc__31_, fe_cmd_li_npc__30_, fe_cmd_li_npc__29_, fe_cmd_li_npc__28_, fe_cmd_li_npc__27_, fe_cmd_li_npc__26_, fe_cmd_li_npc__25_, fe_cmd_li_npc__24_, fe_cmd_li_npc__23_, fe_cmd_li_npc__22_, fe_cmd_li_npc__21_, fe_cmd_li_npc__20_, fe_cmd_li_npc__19_, fe_cmd_li_npc__18_, fe_cmd_li_npc__17_, fe_cmd_li_npc__16_, fe_cmd_li_npc__15_, fe_cmd_li_npc__14_, fe_cmd_li_npc__13_, fe_cmd_li_npc__12_, fe_cmd_li_npc__11_, fe_cmd_li_npc__10_, fe_cmd_li_npc__9_, fe_cmd_li_npc__8_, fe_cmd_li_npc__7_, fe_cmd_li_npc__6_, fe_cmd_li_npc__5_, fe_cmd_li_npc__4_, fe_cmd_li_npc__3_, fe_cmd_li_npc__2_, fe_cmd_li_npc__1_, fe_cmd_li_npc__0_, fe_cmd_li_opcode__2_, fe_cmd_li_opcode__1_, fe_cmd_li_opcode__0_, fe_cmd_li_operands__71_, fe_cmd_li_operands__70_, fe_cmd_li_operands__69_, fe_cmd_li_operands__68_, fe_cmd_li_operands__67_, fe_cmd_li_operands__66_, fe_cmd_li_operands__65_, fe_cmd_li_operands__64_, fe_cmd_li_operands__63_, fe_cmd_li_operands__62_, fe_cmd_li_operands__61_, fe_cmd_li_operands__60_, fe_cmd_li_operands__59_, fe_cmd_li_operands__58_, fe_cmd_li_operands__57_, fe_cmd_li_operands__56_, fe_cmd_li_operands__55_, fe_cmd_li_operands__54_, fe_cmd_li_operands__53_, fe_cmd_li_operands__52_, fe_cmd_li_operands__51_, fe_cmd_li_operands__50_, fe_cmd_li_operands__49_, fe_cmd_li_operands__48_, fe_cmd_li_operands__47_, fe_cmd_li_operands__46_, fe_cmd_li_operands__45_, fe_cmd_li_operands__44_, fe_cmd_li_operands__43_, fe_cmd_li_operands__42_, fe_cmd_li_operands__41_, fe_cmd_li_operands__40_, fe_cmd_li_operands__39_, fe_cmd_li_operands__38_, fe_cmd_li_operands__37_, fe_cmd_li_operands__36_, fe_cmd_li_operands__35_, fe_cmd_li_operands__34_, fe_cmd_li_operands__33_, fe_cmd_li_operands__32_, fe_cmd_li_operands__31_, fe_cmd_li_operands__30_, fe_cmd_li_operands__29_, fe_cmd_li_operands__28_, fe_cmd_li_operands__27_, fe_cmd_li_operands__26_, fe_cmd_li_operands__25_, fe_cmd_li_operands__24_, fe_cmd_li_operands__23_, fe_cmd_li_operands__22_, fe_cmd_li_operands__21_, fe_cmd_li_operands__20_, fe_cmd_li_operands__19_, fe_cmd_li_operands__18_, fe_cmd_li_operands__17_, fe_cmd_li_operands__16_, fe_cmd_li_operands__15_, fe_cmd_li_operands__14_, fe_cmd_li_operands__13_, fe_cmd_li_operands__12_, fe_cmd_li_operands__11_, fe_cmd_li_operands__10_, fe_cmd_li_operands__9_, fe_cmd_li_operands__8_, fe_cmd_li_operands__7_, fe_cmd_li_operands__6_, fe_cmd_li_operands__5_, fe_cmd_li_operands__4_, fe_cmd_li_operands__3_, fe_cmd_li_operands__2_, fe_cmd_li_operands__1_, 1'b0 }),
    .fe_cmd_v_i(fe_cmd_v_li),
    .fe_cmd_o(fe_cmd_o),
    .fe_cmd_v_o(fe_cmd_v_o),
    .fe_cmd_yumi_i(fe_cmd_yumi_i),
    .empty_n_o(cmd_empty_n_lo),
    .empty_r_o(cmd_empty_r_lo),
    .full_n_o(cmd_full_n_o),
    .full_r_o(cmd_full_r_o)
  );

  assign N111 = ~state_r[1];
  assign N112 = ~state_r[0];
  assign N113 = state_r[2] | state_r[3];
  assign N114 = N111 | N113;
  assign N115 = N112 | N114;
  assign N116 = ~N115;
  assign N117 = state_r[2] | state_r[3];
  assign N118 = N111 | N117;
  assign N119 = state_r[0] | N118;
  assign N120 = ~state_r[2];
  assign N121 = N120 | state_r[3];
  assign N122 = state_r[1] | N121;
  assign N123 = state_r[0] | N122;
  assign N124 = ~N123;
  assign N125 = ~fe_cmd_li_opcode__1_;
  assign N126 = N125 | fe_cmd_li_opcode__2_;
  assign N127 = fe_cmd_li_opcode__0_ | N126;
  assign N128 = state_r[2] | state_r[3];
  assign N129 = state_r[1] | N128;
  assign N130 = N112 | N129;
  assign N131 = ~N130;
  assign N132 = state_r[2] | state_r[3];
  assign N133 = state_r[1] | N132;
  assign N134 = state_r[0] | N133;
  assign N135 = ~N134;
  assign npc_n = (N0)? commit_pkt_i[166:128] : 
                 (N15)? issue_pkt_i[244:206] : 
                 (N13)? br_pkt_i[38:0] : 1'b0;
  assign N0 = commit_pkt_i[213];
  assign { N44, N43, N42, N41 } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N52)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                  (N55)? { 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                  (N58)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                  (N40)? state_r : 1'b0;
  assign N1 = freeze_li;
  assign { N50, N49, N48, N47 } = (N2)? { 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                  (N3)? state_r : 1'b0;
  assign N2 = cmd_empty_r_lo;
  assign N3 = N46;
  assign state_n = (N4)? { N44, N43, N42, N41 } : 
                   (N5)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                   (N6)? { N50, N49, N48, N47 } : 1'b0;
  assign N4 = N21;
  assign N5 = N32;
  assign N6 = N36;
  assign { N74, N73 } = (N7)? { 1'b0, 1'b0 } : 
                        (N108)? { 1'b1, 1'b0 } : 
                        (N72)? { 1'b0, 1'b1 } : 1'b0;
  assign N7 = N135;
  assign { N78, N77 } = (N8)? { N76, last_instr_was_btaken } : 
                        (N9)? { 1'b0, 1'b0 } : 1'b0;
  assign N8 = last_instr_was_branch;
  assign N9 = N75;
  assign { fe_cmd_li_operands__14_, fe_cmd_li_operands__13_, fe_cmd_li_operands__12_, fe_cmd_li_operands__11_, fe_cmd_li_operands__10_, fe_cmd_li_operands__9_, fe_cmd_li_operands__8_, fe_cmd_li_operands__7_, fe_cmd_li_operands__6_, fe_cmd_li_operands__5_, fe_cmd_li_operands__4_, fe_cmd_li_operands__3_, fe_cmd_li_operands__2_, fe_cmd_li_operands__1_ } = (N84)? { commit_pkt_i[67:57], commit_pkt_i[210:208] } : 
                                                                                                                                                                                                                                                                                                                                                                   (N80)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { fe_cmd_li_operands__17_, fe_cmd_li_operands__16_, fe_cmd_li_operands__15_ } = (N10)? { commit_pkt_i[18:18], commit_pkt_i[20:19] } : 
                                                                                         (N84)? commit_pkt_i[70:68] : 
                                                                                         (N87)? { 1'b0, 1'b0, 1'b0 } : 
                                                                                         (N90)? { commit_pkt_i[18:18], 1'b0, 1'b0 } : 
                                                                                         (N93)? { 1'b0, 1'b0, 1'b0 } : 
                                                                                         (N95)? { 1'b0, 1'b0, 1'b0 } : 
                                                                                         (N98)? { commit_pkt_i[18:18], commit_pkt_i[20:19] } : 
                                                                                         (N101)? { commit_pkt_i[18:18], commit_pkt_i[20:19] } : 
                                                                                         (N81)? { 1'b0, 1'b0, 1'b0 } : 
                                                                                         (N11)? { 1'b0, 1'b0, 1'b0 } : 
                                                                                         (N11)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = commit_pkt_i[15];
  assign N11 = 1'b0;
  assign { fe_cmd_li_opcode__0_, fe_cmd_li_operands__21_, fe_cmd_li_operands__20_, fe_cmd_li_operands__19_, fe_cmd_li_operands__18_ } = (N10)? { N73, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                        (N84)? { 1'b1, commit_pkt_i[74:71] } : 
                                                                                                                                        (N87)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                        (N90)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                        (N93)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                        (N95)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                        (N98)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                        (N101)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                        (N104)? { 1'b1, issue_pkt_i[1:0], N78, N77 } : 
                                                                                                                                        (N82)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                        (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { fe_cmd_li_npc__38_, fe_cmd_li_npc__37_, fe_cmd_li_npc__36_, fe_cmd_li_npc__35_, fe_cmd_li_npc__34_, fe_cmd_li_npc__33_, fe_cmd_li_npc__32_, fe_cmd_li_npc__31_, fe_cmd_li_npc__30_, fe_cmd_li_npc__29_, fe_cmd_li_npc__28_, fe_cmd_li_npc__27_, fe_cmd_li_npc__26_, fe_cmd_li_npc__25_, fe_cmd_li_npc__24_, fe_cmd_li_npc__23_, fe_cmd_li_npc__22_, fe_cmd_li_npc__21_, fe_cmd_li_npc__20_, fe_cmd_li_npc__19_, fe_cmd_li_npc__18_, fe_cmd_li_npc__17_, fe_cmd_li_npc__16_, fe_cmd_li_npc__15_, fe_cmd_li_npc__14_, fe_cmd_li_npc__13_, fe_cmd_li_npc__12_, fe_cmd_li_npc__11_, fe_cmd_li_npc__10_, fe_cmd_li_npc__9_, fe_cmd_li_npc__8_, fe_cmd_li_npc__7_, fe_cmd_li_npc__6_, fe_cmd_li_npc__5_, fe_cmd_li_npc__4_, fe_cmd_li_npc__3_, fe_cmd_li_npc__2_, fe_cmd_li_npc__1_, fe_cmd_li_npc__0_, fe_cmd_li_opcode__1_, fe_cmd_li_operands__71_, fe_cmd_li_operands__70_, fe_cmd_li_operands__69_, fe_cmd_li_operands__68_, fe_cmd_li_operands__67_, fe_cmd_li_operands__66_, fe_cmd_li_operands__65_, fe_cmd_li_operands__64_, fe_cmd_li_operands__63_, fe_cmd_li_operands__62_, fe_cmd_li_operands__61_, fe_cmd_li_operands__60_, fe_cmd_li_operands__59_, fe_cmd_li_operands__58_, fe_cmd_li_operands__57_, fe_cmd_li_operands__56_, fe_cmd_li_operands__55_, fe_cmd_li_operands__54_, fe_cmd_li_operands__53_, fe_cmd_li_operands__52_, fe_cmd_li_operands__51_, fe_cmd_li_operands__50_, fe_cmd_li_operands__49_, fe_cmd_li_operands__48_, fe_cmd_li_operands__47_, fe_cmd_li_operands__46_, fe_cmd_li_operands__45_, fe_cmd_li_operands__44_, fe_cmd_li_operands__43_, fe_cmd_li_operands__42_, fe_cmd_li_operands__41_, fe_cmd_li_operands__40_, fe_cmd_li_operands__39_, fe_cmd_li_operands__38_, fe_cmd_li_operands__37_, fe_cmd_li_operands__36_, fe_cmd_li_operands__35_, fe_cmd_li_operands__34_, fe_cmd_li_operands__33_, fe_cmd_li_operands__32_, fe_cmd_li_operands__31_, fe_cmd_li_operands__30_, fe_cmd_li_operands__29_, fe_cmd_li_operands__28_, fe_cmd_li_operands__27_, fe_cmd_li_operands__26_, fe_cmd_li_operands__25_, fe_cmd_li_operands__24_, fe_cmd_li_operands__23_, fe_cmd_li_operands__22_ } = (N10)? { npc_n, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N84)? { commit_pkt_i[127:89], 1'b0, commit_pkt_i[56:21], commit_pkt_i[88:75] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N87)? { commit_pkt_i[166:128], 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N90)? { commit_pkt_i[166:128], 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N93)? { commit_pkt_i[166:128], 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N95)? { commit_pkt_i[127:89], 1'b1, commit_pkt_i[88:57], commit_pkt_i[210:208], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N98)? { commit_pkt_i[166:128], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N101)? { commit_pkt_i[166:128], 1'b0, 1'b0, commit_pkt_i[17:17], 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N104)? { expected_npc_o, 1'b0, 1'b0, 1'b1, 1'b0, issue_pkt_i[48:2] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N107)? { expected_npc_o, 1'b1, last_instr_was_btaken, issue_pkt_i[48:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N70)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign fe_cmd_li_opcode__2_ = (N10)? N74 : 
                                (N84)? 1'b1 : 
                                (N87)? 1'b1 : 
                                (N90)? 1'b0 : 
                                (N93)? 1'b1 : 
                                (N83)? 1'b0 : 
                                (N11)? 1'b0 : 
                                (N11)? 1'b0 : 
                                (N11)? 1'b0 : 
                                (N11)? 1'b0 : 
                                (N11)? 1'b0 : 1'b0;
  assign fe_cmd_v_li = (N10)? 1'b1 : 
                       (N84)? 1'b1 : 
                       (N87)? 1'b1 : 
                       (N90)? 1'b1 : 
                       (N93)? 1'b1 : 
                       (N95)? 1'b1 : 
                       (N98)? 1'b1 : 
                       (N101)? 1'b1 : 
                       (N104)? 1'b1 : 
                       (N107)? 1'b1 : 
                       (N70)? 1'b0 : 1'b0;
  assign npc_w_v = commit_pkt_i[213] | br_pkt_i[42];
  assign N12 = br_pkt_i[39] | commit_pkt_i[213];
  assign N13 = ~N12;
  assign N14 = ~commit_pkt_i[213];
  assign N15 = br_pkt_i[39] & N14;
  assign poison_isd_o = issue_pkt_i[263] & N16;
  assign npc_match_v = issue_pkt_i[263] & N17;
  assign last_instr_was_branch = attaboy_pending | br_pkt_i[41];
  assign last_instr_was_btaken = btaken_pending | br_pkt_i[40];
  assign fe_cmd_nonattaboy_v = fe_cmd_v_li & N127;
  assign freeze_li = cfg_bus_i[60] | reset_i;
  assign N21 = ~N20;
  assign N22 = ~state_r[3];
  assign N32 = N137 | N138;
  assign N137 = N25 | N136;
  assign N136 = ~N28;
  assign N138 = ~N31;
  assign N36 = state_r[3] | N140;
  assign N140 = N33 | N139;
  assign N139 = N34 | N35;
  assign N37 = commit_pkt_i[10] | freeze_li;
  assign N38 = commit_pkt_i[13] | N37;
  assign N39 = fe_cmd_nonattaboy_v | N38;
  assign N40 = ~N39;
  assign N45 = ~commit_pkt_i[15];
  assign N46 = ~cmd_empty_r_lo;
  assign N51 = ~freeze_li;
  assign N52 = commit_pkt_i[10] & N51;
  assign N53 = ~commit_pkt_i[10];
  assign N54 = N51 & N53;
  assign N55 = commit_pkt_i[13] & N54;
  assign N56 = ~commit_pkt_i[13];
  assign N57 = N54 & N56;
  assign N58 = fe_cmd_nonattaboy_v & N57;
  assign suppress_iss_o = N141 | commit_pkt_i[213];
  assign N141 = N119 | cmd_full_r_o;
  assign clear_iss_o = N116 & cmd_empty_r_lo;
  assign resume_o = N145 | N147;
  assign N145 = N143 | N144;
  assign N143 = N135 & N142;
  assign N142 = ~freeze_li;
  assign N144 = N124 & irq_waiting_i;
  assign N147 = N131 & N146;
  assign N146 = ~mem_busy_i;
  assign N59 = commit_pkt_i[17] | commit_pkt_i[16];
  assign N60 = npc_match_v & last_instr_was_branch;
  assign N61 = commit_pkt_i[3] | commit_pkt_i[15];
  assign N62 = commit_pkt_i[12] | N61;
  assign N63 = commit_pkt_i[11] | N62;
  assign N64 = commit_pkt_i[10] | N63;
  assign N65 = commit_pkt_i[8] | N64;
  assign N66 = commit_pkt_i[14] | N65;
  assign N67 = N59 | N66;
  assign N68 = poison_isd_o | N67;
  assign N69 = N60 | N68;
  assign N70 = ~N69;
  assign N71 = N131 | N135;
  assign N72 = ~N71;
  assign N75 = ~last_instr_was_branch;
  assign N76 = ~last_instr_was_btaken;
  assign N79 = ~N84;
  assign N80 = N79;
  assign N81 = ~N67;
  assign N82 = ~N68;
  assign N83 = ~N64;
  assign N84 = commit_pkt_i[3] & N45;
  assign N85 = ~commit_pkt_i[3];
  assign N86 = N45 & N85;
  assign N87 = commit_pkt_i[12] & N86;
  assign N88 = ~commit_pkt_i[12];
  assign N89 = N86 & N88;
  assign N90 = commit_pkt_i[11] & N89;
  assign N91 = ~commit_pkt_i[11];
  assign N92 = N89 & N91;
  assign N93 = commit_pkt_i[10] & N92;
  assign N94 = N92 & N53;
  assign N95 = commit_pkt_i[8] & N94;
  assign N96 = ~commit_pkt_i[8];
  assign N97 = N94 & N96;
  assign N98 = commit_pkt_i[14] & N97;
  assign N99 = ~commit_pkt_i[14];
  assign N100 = N97 & N99;
  assign N101 = N59 & N100;
  assign N102 = ~N59;
  assign N103 = N100 & N102;
  assign N104 = poison_isd_o & N103;
  assign N105 = ~poison_isd_o;
  assign N106 = N103 & N105;
  assign N107 = N60 & N106;
  assign N108 = N131 & N134;
  assign N109 = N45 & N32;
  assign N110 = ~N109;

  always @(posedge clk_i) begin
    if(reset_i) begin
      state_r_3_sv2v_reg <= 1'b0;
      state_r_2_sv2v_reg <= 1'b0;
      state_r_1_sv2v_reg <= 1'b0;
      state_r_0_sv2v_reg <= 1'b0;
    end else if(N110) begin
      state_r_3_sv2v_reg <= state_n[3];
      state_r_2_sv2v_reg <= state_n[2];
      state_r_1_sv2v_reg <= state_n[1];
      state_r_0_sv2v_reg <= state_n[0];
    end 
  end


endmodule



module bsg_decode_num_out_p32
(
  i,
  o
);

  input [4:0] i;
  output [31:0] o;
  wire [31:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_decode_with_v_num_out_p32
(
  i,
  v_i,
  o
);

  input [4:0] i;
  output [31:0] o;
  input v_i;
  wire [31:0] o,lo;

  bsg_decode_num_out_p32
  bd
  (
    .i(i),
    .o(lo)
  );

  assign o[31] = v_i & lo[31];
  assign o[30] = v_i & lo[30];
  assign o[29] = v_i & lo[29];
  assign o[28] = v_i & lo[28];
  assign o[27] = v_i & lo[27];
  assign o[26] = v_i & lo[26];
  assign o[25] = v_i & lo[25];
  assign o[24] = v_i & lo[24];
  assign o[23] = v_i & lo[23];
  assign o[22] = v_i & lo[22];
  assign o[21] = v_i & lo[21];
  assign o[20] = v_i & lo[20];
  assign o[19] = v_i & lo[19];
  assign o[18] = v_i & lo[18];
  assign o[17] = v_i & lo[17];
  assign o[16] = v_i & lo[16];
  assign o[15] = v_i & lo[15];
  assign o[14] = v_i & lo[14];
  assign o[13] = v_i & lo[13];
  assign o[12] = v_i & lo[12];
  assign o[11] = v_i & lo[11];
  assign o[10] = v_i & lo[10];
  assign o[9] = v_i & lo[9];
  assign o[8] = v_i & lo[8];
  assign o[7] = v_i & lo[7];
  assign o[6] = v_i & lo[6];
  assign o[5] = v_i & lo[5];
  assign o[4] = v_i & lo[4];
  assign o[3] = v_i & lo[3];
  assign o[2] = v_i & lo[2];
  assign o[1] = v_i & lo[1];
  assign o[0] = v_i & lo[0];

endmodule



module bsg_dff_reset_set_clear_width_p32_clear_over_set_p1
(
  clk_i,
  reset_i,
  set_i,
  clear_i,
  data_o
);

  input [31:0] set_i;
  input [31:0] clear_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  wire [31:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95;
  reg data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,
  data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,
  data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,
  data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N0 = N32 & N33;
  assign N32 = data_o[31] | set_i[31];
  assign N33 = ~clear_i[31];
  assign N1 = N34 & N35;
  assign N34 = data_o[30] | set_i[30];
  assign N35 = ~clear_i[30];
  assign N2 = N36 & N37;
  assign N36 = data_o[29] | set_i[29];
  assign N37 = ~clear_i[29];
  assign N3 = N38 & N39;
  assign N38 = data_o[28] | set_i[28];
  assign N39 = ~clear_i[28];
  assign N4 = N40 & N41;
  assign N40 = data_o[27] | set_i[27];
  assign N41 = ~clear_i[27];
  assign N5 = N42 & N43;
  assign N42 = data_o[26] | set_i[26];
  assign N43 = ~clear_i[26];
  assign N6 = N44 & N45;
  assign N44 = data_o[25] | set_i[25];
  assign N45 = ~clear_i[25];
  assign N7 = N46 & N47;
  assign N46 = data_o[24] | set_i[24];
  assign N47 = ~clear_i[24];
  assign N8 = N48 & N49;
  assign N48 = data_o[23] | set_i[23];
  assign N49 = ~clear_i[23];
  assign N9 = N50 & N51;
  assign N50 = data_o[22] | set_i[22];
  assign N51 = ~clear_i[22];
  assign N10 = N52 & N53;
  assign N52 = data_o[21] | set_i[21];
  assign N53 = ~clear_i[21];
  assign N11 = N54 & N55;
  assign N54 = data_o[20] | set_i[20];
  assign N55 = ~clear_i[20];
  assign N12 = N56 & N57;
  assign N56 = data_o[19] | set_i[19];
  assign N57 = ~clear_i[19];
  assign N13 = N58 & N59;
  assign N58 = data_o[18] | set_i[18];
  assign N59 = ~clear_i[18];
  assign N14 = N60 & N61;
  assign N60 = data_o[17] | set_i[17];
  assign N61 = ~clear_i[17];
  assign N15 = N62 & N63;
  assign N62 = data_o[16] | set_i[16];
  assign N63 = ~clear_i[16];
  assign N16 = N64 & N65;
  assign N64 = data_o[15] | set_i[15];
  assign N65 = ~clear_i[15];
  assign N17 = N66 & N67;
  assign N66 = data_o[14] | set_i[14];
  assign N67 = ~clear_i[14];
  assign N18 = N68 & N69;
  assign N68 = data_o[13] | set_i[13];
  assign N69 = ~clear_i[13];
  assign N19 = N70 & N71;
  assign N70 = data_o[12] | set_i[12];
  assign N71 = ~clear_i[12];
  assign N20 = N72 & N73;
  assign N72 = data_o[11] | set_i[11];
  assign N73 = ~clear_i[11];
  assign N21 = N74 & N75;
  assign N74 = data_o[10] | set_i[10];
  assign N75 = ~clear_i[10];
  assign N22 = N76 & N77;
  assign N76 = data_o[9] | set_i[9];
  assign N77 = ~clear_i[9];
  assign N23 = N78 & N79;
  assign N78 = data_o[8] | set_i[8];
  assign N79 = ~clear_i[8];
  assign N24 = N80 & N81;
  assign N80 = data_o[7] | set_i[7];
  assign N81 = ~clear_i[7];
  assign N25 = N82 & N83;
  assign N82 = data_o[6] | set_i[6];
  assign N83 = ~clear_i[6];
  assign N26 = N84 & N85;
  assign N84 = data_o[5] | set_i[5];
  assign N85 = ~clear_i[5];
  assign N27 = N86 & N87;
  assign N86 = data_o[4] | set_i[4];
  assign N87 = ~clear_i[4];
  assign N28 = N88 & N89;
  assign N88 = data_o[3] | set_i[3];
  assign N89 = ~clear_i[3];
  assign N29 = N90 & N91;
  assign N90 = data_o[2] | set_i[2];
  assign N91 = ~clear_i[2];
  assign N30 = N92 & N93;
  assign N92 = data_o[1] | set_i[1];
  assign N93 = ~clear_i[1];
  assign N31 = N94 & N95;
  assign N94 = data_o[0] | set_i[0];
  assign N95 = ~clear_i[0];

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_31_sv2v_reg <= N0;
      data_o_30_sv2v_reg <= N1;
      data_o_29_sv2v_reg <= N2;
      data_o_28_sv2v_reg <= N3;
      data_o_27_sv2v_reg <= N4;
      data_o_26_sv2v_reg <= N5;
      data_o_25_sv2v_reg <= N6;
      data_o_24_sv2v_reg <= N7;
      data_o_23_sv2v_reg <= N8;
      data_o_22_sv2v_reg <= N9;
      data_o_21_sv2v_reg <= N10;
      data_o_20_sv2v_reg <= N11;
      data_o_19_sv2v_reg <= N12;
      data_o_18_sv2v_reg <= N13;
      data_o_17_sv2v_reg <= N14;
      data_o_16_sv2v_reg <= N15;
      data_o_15_sv2v_reg <= N16;
      data_o_14_sv2v_reg <= N17;
      data_o_13_sv2v_reg <= N18;
      data_o_12_sv2v_reg <= N19;
      data_o_11_sv2v_reg <= N20;
      data_o_10_sv2v_reg <= N21;
      data_o_9_sv2v_reg <= N22;
      data_o_8_sv2v_reg <= N23;
      data_o_7_sv2v_reg <= N24;
      data_o_6_sv2v_reg <= N25;
      data_o_5_sv2v_reg <= N26;
      data_o_4_sv2v_reg <= N27;
      data_o_3_sv2v_reg <= N28;
      data_o_2_sv2v_reg <= N29;
      data_o_1_sv2v_reg <= N30;
      data_o_0_sv2v_reg <= N31;
    end 
  end


endmodule



module bp_be_scoreboard_00_2
(
  clk_i,
  reset_i,
  score_v_i,
  score_rd_i,
  clear_v_i,
  clear_rd_i,
  check_rs_i,
  check_rd_i,
  rs_match_o,
  rd_match_o
);

  input [4:0] score_rd_i;
  input [4:0] clear_rd_i;
  input [9:0] check_rs_i;
  input [4:0] check_rd_i;
  output [1:0] rs_match_o;
  input clk_i;
  input reset_i;
  input score_v_i;
  input clear_v_i;
  output rd_match_o;
  wire [1:0] rs_match_o;
  wire rd_match_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,
  N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,
  N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,
  N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194;
  wire [31:0] score_onehot_li,clear_onehot_li,scoreboard_r;

  bsg_decode_with_v_num_out_p32
  score_decode
  (
    .i(score_rd_i),
    .v_i(score_v_i),
    .o(score_onehot_li)
  );


  bsg_decode_with_v_num_out_p32
  clear_decode
  (
    .i(clear_rd_i),
    .v_i(clear_v_i),
    .o(clear_onehot_li)
  );


  bsg_dff_reset_set_clear_width_p32_clear_over_set_p1
  scoreboard_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .set_i(score_onehot_li),
    .clear_i(clear_onehot_li),
    .data_o(scoreboard_r)
  );

  assign rs_match_o[0] = (N33)? scoreboard_r[0] : 
                         (N35)? scoreboard_r[1] : 
                         (N37)? scoreboard_r[2] : 
                         (N39)? scoreboard_r[3] : 
                         (N41)? scoreboard_r[4] : 
                         (N43)? scoreboard_r[5] : 
                         (N45)? scoreboard_r[6] : 
                         (N47)? scoreboard_r[7] : 
                         (N49)? scoreboard_r[8] : 
                         (N51)? scoreboard_r[9] : 
                         (N53)? scoreboard_r[10] : 
                         (N55)? scoreboard_r[11] : 
                         (N57)? scoreboard_r[12] : 
                         (N59)? scoreboard_r[13] : 
                         (N61)? scoreboard_r[14] : 
                         (N63)? scoreboard_r[15] : 
                         (N34)? scoreboard_r[16] : 
                         (N36)? scoreboard_r[17] : 
                         (N38)? scoreboard_r[18] : 
                         (N40)? scoreboard_r[19] : 
                         (N42)? scoreboard_r[20] : 
                         (N44)? scoreboard_r[21] : 
                         (N46)? scoreboard_r[22] : 
                         (N48)? scoreboard_r[23] : 
                         (N50)? scoreboard_r[24] : 
                         (N52)? scoreboard_r[25] : 
                         (N54)? scoreboard_r[26] : 
                         (N56)? scoreboard_r[27] : 
                         (N58)? scoreboard_r[28] : 
                         (N60)? scoreboard_r[29] : 
                         (N62)? scoreboard_r[30] : 
                         (N64)? scoreboard_r[31] : 1'b0;
  assign rs_match_o[1] = (N98)? scoreboard_r[0] : 
                         (N100)? scoreboard_r[1] : 
                         (N102)? scoreboard_r[2] : 
                         (N104)? scoreboard_r[3] : 
                         (N106)? scoreboard_r[4] : 
                         (N108)? scoreboard_r[5] : 
                         (N110)? scoreboard_r[6] : 
                         (N112)? scoreboard_r[7] : 
                         (N114)? scoreboard_r[8] : 
                         (N116)? scoreboard_r[9] : 
                         (N118)? scoreboard_r[10] : 
                         (N120)? scoreboard_r[11] : 
                         (N122)? scoreboard_r[12] : 
                         (N124)? scoreboard_r[13] : 
                         (N126)? scoreboard_r[14] : 
                         (N128)? scoreboard_r[15] : 
                         (N99)? scoreboard_r[16] : 
                         (N101)? scoreboard_r[17] : 
                         (N103)? scoreboard_r[18] : 
                         (N105)? scoreboard_r[19] : 
                         (N107)? scoreboard_r[20] : 
                         (N109)? scoreboard_r[21] : 
                         (N111)? scoreboard_r[22] : 
                         (N113)? scoreboard_r[23] : 
                         (N115)? scoreboard_r[24] : 
                         (N117)? scoreboard_r[25] : 
                         (N119)? scoreboard_r[26] : 
                         (N121)? scoreboard_r[27] : 
                         (N123)? scoreboard_r[28] : 
                         (N125)? scoreboard_r[29] : 
                         (N127)? scoreboard_r[30] : 
                         (N129)? scoreboard_r[31] : 1'b0;
  assign rd_match_o = (N163)? scoreboard_r[0] : 
                      (N165)? scoreboard_r[1] : 
                      (N167)? scoreboard_r[2] : 
                      (N169)? scoreboard_r[3] : 
                      (N171)? scoreboard_r[4] : 
                      (N173)? scoreboard_r[5] : 
                      (N175)? scoreboard_r[6] : 
                      (N177)? scoreboard_r[7] : 
                      (N179)? scoreboard_r[8] : 
                      (N181)? scoreboard_r[9] : 
                      (N183)? scoreboard_r[10] : 
                      (N185)? scoreboard_r[11] : 
                      (N187)? scoreboard_r[12] : 
                      (N189)? scoreboard_r[13] : 
                      (N191)? scoreboard_r[14] : 
                      (N193)? scoreboard_r[15] : 
                      (N164)? scoreboard_r[16] : 
                      (N166)? scoreboard_r[17] : 
                      (N168)? scoreboard_r[18] : 
                      (N170)? scoreboard_r[19] : 
                      (N172)? scoreboard_r[20] : 
                      (N174)? scoreboard_r[21] : 
                      (N176)? scoreboard_r[22] : 
                      (N178)? scoreboard_r[23] : 
                      (N180)? scoreboard_r[24] : 
                      (N182)? scoreboard_r[25] : 
                      (N184)? scoreboard_r[26] : 
                      (N186)? scoreboard_r[27] : 
                      (N188)? scoreboard_r[28] : 
                      (N190)? scoreboard_r[29] : 
                      (N192)? scoreboard_r[30] : 
                      (N194)? scoreboard_r[31] : 1'b0;
  assign N0 = ~check_rs_i[0];
  assign N1 = ~check_rs_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & check_rs_i[1];
  assign N4 = check_rs_i[0] & N1;
  assign N5 = check_rs_i[0] & check_rs_i[1];
  assign N6 = ~check_rs_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & check_rs_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & check_rs_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & check_rs_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & check_rs_i[2];
  assign N15 = ~check_rs_i[3];
  assign N16 = N7 & N15;
  assign N17 = N7 & check_rs_i[3];
  assign N18 = N9 & N15;
  assign N19 = N9 & check_rs_i[3];
  assign N20 = N11 & N15;
  assign N21 = N11 & check_rs_i[3];
  assign N22 = N13 & N15;
  assign N23 = N13 & check_rs_i[3];
  assign N24 = N8 & N15;
  assign N25 = N8 & check_rs_i[3];
  assign N26 = N10 & N15;
  assign N27 = N10 & check_rs_i[3];
  assign N28 = N12 & N15;
  assign N29 = N12 & check_rs_i[3];
  assign N30 = N14 & N15;
  assign N31 = N14 & check_rs_i[3];
  assign N32 = ~check_rs_i[4];
  assign N33 = N16 & N32;
  assign N34 = N16 & check_rs_i[4];
  assign N35 = N18 & N32;
  assign N36 = N18 & check_rs_i[4];
  assign N37 = N20 & N32;
  assign N38 = N20 & check_rs_i[4];
  assign N39 = N22 & N32;
  assign N40 = N22 & check_rs_i[4];
  assign N41 = N24 & N32;
  assign N42 = N24 & check_rs_i[4];
  assign N43 = N26 & N32;
  assign N44 = N26 & check_rs_i[4];
  assign N45 = N28 & N32;
  assign N46 = N28 & check_rs_i[4];
  assign N47 = N30 & N32;
  assign N48 = N30 & check_rs_i[4];
  assign N49 = N17 & N32;
  assign N50 = N17 & check_rs_i[4];
  assign N51 = N19 & N32;
  assign N52 = N19 & check_rs_i[4];
  assign N53 = N21 & N32;
  assign N54 = N21 & check_rs_i[4];
  assign N55 = N23 & N32;
  assign N56 = N23 & check_rs_i[4];
  assign N57 = N25 & N32;
  assign N58 = N25 & check_rs_i[4];
  assign N59 = N27 & N32;
  assign N60 = N27 & check_rs_i[4];
  assign N61 = N29 & N32;
  assign N62 = N29 & check_rs_i[4];
  assign N63 = N31 & N32;
  assign N64 = N31 & check_rs_i[4];
  assign N65 = ~check_rs_i[5];
  assign N66 = ~check_rs_i[6];
  assign N67 = N65 & N66;
  assign N68 = N65 & check_rs_i[6];
  assign N69 = check_rs_i[5] & N66;
  assign N70 = check_rs_i[5] & check_rs_i[6];
  assign N71 = ~check_rs_i[7];
  assign N72 = N67 & N71;
  assign N73 = N67 & check_rs_i[7];
  assign N74 = N69 & N71;
  assign N75 = N69 & check_rs_i[7];
  assign N76 = N68 & N71;
  assign N77 = N68 & check_rs_i[7];
  assign N78 = N70 & N71;
  assign N79 = N70 & check_rs_i[7];
  assign N80 = ~check_rs_i[8];
  assign N81 = N72 & N80;
  assign N82 = N72 & check_rs_i[8];
  assign N83 = N74 & N80;
  assign N84 = N74 & check_rs_i[8];
  assign N85 = N76 & N80;
  assign N86 = N76 & check_rs_i[8];
  assign N87 = N78 & N80;
  assign N88 = N78 & check_rs_i[8];
  assign N89 = N73 & N80;
  assign N90 = N73 & check_rs_i[8];
  assign N91 = N75 & N80;
  assign N92 = N75 & check_rs_i[8];
  assign N93 = N77 & N80;
  assign N94 = N77 & check_rs_i[8];
  assign N95 = N79 & N80;
  assign N96 = N79 & check_rs_i[8];
  assign N97 = ~check_rs_i[9];
  assign N98 = N81 & N97;
  assign N99 = N81 & check_rs_i[9];
  assign N100 = N83 & N97;
  assign N101 = N83 & check_rs_i[9];
  assign N102 = N85 & N97;
  assign N103 = N85 & check_rs_i[9];
  assign N104 = N87 & N97;
  assign N105 = N87 & check_rs_i[9];
  assign N106 = N89 & N97;
  assign N107 = N89 & check_rs_i[9];
  assign N108 = N91 & N97;
  assign N109 = N91 & check_rs_i[9];
  assign N110 = N93 & N97;
  assign N111 = N93 & check_rs_i[9];
  assign N112 = N95 & N97;
  assign N113 = N95 & check_rs_i[9];
  assign N114 = N82 & N97;
  assign N115 = N82 & check_rs_i[9];
  assign N116 = N84 & N97;
  assign N117 = N84 & check_rs_i[9];
  assign N118 = N86 & N97;
  assign N119 = N86 & check_rs_i[9];
  assign N120 = N88 & N97;
  assign N121 = N88 & check_rs_i[9];
  assign N122 = N90 & N97;
  assign N123 = N90 & check_rs_i[9];
  assign N124 = N92 & N97;
  assign N125 = N92 & check_rs_i[9];
  assign N126 = N94 & N97;
  assign N127 = N94 & check_rs_i[9];
  assign N128 = N96 & N97;
  assign N129 = N96 & check_rs_i[9];
  assign N130 = ~check_rd_i[0];
  assign N131 = ~check_rd_i[1];
  assign N132 = N130 & N131;
  assign N133 = N130 & check_rd_i[1];
  assign N134 = check_rd_i[0] & N131;
  assign N135 = check_rd_i[0] & check_rd_i[1];
  assign N136 = ~check_rd_i[2];
  assign N137 = N132 & N136;
  assign N138 = N132 & check_rd_i[2];
  assign N139 = N134 & N136;
  assign N140 = N134 & check_rd_i[2];
  assign N141 = N133 & N136;
  assign N142 = N133 & check_rd_i[2];
  assign N143 = N135 & N136;
  assign N144 = N135 & check_rd_i[2];
  assign N145 = ~check_rd_i[3];
  assign N146 = N137 & N145;
  assign N147 = N137 & check_rd_i[3];
  assign N148 = N139 & N145;
  assign N149 = N139 & check_rd_i[3];
  assign N150 = N141 & N145;
  assign N151 = N141 & check_rd_i[3];
  assign N152 = N143 & N145;
  assign N153 = N143 & check_rd_i[3];
  assign N154 = N138 & N145;
  assign N155 = N138 & check_rd_i[3];
  assign N156 = N140 & N145;
  assign N157 = N140 & check_rd_i[3];
  assign N158 = N142 & N145;
  assign N159 = N142 & check_rd_i[3];
  assign N160 = N144 & N145;
  assign N161 = N144 & check_rd_i[3];
  assign N162 = ~check_rd_i[4];
  assign N163 = N146 & N162;
  assign N164 = N146 & check_rd_i[4];
  assign N165 = N148 & N162;
  assign N166 = N148 & check_rd_i[4];
  assign N167 = N150 & N162;
  assign N168 = N150 & check_rd_i[4];
  assign N169 = N152 & N162;
  assign N170 = N152 & check_rd_i[4];
  assign N171 = N154 & N162;
  assign N172 = N154 & check_rd_i[4];
  assign N173 = N156 & N162;
  assign N174 = N156 & check_rd_i[4];
  assign N175 = N158 & N162;
  assign N176 = N158 & check_rd_i[4];
  assign N177 = N160 & N162;
  assign N178 = N160 & check_rd_i[4];
  assign N179 = N147 & N162;
  assign N180 = N147 & check_rd_i[4];
  assign N181 = N149 & N162;
  assign N182 = N149 & check_rd_i[4];
  assign N183 = N151 & N162;
  assign N184 = N151 & check_rd_i[4];
  assign N185 = N153 & N162;
  assign N186 = N153 & check_rd_i[4];
  assign N187 = N155 & N162;
  assign N188 = N155 & check_rd_i[4];
  assign N189 = N157 & N162;
  assign N190 = N157 & check_rd_i[4];
  assign N191 = N159 & N162;
  assign N192 = N159 & check_rd_i[4];
  assign N193 = N161 & N162;
  assign N194 = N161 & check_rd_i[4];

endmodule



module bp_be_scoreboard_00_3
(
  clk_i,
  reset_i,
  score_v_i,
  score_rd_i,
  clear_v_i,
  clear_rd_i,
  check_rs_i,
  check_rd_i,
  rs_match_o,
  rd_match_o
);

  input [4:0] score_rd_i;
  input [4:0] clear_rd_i;
  input [14:0] check_rs_i;
  input [4:0] check_rd_i;
  output [2:0] rs_match_o;
  input clk_i;
  input reset_i;
  input score_v_i;
  input clear_v_i;
  output rd_match_o;
  wire [2:0] rs_match_o;
  wire rd_match_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,
  N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,
  N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,
  N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,
  N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,
  N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
  N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,
  N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,
  N259;
  wire [31:0] score_onehot_li,clear_onehot_li,scoreboard_r;

  bsg_decode_with_v_num_out_p32
  score_decode
  (
    .i(score_rd_i),
    .v_i(score_v_i),
    .o(score_onehot_li)
  );


  bsg_decode_with_v_num_out_p32
  clear_decode
  (
    .i(clear_rd_i),
    .v_i(clear_v_i),
    .o(clear_onehot_li)
  );


  bsg_dff_reset_set_clear_width_p32_clear_over_set_p1
  scoreboard_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .set_i(score_onehot_li),
    .clear_i(clear_onehot_li),
    .data_o(scoreboard_r)
  );

  assign rs_match_o[0] = (N33)? scoreboard_r[0] : 
                         (N35)? scoreboard_r[1] : 
                         (N37)? scoreboard_r[2] : 
                         (N39)? scoreboard_r[3] : 
                         (N41)? scoreboard_r[4] : 
                         (N43)? scoreboard_r[5] : 
                         (N45)? scoreboard_r[6] : 
                         (N47)? scoreboard_r[7] : 
                         (N49)? scoreboard_r[8] : 
                         (N51)? scoreboard_r[9] : 
                         (N53)? scoreboard_r[10] : 
                         (N55)? scoreboard_r[11] : 
                         (N57)? scoreboard_r[12] : 
                         (N59)? scoreboard_r[13] : 
                         (N61)? scoreboard_r[14] : 
                         (N63)? scoreboard_r[15] : 
                         (N34)? scoreboard_r[16] : 
                         (N36)? scoreboard_r[17] : 
                         (N38)? scoreboard_r[18] : 
                         (N40)? scoreboard_r[19] : 
                         (N42)? scoreboard_r[20] : 
                         (N44)? scoreboard_r[21] : 
                         (N46)? scoreboard_r[22] : 
                         (N48)? scoreboard_r[23] : 
                         (N50)? scoreboard_r[24] : 
                         (N52)? scoreboard_r[25] : 
                         (N54)? scoreboard_r[26] : 
                         (N56)? scoreboard_r[27] : 
                         (N58)? scoreboard_r[28] : 
                         (N60)? scoreboard_r[29] : 
                         (N62)? scoreboard_r[30] : 
                         (N64)? scoreboard_r[31] : 1'b0;
  assign rs_match_o[1] = (N98)? scoreboard_r[0] : 
                         (N100)? scoreboard_r[1] : 
                         (N102)? scoreboard_r[2] : 
                         (N104)? scoreboard_r[3] : 
                         (N106)? scoreboard_r[4] : 
                         (N108)? scoreboard_r[5] : 
                         (N110)? scoreboard_r[6] : 
                         (N112)? scoreboard_r[7] : 
                         (N114)? scoreboard_r[8] : 
                         (N116)? scoreboard_r[9] : 
                         (N118)? scoreboard_r[10] : 
                         (N120)? scoreboard_r[11] : 
                         (N122)? scoreboard_r[12] : 
                         (N124)? scoreboard_r[13] : 
                         (N126)? scoreboard_r[14] : 
                         (N128)? scoreboard_r[15] : 
                         (N99)? scoreboard_r[16] : 
                         (N101)? scoreboard_r[17] : 
                         (N103)? scoreboard_r[18] : 
                         (N105)? scoreboard_r[19] : 
                         (N107)? scoreboard_r[20] : 
                         (N109)? scoreboard_r[21] : 
                         (N111)? scoreboard_r[22] : 
                         (N113)? scoreboard_r[23] : 
                         (N115)? scoreboard_r[24] : 
                         (N117)? scoreboard_r[25] : 
                         (N119)? scoreboard_r[26] : 
                         (N121)? scoreboard_r[27] : 
                         (N123)? scoreboard_r[28] : 
                         (N125)? scoreboard_r[29] : 
                         (N127)? scoreboard_r[30] : 
                         (N129)? scoreboard_r[31] : 1'b0;
  assign rs_match_o[2] = (N163)? scoreboard_r[0] : 
                         (N165)? scoreboard_r[1] : 
                         (N167)? scoreboard_r[2] : 
                         (N169)? scoreboard_r[3] : 
                         (N171)? scoreboard_r[4] : 
                         (N173)? scoreboard_r[5] : 
                         (N175)? scoreboard_r[6] : 
                         (N177)? scoreboard_r[7] : 
                         (N179)? scoreboard_r[8] : 
                         (N181)? scoreboard_r[9] : 
                         (N183)? scoreboard_r[10] : 
                         (N185)? scoreboard_r[11] : 
                         (N187)? scoreboard_r[12] : 
                         (N189)? scoreboard_r[13] : 
                         (N191)? scoreboard_r[14] : 
                         (N193)? scoreboard_r[15] : 
                         (N164)? scoreboard_r[16] : 
                         (N166)? scoreboard_r[17] : 
                         (N168)? scoreboard_r[18] : 
                         (N170)? scoreboard_r[19] : 
                         (N172)? scoreboard_r[20] : 
                         (N174)? scoreboard_r[21] : 
                         (N176)? scoreboard_r[22] : 
                         (N178)? scoreboard_r[23] : 
                         (N180)? scoreboard_r[24] : 
                         (N182)? scoreboard_r[25] : 
                         (N184)? scoreboard_r[26] : 
                         (N186)? scoreboard_r[27] : 
                         (N188)? scoreboard_r[28] : 
                         (N190)? scoreboard_r[29] : 
                         (N192)? scoreboard_r[30] : 
                         (N194)? scoreboard_r[31] : 1'b0;
  assign rd_match_o = (N228)? scoreboard_r[0] : 
                      (N230)? scoreboard_r[1] : 
                      (N232)? scoreboard_r[2] : 
                      (N234)? scoreboard_r[3] : 
                      (N236)? scoreboard_r[4] : 
                      (N238)? scoreboard_r[5] : 
                      (N240)? scoreboard_r[6] : 
                      (N242)? scoreboard_r[7] : 
                      (N244)? scoreboard_r[8] : 
                      (N246)? scoreboard_r[9] : 
                      (N248)? scoreboard_r[10] : 
                      (N250)? scoreboard_r[11] : 
                      (N252)? scoreboard_r[12] : 
                      (N254)? scoreboard_r[13] : 
                      (N256)? scoreboard_r[14] : 
                      (N258)? scoreboard_r[15] : 
                      (N229)? scoreboard_r[16] : 
                      (N231)? scoreboard_r[17] : 
                      (N233)? scoreboard_r[18] : 
                      (N235)? scoreboard_r[19] : 
                      (N237)? scoreboard_r[20] : 
                      (N239)? scoreboard_r[21] : 
                      (N241)? scoreboard_r[22] : 
                      (N243)? scoreboard_r[23] : 
                      (N245)? scoreboard_r[24] : 
                      (N247)? scoreboard_r[25] : 
                      (N249)? scoreboard_r[26] : 
                      (N251)? scoreboard_r[27] : 
                      (N253)? scoreboard_r[28] : 
                      (N255)? scoreboard_r[29] : 
                      (N257)? scoreboard_r[30] : 
                      (N259)? scoreboard_r[31] : 1'b0;
  assign N0 = ~check_rs_i[0];
  assign N1 = ~check_rs_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & check_rs_i[1];
  assign N4 = check_rs_i[0] & N1;
  assign N5 = check_rs_i[0] & check_rs_i[1];
  assign N6 = ~check_rs_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & check_rs_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & check_rs_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & check_rs_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & check_rs_i[2];
  assign N15 = ~check_rs_i[3];
  assign N16 = N7 & N15;
  assign N17 = N7 & check_rs_i[3];
  assign N18 = N9 & N15;
  assign N19 = N9 & check_rs_i[3];
  assign N20 = N11 & N15;
  assign N21 = N11 & check_rs_i[3];
  assign N22 = N13 & N15;
  assign N23 = N13 & check_rs_i[3];
  assign N24 = N8 & N15;
  assign N25 = N8 & check_rs_i[3];
  assign N26 = N10 & N15;
  assign N27 = N10 & check_rs_i[3];
  assign N28 = N12 & N15;
  assign N29 = N12 & check_rs_i[3];
  assign N30 = N14 & N15;
  assign N31 = N14 & check_rs_i[3];
  assign N32 = ~check_rs_i[4];
  assign N33 = N16 & N32;
  assign N34 = N16 & check_rs_i[4];
  assign N35 = N18 & N32;
  assign N36 = N18 & check_rs_i[4];
  assign N37 = N20 & N32;
  assign N38 = N20 & check_rs_i[4];
  assign N39 = N22 & N32;
  assign N40 = N22 & check_rs_i[4];
  assign N41 = N24 & N32;
  assign N42 = N24 & check_rs_i[4];
  assign N43 = N26 & N32;
  assign N44 = N26 & check_rs_i[4];
  assign N45 = N28 & N32;
  assign N46 = N28 & check_rs_i[4];
  assign N47 = N30 & N32;
  assign N48 = N30 & check_rs_i[4];
  assign N49 = N17 & N32;
  assign N50 = N17 & check_rs_i[4];
  assign N51 = N19 & N32;
  assign N52 = N19 & check_rs_i[4];
  assign N53 = N21 & N32;
  assign N54 = N21 & check_rs_i[4];
  assign N55 = N23 & N32;
  assign N56 = N23 & check_rs_i[4];
  assign N57 = N25 & N32;
  assign N58 = N25 & check_rs_i[4];
  assign N59 = N27 & N32;
  assign N60 = N27 & check_rs_i[4];
  assign N61 = N29 & N32;
  assign N62 = N29 & check_rs_i[4];
  assign N63 = N31 & N32;
  assign N64 = N31 & check_rs_i[4];
  assign N65 = ~check_rs_i[5];
  assign N66 = ~check_rs_i[6];
  assign N67 = N65 & N66;
  assign N68 = N65 & check_rs_i[6];
  assign N69 = check_rs_i[5] & N66;
  assign N70 = check_rs_i[5] & check_rs_i[6];
  assign N71 = ~check_rs_i[7];
  assign N72 = N67 & N71;
  assign N73 = N67 & check_rs_i[7];
  assign N74 = N69 & N71;
  assign N75 = N69 & check_rs_i[7];
  assign N76 = N68 & N71;
  assign N77 = N68 & check_rs_i[7];
  assign N78 = N70 & N71;
  assign N79 = N70 & check_rs_i[7];
  assign N80 = ~check_rs_i[8];
  assign N81 = N72 & N80;
  assign N82 = N72 & check_rs_i[8];
  assign N83 = N74 & N80;
  assign N84 = N74 & check_rs_i[8];
  assign N85 = N76 & N80;
  assign N86 = N76 & check_rs_i[8];
  assign N87 = N78 & N80;
  assign N88 = N78 & check_rs_i[8];
  assign N89 = N73 & N80;
  assign N90 = N73 & check_rs_i[8];
  assign N91 = N75 & N80;
  assign N92 = N75 & check_rs_i[8];
  assign N93 = N77 & N80;
  assign N94 = N77 & check_rs_i[8];
  assign N95 = N79 & N80;
  assign N96 = N79 & check_rs_i[8];
  assign N97 = ~check_rs_i[9];
  assign N98 = N81 & N97;
  assign N99 = N81 & check_rs_i[9];
  assign N100 = N83 & N97;
  assign N101 = N83 & check_rs_i[9];
  assign N102 = N85 & N97;
  assign N103 = N85 & check_rs_i[9];
  assign N104 = N87 & N97;
  assign N105 = N87 & check_rs_i[9];
  assign N106 = N89 & N97;
  assign N107 = N89 & check_rs_i[9];
  assign N108 = N91 & N97;
  assign N109 = N91 & check_rs_i[9];
  assign N110 = N93 & N97;
  assign N111 = N93 & check_rs_i[9];
  assign N112 = N95 & N97;
  assign N113 = N95 & check_rs_i[9];
  assign N114 = N82 & N97;
  assign N115 = N82 & check_rs_i[9];
  assign N116 = N84 & N97;
  assign N117 = N84 & check_rs_i[9];
  assign N118 = N86 & N97;
  assign N119 = N86 & check_rs_i[9];
  assign N120 = N88 & N97;
  assign N121 = N88 & check_rs_i[9];
  assign N122 = N90 & N97;
  assign N123 = N90 & check_rs_i[9];
  assign N124 = N92 & N97;
  assign N125 = N92 & check_rs_i[9];
  assign N126 = N94 & N97;
  assign N127 = N94 & check_rs_i[9];
  assign N128 = N96 & N97;
  assign N129 = N96 & check_rs_i[9];
  assign N130 = ~check_rs_i[10];
  assign N131 = ~check_rs_i[11];
  assign N132 = N130 & N131;
  assign N133 = N130 & check_rs_i[11];
  assign N134 = check_rs_i[10] & N131;
  assign N135 = check_rs_i[10] & check_rs_i[11];
  assign N136 = ~check_rs_i[12];
  assign N137 = N132 & N136;
  assign N138 = N132 & check_rs_i[12];
  assign N139 = N134 & N136;
  assign N140 = N134 & check_rs_i[12];
  assign N141 = N133 & N136;
  assign N142 = N133 & check_rs_i[12];
  assign N143 = N135 & N136;
  assign N144 = N135 & check_rs_i[12];
  assign N145 = ~check_rs_i[13];
  assign N146 = N137 & N145;
  assign N147 = N137 & check_rs_i[13];
  assign N148 = N139 & N145;
  assign N149 = N139 & check_rs_i[13];
  assign N150 = N141 & N145;
  assign N151 = N141 & check_rs_i[13];
  assign N152 = N143 & N145;
  assign N153 = N143 & check_rs_i[13];
  assign N154 = N138 & N145;
  assign N155 = N138 & check_rs_i[13];
  assign N156 = N140 & N145;
  assign N157 = N140 & check_rs_i[13];
  assign N158 = N142 & N145;
  assign N159 = N142 & check_rs_i[13];
  assign N160 = N144 & N145;
  assign N161 = N144 & check_rs_i[13];
  assign N162 = ~check_rs_i[14];
  assign N163 = N146 & N162;
  assign N164 = N146 & check_rs_i[14];
  assign N165 = N148 & N162;
  assign N166 = N148 & check_rs_i[14];
  assign N167 = N150 & N162;
  assign N168 = N150 & check_rs_i[14];
  assign N169 = N152 & N162;
  assign N170 = N152 & check_rs_i[14];
  assign N171 = N154 & N162;
  assign N172 = N154 & check_rs_i[14];
  assign N173 = N156 & N162;
  assign N174 = N156 & check_rs_i[14];
  assign N175 = N158 & N162;
  assign N176 = N158 & check_rs_i[14];
  assign N177 = N160 & N162;
  assign N178 = N160 & check_rs_i[14];
  assign N179 = N147 & N162;
  assign N180 = N147 & check_rs_i[14];
  assign N181 = N149 & N162;
  assign N182 = N149 & check_rs_i[14];
  assign N183 = N151 & N162;
  assign N184 = N151 & check_rs_i[14];
  assign N185 = N153 & N162;
  assign N186 = N153 & check_rs_i[14];
  assign N187 = N155 & N162;
  assign N188 = N155 & check_rs_i[14];
  assign N189 = N157 & N162;
  assign N190 = N157 & check_rs_i[14];
  assign N191 = N159 & N162;
  assign N192 = N159 & check_rs_i[14];
  assign N193 = N161 & N162;
  assign N194 = N161 & check_rs_i[14];
  assign N195 = ~check_rd_i[0];
  assign N196 = ~check_rd_i[1];
  assign N197 = N195 & N196;
  assign N198 = N195 & check_rd_i[1];
  assign N199 = check_rd_i[0] & N196;
  assign N200 = check_rd_i[0] & check_rd_i[1];
  assign N201 = ~check_rd_i[2];
  assign N202 = N197 & N201;
  assign N203 = N197 & check_rd_i[2];
  assign N204 = N199 & N201;
  assign N205 = N199 & check_rd_i[2];
  assign N206 = N198 & N201;
  assign N207 = N198 & check_rd_i[2];
  assign N208 = N200 & N201;
  assign N209 = N200 & check_rd_i[2];
  assign N210 = ~check_rd_i[3];
  assign N211 = N202 & N210;
  assign N212 = N202 & check_rd_i[3];
  assign N213 = N204 & N210;
  assign N214 = N204 & check_rd_i[3];
  assign N215 = N206 & N210;
  assign N216 = N206 & check_rd_i[3];
  assign N217 = N208 & N210;
  assign N218 = N208 & check_rd_i[3];
  assign N219 = N203 & N210;
  assign N220 = N203 & check_rd_i[3];
  assign N221 = N205 & N210;
  assign N222 = N205 & check_rd_i[3];
  assign N223 = N207 & N210;
  assign N224 = N207 & check_rd_i[3];
  assign N225 = N209 & N210;
  assign N226 = N209 & check_rd_i[3];
  assign N227 = ~check_rd_i[4];
  assign N228 = N211 & N227;
  assign N229 = N211 & check_rd_i[4];
  assign N230 = N213 & N227;
  assign N231 = N213 & check_rd_i[4];
  assign N232 = N215 & N227;
  assign N233 = N215 & check_rd_i[4];
  assign N234 = N217 & N227;
  assign N235 = N217 & check_rd_i[4];
  assign N236 = N219 & N227;
  assign N237 = N219 & check_rd_i[4];
  assign N238 = N221 & N227;
  assign N239 = N221 & check_rd_i[4];
  assign N240 = N223 & N227;
  assign N241 = N223 & check_rd_i[4];
  assign N242 = N225 & N227;
  assign N243 = N225 & check_rd_i[4];
  assign N244 = N212 & N227;
  assign N245 = N212 & check_rd_i[4];
  assign N246 = N214 & N227;
  assign N247 = N214 & check_rd_i[4];
  assign N248 = N216 & N227;
  assign N249 = N216 & check_rd_i[4];
  assign N250 = N218 & N227;
  assign N251 = N218 & check_rd_i[4];
  assign N252 = N220 & N227;
  assign N253 = N220 & check_rd_i[4];
  assign N254 = N222 & N227;
  assign N255 = N222 & check_rd_i[4];
  assign N256 = N224 & N227;
  assign N257 = N224 & check_rd_i[4];
  assign N258 = N226 & N227;
  assign N259 = N226 & check_rd_i[4];

endmodule



module bp_be_detector_00
(
  clk_i,
  reset_i,
  issue_pkt_i,
  cmd_full_i,
  credits_full_i,
  credits_empty_i,
  idiv_busy_i,
  fdiv_busy_i,
  mem_busy_i,
  mem_ordered_i,
  hazard_v_o,
  ordered_v_o,
  dispatch_pkt_i,
  commit_pkt_i,
  late_wb_pkt_i,
  late_wb_yumi_i,
  ispec_v_o
);

  input [263:0] issue_pkt_i;
  input [365:0] dispatch_pkt_i;
  input [213:0] commit_pkt_i;
  input [78:0] late_wb_pkt_i;
  input clk_i;
  input reset_i;
  input cmd_full_i;
  input credits_full_i;
  input credits_empty_i;
  input idiv_busy_i;
  input fdiv_busy_i;
  input mem_busy_i;
  input mem_ordered_i;
  input late_wb_yumi_i;
  output hazard_v_o;
  output ordered_v_o;
  output ispec_v_o;
  wire hazard_v_o,ordered_v_o,ispec_v_o,N0,dep_status_r_3__fflags_v_,
  dep_status_r_2__fflags_v_,dep_status_r_2__fma_fwb_v_,dep_status_r_2__long_iwb_v_,
  dep_status_r_2__long_fwb_v_,dep_status_r_2__rd_addr__4_,dep_status_r_2__rd_addr__3_,
  dep_status_r_2__rd_addr__2_,dep_status_r_2__rd_addr__1_,dep_status_r_2__rd_addr__0_,
  dep_status_r_1__fflags_v_,dep_status_r_1__fmem_iwb_v_,dep_status_r_1__fmem_fwb_v_,
  dep_status_r_1__mul_iwb_v_,dep_status_r_1__fma_fwb_v_,dep_status_r_1__long_iwb_v_,
  dep_status_r_1__long_fwb_v_,dep_status_r_1__rd_addr__4_,dep_status_r_1__rd_addr__3_,
  dep_status_r_1__rd_addr__2_,dep_status_r_1__rd_addr__1_,
  dep_status_r_1__rd_addr__0_,dep_status_r_0__fflags_v_,dep_status_r_0__aux_iwb_v_,
  dep_status_r_0__aux_fwb_v_,dep_status_r_0__fint_iwb_v_,dep_status_r_0__fint_fwb_v_,
  dep_status_r_0__emem_iwb_v_,dep_status_r_0__emem_fwb_v_,dep_status_r_0__fmem_iwb_v_,
  dep_status_r_0__fmem_fwb_v_,dep_status_r_0__mul_iwb_v_,dep_status_r_0__fma_fwb_v_,
  dep_status_r_0__long_iwb_v_,dep_status_r_0__long_fwb_v_,dep_status_r_0__rd_addr__4_,
  dep_status_r_0__rd_addr__3_,dep_status_r_0__rd_addr__2_,dep_status_r_0__rd_addr__1_,
  dep_status_r_0__rd_addr__0_,irs1_ispec_v,irs2_ispec_v,irs2_store_v,clear_int_v_li,
  ird_match_lo,clear_fp_v_li,frd_match_lo,irs1_sb_raw_haz_v,irs2_sb_raw_haz_v,
  ird_sb_waw_haz_v,frs1_sb_raw_haz_v,frs2_sb_raw_haz_v,frs3_sb_raw_haz_v,frd_sb_waw_haz_v,
  iscore_haz_v,fscore_haz_v,fence_haz_v,fflags_haz_v,control_haz_v,data_haz_v,
  struct_haz_v,dep_status_n_fflags_v_,dep_status_n_aux_iwb_v_,dep_status_n_aux_fwb_v_,
  dep_status_n_fint_iwb_v_,dep_status_n_fint_fwb_v_,dep_status_n_emem_iwb_v_,
  dep_status_n_emem_fwb_v_,dep_status_n_fmem_iwb_v_,dep_status_n_fmem_fwb_v_,
  dep_status_n_mul_iwb_v_,dep_status_n_fma_fwb_v_,dep_status_n_long_iwb_v_,
  dep_status_n_long_fwb_v_,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,
  N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,
  N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,
  N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145;
  wire [2:0] rs1_match_vector,rs2_match_vector,frs_match_lo,rs3_match_vector,rd_match_vector,
  irs1_data_haz_v,irs2_data_haz_v,frs1_data_haz_v,frs2_data_haz_v,frs3_data_haz_v;
  wire [1:0] irs_match_lo;
  reg dep_status_r_3__fflags_v__sv2v_reg,dep_status_r_2__fflags_v__sv2v_reg,
  dep_status_r_2__fma_fwb_v__sv2v_reg,dep_status_r_2__long_iwb_v__sv2v_reg,
  dep_status_r_2__long_fwb_v__sv2v_reg,dep_status_r_2__rd_addr__4__sv2v_reg,
  dep_status_r_2__rd_addr__3__sv2v_reg,dep_status_r_2__rd_addr__2__sv2v_reg,
  dep_status_r_2__rd_addr__1__sv2v_reg,dep_status_r_2__rd_addr__0__sv2v_reg,dep_status_r_1__fflags_v__sv2v_reg,
  dep_status_r_1__fmem_iwb_v__sv2v_reg,dep_status_r_1__fmem_fwb_v__sv2v_reg,
  dep_status_r_1__mul_iwb_v__sv2v_reg,dep_status_r_1__fma_fwb_v__sv2v_reg,
  dep_status_r_1__long_iwb_v__sv2v_reg,dep_status_r_1__long_fwb_v__sv2v_reg,
  dep_status_r_1__rd_addr__4__sv2v_reg,dep_status_r_1__rd_addr__3__sv2v_reg,
  dep_status_r_1__rd_addr__2__sv2v_reg,dep_status_r_1__rd_addr__1__sv2v_reg,
  dep_status_r_1__rd_addr__0__sv2v_reg,dep_status_r_0__fflags_v__sv2v_reg,dep_status_r_0__aux_iwb_v__sv2v_reg,
  dep_status_r_0__aux_fwb_v__sv2v_reg,dep_status_r_0__fint_iwb_v__sv2v_reg,
  dep_status_r_0__fint_fwb_v__sv2v_reg,dep_status_r_0__emem_iwb_v__sv2v_reg,
  dep_status_r_0__emem_fwb_v__sv2v_reg,dep_status_r_0__fmem_iwb_v__sv2v_reg,
  dep_status_r_0__fmem_fwb_v__sv2v_reg,dep_status_r_0__mul_iwb_v__sv2v_reg,
  dep_status_r_0__fma_fwb_v__sv2v_reg,dep_status_r_0__long_iwb_v__sv2v_reg,dep_status_r_0__long_fwb_v__sv2v_reg,
  dep_status_r_0__rd_addr__4__sv2v_reg,dep_status_r_0__rd_addr__3__sv2v_reg,
  dep_status_r_0__rd_addr__2__sv2v_reg,dep_status_r_0__rd_addr__1__sv2v_reg,
  dep_status_r_0__rd_addr__0__sv2v_reg;
  assign dep_status_r_3__fflags_v_ = dep_status_r_3__fflags_v__sv2v_reg;
  assign dep_status_r_2__fflags_v_ = dep_status_r_2__fflags_v__sv2v_reg;
  assign dep_status_r_2__fma_fwb_v_ = dep_status_r_2__fma_fwb_v__sv2v_reg;
  assign dep_status_r_2__long_iwb_v_ = dep_status_r_2__long_iwb_v__sv2v_reg;
  assign dep_status_r_2__long_fwb_v_ = dep_status_r_2__long_fwb_v__sv2v_reg;
  assign dep_status_r_2__rd_addr__4_ = dep_status_r_2__rd_addr__4__sv2v_reg;
  assign dep_status_r_2__rd_addr__3_ = dep_status_r_2__rd_addr__3__sv2v_reg;
  assign dep_status_r_2__rd_addr__2_ = dep_status_r_2__rd_addr__2__sv2v_reg;
  assign dep_status_r_2__rd_addr__1_ = dep_status_r_2__rd_addr__1__sv2v_reg;
  assign dep_status_r_2__rd_addr__0_ = dep_status_r_2__rd_addr__0__sv2v_reg;
  assign dep_status_r_1__fflags_v_ = dep_status_r_1__fflags_v__sv2v_reg;
  assign dep_status_r_1__fmem_iwb_v_ = dep_status_r_1__fmem_iwb_v__sv2v_reg;
  assign dep_status_r_1__fmem_fwb_v_ = dep_status_r_1__fmem_fwb_v__sv2v_reg;
  assign dep_status_r_1__mul_iwb_v_ = dep_status_r_1__mul_iwb_v__sv2v_reg;
  assign dep_status_r_1__fma_fwb_v_ = dep_status_r_1__fma_fwb_v__sv2v_reg;
  assign dep_status_r_1__long_iwb_v_ = dep_status_r_1__long_iwb_v__sv2v_reg;
  assign dep_status_r_1__long_fwb_v_ = dep_status_r_1__long_fwb_v__sv2v_reg;
  assign dep_status_r_1__rd_addr__4_ = dep_status_r_1__rd_addr__4__sv2v_reg;
  assign dep_status_r_1__rd_addr__3_ = dep_status_r_1__rd_addr__3__sv2v_reg;
  assign dep_status_r_1__rd_addr__2_ = dep_status_r_1__rd_addr__2__sv2v_reg;
  assign dep_status_r_1__rd_addr__1_ = dep_status_r_1__rd_addr__1__sv2v_reg;
  assign dep_status_r_1__rd_addr__0_ = dep_status_r_1__rd_addr__0__sv2v_reg;
  assign dep_status_r_0__fflags_v_ = dep_status_r_0__fflags_v__sv2v_reg;
  assign dep_status_r_0__aux_iwb_v_ = dep_status_r_0__aux_iwb_v__sv2v_reg;
  assign dep_status_r_0__aux_fwb_v_ = dep_status_r_0__aux_fwb_v__sv2v_reg;
  assign dep_status_r_0__fint_iwb_v_ = dep_status_r_0__fint_iwb_v__sv2v_reg;
  assign dep_status_r_0__fint_fwb_v_ = dep_status_r_0__fint_fwb_v__sv2v_reg;
  assign dep_status_r_0__emem_iwb_v_ = dep_status_r_0__emem_iwb_v__sv2v_reg;
  assign dep_status_r_0__emem_fwb_v_ = dep_status_r_0__emem_fwb_v__sv2v_reg;
  assign dep_status_r_0__fmem_iwb_v_ = dep_status_r_0__fmem_iwb_v__sv2v_reg;
  assign dep_status_r_0__fmem_fwb_v_ = dep_status_r_0__fmem_fwb_v__sv2v_reg;
  assign dep_status_r_0__mul_iwb_v_ = dep_status_r_0__mul_iwb_v__sv2v_reg;
  assign dep_status_r_0__fma_fwb_v_ = dep_status_r_0__fma_fwb_v__sv2v_reg;
  assign dep_status_r_0__long_iwb_v_ = dep_status_r_0__long_iwb_v__sv2v_reg;
  assign dep_status_r_0__long_fwb_v_ = dep_status_r_0__long_fwb_v__sv2v_reg;
  assign dep_status_r_0__rd_addr__4_ = dep_status_r_0__rd_addr__4__sv2v_reg;
  assign dep_status_r_0__rd_addr__3_ = dep_status_r_0__rd_addr__3__sv2v_reg;
  assign dep_status_r_0__rd_addr__2_ = dep_status_r_0__rd_addr__2__sv2v_reg;
  assign dep_status_r_0__rd_addr__1_ = dep_status_r_0__rd_addr__1__sv2v_reg;
  assign dep_status_r_0__rd_addr__0_ = dep_status_r_0__rd_addr__0__sv2v_reg;

  bp_be_scoreboard_00_2
  int_scoreboard
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .score_v_i(commit_pkt_i[1]),
    .score_rd_i(commit_pkt_i[68:64]),
    .clear_v_i(clear_int_v_li),
    .clear_rd_i(late_wb_pkt_i[75:71]),
    .check_rs_i(issue_pkt_i[198:189]),
    .check_rd_i(issue_pkt_i[185:181]),
    .rs_match_o(irs_match_lo),
    .rd_match_o(ird_match_lo)
  );


  bp_be_scoreboard_00_3
  fp_scoreboard
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .score_v_i(commit_pkt_i[0]),
    .score_rd_i(commit_pkt_i[68:64]),
    .clear_v_i(clear_fp_v_li),
    .clear_rd_i(late_wb_pkt_i[75:71]),
    .check_rs_i({ issue_pkt_i[205:201], issue_pkt_i[198:189] }),
    .check_rd_i(issue_pkt_i[185:181]),
    .rs_match_o(frs_match_lo),
    .rd_match_o(frd_match_lo)
  );

  assign rs1_match_vector[0] = issue_pkt_i[193:189] == { dep_status_r_0__rd_addr__4_, dep_status_r_0__rd_addr__3_, dep_status_r_0__rd_addr__2_, dep_status_r_0__rd_addr__1_, dep_status_r_0__rd_addr__0_ };
  assign rs2_match_vector[0] = issue_pkt_i[198:194] == { dep_status_r_0__rd_addr__4_, dep_status_r_0__rd_addr__3_, dep_status_r_0__rd_addr__2_, dep_status_r_0__rd_addr__1_, dep_status_r_0__rd_addr__0_ };
  assign rs3_match_vector[0] = issue_pkt_i[205:201] == { dep_status_r_0__rd_addr__4_, dep_status_r_0__rd_addr__3_, dep_status_r_0__rd_addr__2_, dep_status_r_0__rd_addr__1_, dep_status_r_0__rd_addr__0_ };
  assign rd_match_vector[0] = issue_pkt_i[185:181] == { dep_status_r_0__rd_addr__4_, dep_status_r_0__rd_addr__3_, dep_status_r_0__rd_addr__2_, dep_status_r_0__rd_addr__1_, dep_status_r_0__rd_addr__0_ };
  assign rs1_match_vector[1] = issue_pkt_i[193:189] == { dep_status_r_1__rd_addr__4_, dep_status_r_1__rd_addr__3_, dep_status_r_1__rd_addr__2_, dep_status_r_1__rd_addr__1_, dep_status_r_1__rd_addr__0_ };
  assign rs2_match_vector[1] = issue_pkt_i[198:194] == { dep_status_r_1__rd_addr__4_, dep_status_r_1__rd_addr__3_, dep_status_r_1__rd_addr__2_, dep_status_r_1__rd_addr__1_, dep_status_r_1__rd_addr__0_ };
  assign rs3_match_vector[1] = issue_pkt_i[205:201] == { dep_status_r_1__rd_addr__4_, dep_status_r_1__rd_addr__3_, dep_status_r_1__rd_addr__2_, dep_status_r_1__rd_addr__1_, dep_status_r_1__rd_addr__0_ };
  assign rd_match_vector[1] = issue_pkt_i[185:181] == { dep_status_r_1__rd_addr__4_, dep_status_r_1__rd_addr__3_, dep_status_r_1__rd_addr__2_, dep_status_r_1__rd_addr__1_, dep_status_r_1__rd_addr__0_ };
  assign rs1_match_vector[2] = issue_pkt_i[193:189] == { dep_status_r_2__rd_addr__4_, dep_status_r_2__rd_addr__3_, dep_status_r_2__rd_addr__2_, dep_status_r_2__rd_addr__1_, dep_status_r_2__rd_addr__0_ };
  assign rs2_match_vector[2] = issue_pkt_i[198:194] == { dep_status_r_2__rd_addr__4_, dep_status_r_2__rd_addr__3_, dep_status_r_2__rd_addr__2_, dep_status_r_2__rd_addr__1_, dep_status_r_2__rd_addr__0_ };
  assign rs3_match_vector[2] = issue_pkt_i[205:201] == { dep_status_r_2__rd_addr__4_, dep_status_r_2__rd_addr__3_, dep_status_r_2__rd_addr__2_, dep_status_r_2__rd_addr__1_, dep_status_r_2__rd_addr__0_ };
  assign rd_match_vector[2] = issue_pkt_i[185:181] == { dep_status_r_2__rd_addr__4_, dep_status_r_2__rd_addr__3_, dep_status_r_2__rd_addr__2_, dep_status_r_2__rd_addr__1_, dep_status_r_2__rd_addr__0_ };
  assign { N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2 } = (N0)? { dep_status_n_fflags_v_, dep_status_n_aux_iwb_v_, dep_status_n_aux_fwb_v_, dep_status_n_fint_iwb_v_, dep_status_n_fint_fwb_v_, dep_status_n_emem_iwb_v_, dep_status_n_emem_fwb_v_, dep_status_n_fmem_iwb_v_, dep_status_n_fmem_fwb_v_, dep_status_n_mul_iwb_v_, dep_status_n_fma_fwb_v_, dep_status_n_long_iwb_v_, dep_status_n_long_fwb_v_, dispatch_pkt_i[302:298] } : 
                                                                                                (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = dispatch_pkt_i[365];
  assign irs1_ispec_v = N21 & N23;
  assign N21 = N20 & issue_pkt_i[168];
  assign N20 = issue_pkt_i[160] & rs1_match_vector[0];
  assign N23 = N22 | dep_status_r_0__fint_iwb_v_;
  assign N22 = dep_status_r_0__aux_iwb_v_ | dep_status_r_0__emem_iwb_v_;
  assign irs2_ispec_v = N25 & N27;
  assign N25 = N24 & issue_pkt_i[168];
  assign N24 = issue_pkt_i[159] & rs2_match_vector[0];
  assign N27 = N26 | dep_status_r_0__fint_iwb_v_;
  assign N26 = dep_status_r_0__aux_iwb_v_ | dep_status_r_0__emem_iwb_v_;
  assign irs2_store_v = N29 & N31;
  assign N29 = N28 & issue_pkt_i[148];
  assign N28 = issue_pkt_i[159] & rs2_match_vector[0];
  assign N31 = N30 | dep_status_r_0__fint_iwb_v_;
  assign N30 = dep_status_r_0__aux_iwb_v_ | dep_status_r_0__emem_iwb_v_;
  assign ispec_v_o = irs1_ispec_v | irs2_ispec_v;
  assign clear_int_v_li = late_wb_pkt_i[78] & late_wb_yumi_i;
  assign clear_fp_v_li = late_wb_pkt_i[77] & late_wb_yumi_i;
  assign irs1_sb_raw_haz_v = issue_pkt_i[160] & irs_match_lo[0];
  assign irs2_sb_raw_haz_v = issue_pkt_i[159] & irs_match_lo[1];
  assign ird_sb_waw_haz_v = issue_pkt_i[155] & ird_match_lo;
  assign frs1_sb_raw_haz_v = issue_pkt_i[158] & frs_match_lo[0];
  assign frs2_sb_raw_haz_v = issue_pkt_i[157] & frs_match_lo[1];
  assign frs3_sb_raw_haz_v = issue_pkt_i[156] & frs_match_lo[2];
  assign frd_sb_waw_haz_v = issue_pkt_i[154] & frd_match_lo;
  assign iscore_haz_v = N36 | N38;
  assign N36 = N33 | N35;
  assign N33 = N32 & rd_match_vector[0];
  assign N32 = issue_pkt_i[155] & dep_status_r_0__long_iwb_v_;
  assign N35 = N34 & rd_match_vector[1];
  assign N34 = issue_pkt_i[155] & dep_status_r_1__long_iwb_v_;
  assign N38 = N37 & rd_match_vector[2];
  assign N37 = issue_pkt_i[155] & dep_status_r_2__long_iwb_v_;
  assign fscore_haz_v = N43 | N45;
  assign N43 = N40 | N42;
  assign N40 = N39 & rd_match_vector[0];
  assign N39 = issue_pkt_i[154] & dep_status_r_0__long_fwb_v_;
  assign N42 = N41 & rd_match_vector[1];
  assign N41 = issue_pkt_i[154] & dep_status_r_1__long_fwb_v_;
  assign N45 = N44 & rd_match_vector[2];
  assign N44 = issue_pkt_i[154] & dep_status_r_2__long_fwb_v_;
  assign irs1_data_haz_v[0] = N52 & N53;
  assign N52 = N46 & N51;
  assign N46 = issue_pkt_i[160] & rs1_match_vector[0];
  assign N51 = N50 | dep_status_r_0__long_iwb_v_;
  assign N50 = N49 | dep_status_r_0__fmem_iwb_v_;
  assign N49 = N48 | dep_status_r_0__emem_iwb_v_;
  assign N48 = N47 | dep_status_r_0__mul_iwb_v_;
  assign N47 = dep_status_r_0__fint_iwb_v_ | dep_status_r_0__aux_iwb_v_;
  assign N53 = ~irs1_ispec_v;
  assign irs2_data_haz_v[0] = N62 & N63;
  assign N62 = N60 & N61;
  assign N60 = N54 & N59;
  assign N54 = issue_pkt_i[159] & rs2_match_vector[0];
  assign N59 = N58 | dep_status_r_0__long_iwb_v_;
  assign N58 = N57 | dep_status_r_0__fmem_iwb_v_;
  assign N57 = N56 | dep_status_r_0__emem_iwb_v_;
  assign N56 = N55 | dep_status_r_0__mul_iwb_v_;
  assign N55 = dep_status_r_0__fint_iwb_v_ | dep_status_r_0__aux_iwb_v_;
  assign N61 = ~irs2_ispec_v;
  assign N63 = ~irs2_store_v;
  assign frs1_data_haz_v[0] = N64 & N69;
  assign N64 = issue_pkt_i[158] & rs1_match_vector[0];
  assign N69 = N68 | dep_status_r_0__long_fwb_v_;
  assign N68 = N67 | dep_status_r_0__fma_fwb_v_;
  assign N67 = N66 | dep_status_r_0__fmem_fwb_v_;
  assign N66 = N65 | dep_status_r_0__emem_fwb_v_;
  assign N65 = dep_status_r_0__fint_fwb_v_ | dep_status_r_0__aux_fwb_v_;
  assign frs2_data_haz_v[0] = N70 & N75;
  assign N70 = issue_pkt_i[157] & rs2_match_vector[0];
  assign N75 = N74 | dep_status_r_0__long_fwb_v_;
  assign N74 = N73 | dep_status_r_0__fma_fwb_v_;
  assign N73 = N72 | dep_status_r_0__fmem_fwb_v_;
  assign N72 = N71 | dep_status_r_0__emem_fwb_v_;
  assign N71 = dep_status_r_0__fint_fwb_v_ | dep_status_r_0__aux_fwb_v_;
  assign frs3_data_haz_v[0] = N76 & N81;
  assign N76 = issue_pkt_i[156] & rs3_match_vector[0];
  assign N81 = N80 | dep_status_r_0__long_fwb_v_;
  assign N80 = N79 | dep_status_r_0__fma_fwb_v_;
  assign N79 = N78 | dep_status_r_0__fmem_fwb_v_;
  assign N78 = N77 | dep_status_r_0__emem_fwb_v_;
  assign N77 = dep_status_r_0__fint_fwb_v_ | dep_status_r_0__aux_fwb_v_;
  assign irs1_data_haz_v[1] = N82 & N84;
  assign N82 = issue_pkt_i[160] & rs1_match_vector[1];
  assign N84 = N83 | dep_status_r_1__long_iwb_v_;
  assign N83 = dep_status_r_1__fmem_iwb_v_ | dep_status_r_1__mul_iwb_v_;
  assign irs2_data_haz_v[1] = N85 & N87;
  assign N85 = issue_pkt_i[159] & rs2_match_vector[1];
  assign N87 = N86 | dep_status_r_1__long_iwb_v_;
  assign N86 = dep_status_r_1__fmem_iwb_v_ | dep_status_r_1__mul_iwb_v_;
  assign frs1_data_haz_v[1] = N88 & N90;
  assign N88 = issue_pkt_i[158] & rs1_match_vector[1];
  assign N90 = N89 | dep_status_r_1__long_fwb_v_;
  assign N89 = dep_status_r_1__fmem_fwb_v_ | dep_status_r_1__fma_fwb_v_;
  assign frs2_data_haz_v[1] = N91 & N93;
  assign N91 = issue_pkt_i[157] & rs2_match_vector[1];
  assign N93 = N92 | dep_status_r_1__long_fwb_v_;
  assign N92 = dep_status_r_1__fmem_fwb_v_ | dep_status_r_1__fma_fwb_v_;
  assign frs3_data_haz_v[1] = N94 & N96;
  assign N94 = issue_pkt_i[156] & rs3_match_vector[1];
  assign N96 = N95 | dep_status_r_1__long_fwb_v_;
  assign N95 = dep_status_r_1__fmem_fwb_v_ | dep_status_r_1__fma_fwb_v_;
  assign irs1_data_haz_v[2] = N97 & dep_status_r_2__long_iwb_v_;
  assign N97 = issue_pkt_i[160] & rs1_match_vector[2];
  assign irs2_data_haz_v[2] = N98 & dep_status_r_2__long_iwb_v_;
  assign N98 = issue_pkt_i[159] & rs2_match_vector[2];
  assign frs1_data_haz_v[2] = N99 & N100;
  assign N99 = issue_pkt_i[158] & rs1_match_vector[2];
  assign N100 = dep_status_r_2__fma_fwb_v_ | dep_status_r_2__long_fwb_v_;
  assign frs2_data_haz_v[2] = N101 & N102;
  assign N101 = issue_pkt_i[157] & rs2_match_vector[2];
  assign N102 = dep_status_r_2__fma_fwb_v_ | dep_status_r_2__long_fwb_v_;
  assign frs3_data_haz_v[2] = N103 & N104;
  assign N103 = issue_pkt_i[156] & rs3_match_vector[2];
  assign N104 = dep_status_r_2__fma_fwb_v_ | dep_status_r_2__long_fwb_v_;
  assign fence_haz_v = issue_pkt_i[150] & N105;
  assign N105 = ~mem_ordered_i;
  assign fflags_haz_v = N106 & N110;
  assign N106 = issue_pkt_i[144] | issue_pkt_i[145];
  assign N110 = N109 | fdiv_busy_i;
  assign N109 = N108 | dep_status_r_3__fflags_v_;
  assign N108 = N107 | dep_status_r_2__fflags_v_;
  assign N107 = dep_status_r_0__fflags_v_ | dep_status_r_1__fflags_v_;
  assign control_haz_v = fence_haz_v | fflags_haz_v;
  assign data_haz_v = N127 | N130;
  assign N127 = N124 | N126;
  assign N124 = N121 | N123;
  assign N121 = N118 | N120;
  assign N118 = N115 | N117;
  assign N115 = N112 | N114;
  assign N112 = N111 | irs1_data_haz_v[0];
  assign N111 = irs1_data_haz_v[2] | irs1_data_haz_v[1];
  assign N114 = N113 | irs2_data_haz_v[0];
  assign N113 = irs2_data_haz_v[2] | irs2_data_haz_v[1];
  assign N117 = N116 | frs1_data_haz_v[0];
  assign N116 = frs1_data_haz_v[2] | frs1_data_haz_v[1];
  assign N120 = N119 | frs2_data_haz_v[0];
  assign N119 = frs2_data_haz_v[2] | frs2_data_haz_v[1];
  assign N123 = N122 | frs3_data_haz_v[0];
  assign N122 = frs3_data_haz_v[2] | frs3_data_haz_v[1];
  assign N126 = N125 | ird_sb_waw_haz_v;
  assign N125 = irs1_sb_raw_haz_v | irs2_sb_raw_haz_v;
  assign N130 = N129 | frd_sb_waw_haz_v;
  assign N129 = N128 | frs3_sb_raw_haz_v;
  assign N128 = frs1_sb_raw_haz_v | frs2_sb_raw_haz_v;
  assign struct_haz_v = N138 | N139;
  assign N138 = N136 | N137;
  assign N136 = N134 | N135;
  assign N134 = N132 | N133;
  assign N132 = N131 | iscore_haz_v;
  assign N131 = cmd_full_i | fscore_haz_v;
  assign N133 = mem_busy_i & issue_pkt_i[167];
  assign N135 = mem_busy_i & issue_pkt_i[165];
  assign N137 = fdiv_busy_i & issue_pkt_i[161];
  assign N139 = idiv_busy_i & issue_pkt_i[161];
  assign hazard_v_o = N140 | data_haz_v;
  assign N140 = struct_haz_v | control_haz_v;
  assign ordered_v_o = N143 & mem_ordered_i;
  assign N143 = ~N142;
  assign N142 = N141 | idiv_busy_i;
  assign N141 = mem_busy_i | fdiv_busy_i;
  assign dep_status_n_fflags_v_ = N144 | dispatch_pkt_i[279];
  assign N144 = dispatch_pkt_i[362] | dispatch_pkt_i[283];
  assign dep_status_n_fint_iwb_v_ = N145 & ispec_v_o;
  assign N145 = dispatch_pkt_i[285] & dispatch_pkt_i[272];
  assign dep_status_n_fint_fwb_v_ = dispatch_pkt_i[285] & dispatch_pkt_i[271];
  assign dep_status_n_aux_iwb_v_ = dispatch_pkt_i[283] & dispatch_pkt_i[272];
  assign dep_status_n_aux_fwb_v_ = dispatch_pkt_i[283] & dispatch_pkt_i[271];
  assign dep_status_n_emem_iwb_v_ = dispatch_pkt_i[284] & dispatch_pkt_i[272];
  assign dep_status_n_emem_fwb_v_ = dispatch_pkt_i[284] & dispatch_pkt_i[271];
  assign dep_status_n_fmem_iwb_v_ = dispatch_pkt_i[282] & dispatch_pkt_i[272];
  assign dep_status_n_fmem_fwb_v_ = dispatch_pkt_i[282] & dispatch_pkt_i[271];
  assign dep_status_n_mul_iwb_v_ = dispatch_pkt_i[280] & dispatch_pkt_i[272];
  assign dep_status_n_fma_fwb_v_ = dispatch_pkt_i[279] & dispatch_pkt_i[271];
  assign dep_status_n_long_iwb_v_ = dispatch_pkt_i[278] & dispatch_pkt_i[272];
  assign dep_status_n_long_fwb_v_ = dispatch_pkt_i[278] & dispatch_pkt_i[271];
  assign N1 = ~dispatch_pkt_i[365];

  always @(posedge clk_i) begin
    if(1'b1) begin
      dep_status_r_3__fflags_v__sv2v_reg <= dep_status_r_2__fflags_v_;
      dep_status_r_2__fflags_v__sv2v_reg <= dep_status_r_1__fflags_v_;
      dep_status_r_2__fma_fwb_v__sv2v_reg <= dep_status_r_1__fma_fwb_v_;
      dep_status_r_2__long_iwb_v__sv2v_reg <= dep_status_r_1__long_iwb_v_;
      dep_status_r_2__long_fwb_v__sv2v_reg <= dep_status_r_1__long_fwb_v_;
      dep_status_r_2__rd_addr__4__sv2v_reg <= dep_status_r_1__rd_addr__4_;
      dep_status_r_2__rd_addr__3__sv2v_reg <= dep_status_r_1__rd_addr__3_;
      dep_status_r_2__rd_addr__2__sv2v_reg <= dep_status_r_1__rd_addr__2_;
      dep_status_r_2__rd_addr__1__sv2v_reg <= dep_status_r_1__rd_addr__1_;
      dep_status_r_2__rd_addr__0__sv2v_reg <= dep_status_r_1__rd_addr__0_;
      dep_status_r_1__fflags_v__sv2v_reg <= dep_status_r_0__fflags_v_;
      dep_status_r_1__fmem_iwb_v__sv2v_reg <= dep_status_r_0__fmem_iwb_v_;
      dep_status_r_1__fmem_fwb_v__sv2v_reg <= dep_status_r_0__fmem_fwb_v_;
      dep_status_r_1__mul_iwb_v__sv2v_reg <= dep_status_r_0__mul_iwb_v_;
      dep_status_r_1__fma_fwb_v__sv2v_reg <= dep_status_r_0__fma_fwb_v_;
      dep_status_r_1__long_iwb_v__sv2v_reg <= dep_status_r_0__long_iwb_v_;
      dep_status_r_1__long_fwb_v__sv2v_reg <= dep_status_r_0__long_fwb_v_;
      dep_status_r_1__rd_addr__4__sv2v_reg <= dep_status_r_0__rd_addr__4_;
      dep_status_r_1__rd_addr__3__sv2v_reg <= dep_status_r_0__rd_addr__3_;
      dep_status_r_1__rd_addr__2__sv2v_reg <= dep_status_r_0__rd_addr__2_;
      dep_status_r_1__rd_addr__1__sv2v_reg <= dep_status_r_0__rd_addr__1_;
      dep_status_r_1__rd_addr__0__sv2v_reg <= dep_status_r_0__rd_addr__0_;
      dep_status_r_0__fflags_v__sv2v_reg <= N19;
      dep_status_r_0__aux_iwb_v__sv2v_reg <= N18;
      dep_status_r_0__aux_fwb_v__sv2v_reg <= N17;
      dep_status_r_0__fint_iwb_v__sv2v_reg <= N16;
      dep_status_r_0__fint_fwb_v__sv2v_reg <= N15;
      dep_status_r_0__emem_iwb_v__sv2v_reg <= N14;
      dep_status_r_0__emem_fwb_v__sv2v_reg <= N13;
      dep_status_r_0__fmem_iwb_v__sv2v_reg <= N12;
      dep_status_r_0__fmem_fwb_v__sv2v_reg <= N11;
      dep_status_r_0__mul_iwb_v__sv2v_reg <= N10;
      dep_status_r_0__fma_fwb_v__sv2v_reg <= N9;
      dep_status_r_0__long_iwb_v__sv2v_reg <= N8;
      dep_status_r_0__long_fwb_v__sv2v_reg <= N7;
      dep_status_r_0__rd_addr__4__sv2v_reg <= N6;
      dep_status_r_0__rd_addr__3__sv2v_reg <= N5;
      dep_status_r_0__rd_addr__2__sv2v_reg <= N4;
      dep_status_r_0__rd_addr__1__sv2v_reg <= N3;
      dep_status_r_0__rd_addr__0__sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_dff_en_0000002d
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [44:0] data_i;
  output [44:0] data_o;
  input clk_i;
  input en_i;
  wire [44:0] data_o;
  reg data_o_44_sv2v_reg,data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,
  data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,
  data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,
  data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,
  data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,
  data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,
  data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,
  data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_0000001e
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [29:0] data_i;
  output [29:0] data_o;
  input clk_i;
  input en_i;
  wire [29:0] data_o;
  reg data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,
  data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,
  data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,
  data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,
  data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bp_be_ptw_00_64_3_8_9
(
  clk_i,
  reset_i,
  busy_o,
  commit_pkt_i,
  trans_info_i,
  ordered_i,
  v_o,
  walk_o,
  itlb_fill_o,
  dtlb_fill_o,
  instr_page_fault_o,
  load_page_fault_o,
  store_page_fault_o,
  count_o,
  addr_o,
  pte_o,
  v_i,
  data_i
);

  input [213:0] commit_pkt_i;
  input [32:0] trans_info_i;
  output [2:0] count_o;
  output [63:0] addr_o;
  output [63:0] pte_o;
  input [63:0] data_i;
  input clk_i;
  input reset_i;
  input ordered_i;
  input v_i;
  output busy_o;
  output v_o;
  output walk_o;
  output itlb_fill_o;
  output dtlb_fill_o;
  output instr_page_fault_o;
  output load_page_fault_o;
  output store_page_fault_o;
  wire [2:0] count_o,count_r;
  wire [63:0] addr_o,pte_o;
  wire busy_o,v_o,walk_o,itlb_fill_o,dtlb_fill_o,instr_page_fault_o,load_page_fault_o,
  store_page_fault_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,
  N18,N19,N20,pte_o_35_,pte_o_5_,pte_o_4_,pte_o_3_,pte_o_2_,pte_o_1_,pte_o_0_,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,pte_is_leaf,pte_invalid,
  leaf_not_found,instr_r,s_priv_req,u_priv_req,priv_fault,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,misaligned_superpage,store_r,ad_fault,common_faults,
  instr_page_fault,load_r,load_page_fault,store_page_fault,page_fault_v,tlb_miss_v,
  walk_start,walk_ready,walk_next,walk_done,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,
  N58,walk_en,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,
  N76,N77,N79,N80,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,
  N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,
  N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,
  N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,
  N146,N147;
  wire [1:0] state_r,level_r,level_n,state_n;
  wire [11:0] vaddr_r;
  wire [26:0] vpn,partial_ppn;
  wire [11:3] walk_offset;
  wire [39:39] walk_addr;
  wire [27:0] ppn_n,ppn_r;
  reg state_r_1_sv2v_reg,state_r_0_sv2v_reg;
  assign state_r[1] = state_r_1_sv2v_reg;
  assign state_r[0] = state_r_0_sv2v_reg;
  assign pte_o[36] = 1'b0;
  assign pte_o[37] = 1'b0;
  assign pte_o[38] = 1'b0;
  assign pte_o[39] = 1'b0;
  assign pte_o[40] = 1'b0;
  assign pte_o[41] = 1'b0;
  assign pte_o[42] = 1'b0;
  assign pte_o[43] = 1'b0;
  assign pte_o[44] = 1'b0;
  assign pte_o[45] = 1'b0;
  assign pte_o[46] = 1'b0;
  assign pte_o[47] = 1'b0;
  assign pte_o[48] = 1'b0;
  assign pte_o[49] = 1'b0;
  assign pte_o[50] = 1'b0;
  assign pte_o[51] = 1'b0;
  assign pte_o[52] = 1'b0;
  assign pte_o[53] = 1'b0;
  assign pte_o[54] = 1'b0;
  assign pte_o[55] = 1'b0;
  assign pte_o[56] = 1'b0;
  assign pte_o[57] = 1'b0;
  assign pte_o[58] = 1'b0;
  assign pte_o[59] = 1'b0;
  assign pte_o[60] = 1'b0;
  assign pte_o[61] = 1'b0;
  assign pte_o[62] = 1'b0;
  assign pte_o[63] = 1'b0;
  assign addr_o[40] = 1'b0;
  assign addr_o[41] = 1'b0;
  assign addr_o[42] = 1'b0;
  assign addr_o[43] = 1'b0;
  assign addr_o[44] = 1'b0;
  assign addr_o[45] = 1'b0;
  assign addr_o[46] = 1'b0;
  assign addr_o[47] = 1'b0;
  assign addr_o[48] = 1'b0;
  assign addr_o[49] = 1'b0;
  assign addr_o[50] = 1'b0;
  assign addr_o[51] = 1'b0;
  assign addr_o[52] = 1'b0;
  assign addr_o[53] = 1'b0;
  assign addr_o[54] = 1'b0;
  assign addr_o[55] = 1'b0;
  assign addr_o[56] = 1'b0;
  assign addr_o[57] = 1'b0;
  assign addr_o[58] = 1'b0;
  assign addr_o[59] = 1'b0;
  assign addr_o[60] = 1'b0;
  assign addr_o[61] = 1'b0;
  assign addr_o[62] = 1'b0;
  assign addr_o[63] = 1'b0;
  assign pte_o_35_ = data_i[37];
  assign pte_o[35] = pte_o_35_;
  assign pte_o_5_ = data_i[6];
  assign pte_o[5] = pte_o_5_;
  assign pte_o_4_ = data_i[7];
  assign pte_o[4] = pte_o_4_;
  assign pte_o_3_ = data_i[4];
  assign pte_o[3] = pte_o_3_;
  assign pte_o_2_ = data_i[3];
  assign pte_o[2] = pte_o_2_;
  assign pte_o_1_ = data_i[2];
  assign pte_o[1] = pte_o_1_;
  assign pte_o_0_ = data_i[1];
  assign pte_o[0] = pte_o_0_;
  assign N21 = level_r > 1'b0;
  assign N23 = level_r > 1'b1;
  assign N25 = level_r > { 1'b1, 1'b0 };

  bsg_dff_en_0000002d
  miss_reg
  (
    .clk_i(clk_i),
    .data_i({ commit_pkt_i[9:9], commit_pkt_i[6:6], commit_pkt_i[7:7], commit_pkt_i[210:208], commit_pkt_i[127:89] }),
    .en_i(walk_start),
    .data_o({ instr_r, load_r, store_r, count_r, vpn, vaddr_r })
  );


  bsg_dff_en_0000001e
  walk_reg
  (
    .clk_i(clk_i),
    .data_i({ level_n, ppn_n }),
    .en_i(walk_en),
    .data_o({ level_r, ppn_r })
  );

  assign N62 = N82 & N85;
  assign N63 = state_r[1] | N85;
  assign N65 = N82 | state_r[0];
  assign N67 = state_r[1] & state_r[0];
  assign N76 = ~level_r[1];
  assign N77 = level_r[0] | N76;
  assign pte_o[7] = ~N77;
  assign N79 = ~level_r[0];
  assign N80 = N79 | level_r[1];
  assign pte_o[6] = ~N80;
  assign N82 = ~state_r[1];
  assign N83 = state_r[0] | N82;
  assign N84 = ~N83;
  assign N85 = ~state_r[0];
  assign N86 = N85 | state_r[1];
  assign N87 = ~N86;
  assign N88 = state_r[0] | state_r[1];
  assign N89 = ~N88;
  assign N90 = level_r[0] | level_r[1];
  assign N91 = ~N90;
  assign N92 = ~trans_info_i[31];
  assign N93 = N92 | trans_info_i[32];
  assign N94 = ~N93;
  assign N95 = trans_info_i[31] | trans_info_i[32];
  assign N96 = ~N95;
  assign { N58, N57 } = level_r - walk_next;
  assign N38 = level_r[0] & level_r[1];
  assign N37 = N0 & level_r[1];
  assign N0 = ~level_r[0];
  assign N36 = level_r[0] & N1;
  assign N1 = ~level_r[1];
  assign pte_o[16:8] = (N2)? vpn[8:0] : 
                       (N22)? partial_ppn[8:0] : 1'b0;
  assign N2 = N21;
  assign pte_o[25:17] = (N3)? vpn[17:9] : 
                        (N24)? partial_ppn[17:9] : 1'b0;
  assign N3 = N23;
  assign { N35, N34, N33, N32, N31, N30, N29, N28, N27 } = (N4)? vpn[26:18] : 
                                                           (N26)? partial_ppn[26:18] : 1'b0;
  assign N4 = N25;
  assign { N47, N46, N45, N44, N43, N42, N41, N40, N39 } = (N5)? data_i[36:28] : 
                                                           (N6)? data_i[27:19] : 
                                                           (N7)? data_i[18:10] : 1'b0;
  assign N5 = N38;
  assign N6 = N37;
  assign N7 = N36;
  assign ppn_n = (N8)? trans_info_i[30:3] : 
                 (N9)? { pte_o_35_, data_i[36:10] } : 1'b0;
  assign N8 = N54;
  assign N9 = N53;
  assign level_n = (N10)? { 1'b1, 1'b0 } : 
                   (N11)? { N58, N57 } : 1'b0;
  assign N10 = N56;
  assign N11 = N55;
  assign { walk_addr[39:39], partial_ppn } = (N12)? ppn_n : 
                                             (N13)? ppn_r : 1'b0;
  assign N12 = N60;
  assign N13 = N59;
  assign count_o = (N14)? count_r : 
                   (N15)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N14 = walk_done;
  assign N15 = N61;
  assign addr_o[39:0] = (N14)? { 1'b0, vpn, vaddr_r } : 
                        (N15)? { walk_addr[39:39], partial_ppn, walk_offset, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N73, N72 } = (N16)? { 1'b0, 1'b1 } : 
                        (N75)? { 1'b0, 1'b0 } : 
                        (N71)? { 1'b1, 1'b1 } : 1'b0;
  assign N16 = commit_pkt_i[4];
  assign state_n = (N17)? { 1'b0, N68 } : 
                   (N18)? { walk_ready, N69 } : 
                   (N19)? { 1'b1, N84 } : 
                   (N20)? { N73, N72 } : 1'b0;
  assign N17 = N62;
  assign N18 = N64;
  assign N19 = N66;
  assign N20 = N67;
  assign walk_offset[11] = (N50)? vpn[8] : 
                           (N52)? vpn[17] : 
                           (N51)? vpn[26] : 1'b0;
  assign walk_offset[10] = (N50)? vpn[7] : 
                           (N52)? vpn[16] : 
                           (N51)? vpn[25] : 1'b0;
  assign walk_offset[9] = (N50)? vpn[6] : 
                          (N52)? vpn[15] : 
                          (N51)? vpn[24] : 1'b0;
  assign walk_offset[8] = (N50)? vpn[5] : 
                          (N52)? vpn[14] : 
                          (N51)? vpn[23] : 1'b0;
  assign walk_offset[7] = (N50)? vpn[4] : 
                          (N52)? vpn[13] : 
                          (N51)? vpn[22] : 1'b0;
  assign walk_offset[6] = (N50)? vpn[3] : 
                          (N52)? vpn[12] : 
                          (N51)? vpn[21] : 1'b0;
  assign walk_offset[5] = (N50)? vpn[2] : 
                          (N52)? vpn[11] : 
                          (N51)? vpn[20] : 1'b0;
  assign walk_offset[4] = (N50)? vpn[1] : 
                          (N52)? vpn[10] : 
                          (N51)? vpn[19] : 1'b0;
  assign walk_offset[3] = (N50)? vpn[0] : 
                          (N52)? vpn[9] : 
                          (N51)? vpn[18] : 1'b0;
  assign N22 = ~N21;
  assign N24 = ~N23;
  assign N26 = ~N25;
  assign pte_o[34] = N35 | data_i[36];
  assign pte_o[33] = N34 | data_i[35];
  assign pte_o[32] = N33 | data_i[34];
  assign pte_o[31] = N32 | data_i[33];
  assign pte_o[30] = N31 | data_i[32];
  assign pte_o[29] = N30 | data_i[31];
  assign pte_o[28] = N29 | data_i[30];
  assign pte_o[27] = N28 | data_i[29];
  assign pte_o[26] = N27 | data_i[28];
  assign busy_o = ~N89;
  assign pte_is_leaf = N97 | pte_o_0_;
  assign N97 = pte_o_2_ | pte_o_1_;
  assign pte_invalid = N98 | N100;
  assign N98 = ~data_i[0];
  assign N100 = N99 & pte_o_1_;
  assign N99 = ~pte_o_0_;
  assign leaf_not_found = N91 & N101;
  assign N101 = ~pte_is_leaf;
  assign s_priv_req = N102 & N104;
  assign N102 = pte_is_leaf & N94;
  assign N104 = instr_r | N103;
  assign N103 = ~trans_info_i[1];
  assign u_priv_req = pte_is_leaf & N96;
  assign priv_fault = pte_is_leaf & N108;
  assign N108 = N105 | N107;
  assign N105 = pte_o_3_ & s_priv_req;
  assign N107 = N106 & u_priv_req;
  assign N106 = ~pte_o_3_;
  assign misaligned_superpage = N110 & N118;
  assign N110 = pte_is_leaf & N109;
  assign N109 = level_r[1] | level_r[0];
  assign N118 = N117 | N39;
  assign N117 = N116 | N40;
  assign N116 = N115 | N41;
  assign N115 = N114 | N42;
  assign N114 = N113 | N43;
  assign N113 = N112 | N44;
  assign N112 = N111 | N45;
  assign N111 = N47 | N46;
  assign ad_fault = pte_is_leaf & N122;
  assign N122 = N119 | N121;
  assign N119 = ~pte_o_5_;
  assign N121 = store_r & N120;
  assign N120 = ~pte_o_4_;
  assign common_faults = N125 | ad_fault;
  assign N125 = N124 | misaligned_superpage;
  assign N124 = N123 | priv_fault;
  assign N123 = pte_invalid | leaf_not_found;
  assign instr_page_fault = instr_r & N128;
  assign N128 = common_faults | N127;
  assign N127 = pte_is_leaf & N126;
  assign N126 = ~pte_o_2_;
  assign load_page_fault = load_r & N133;
  assign N133 = common_faults | N132;
  assign N132 = pte_is_leaf & N131;
  assign N131 = ~N130;
  assign N130 = pte_o_0_ | N129;
  assign N129 = pte_o_2_ & trans_info_i[0];
  assign store_page_fault = store_r & N136;
  assign N136 = common_faults | N135;
  assign N135 = pte_is_leaf & N134;
  assign N134 = ~pte_o_1_;
  assign page_fault_v = N137 | store_page_fault;
  assign N137 = instr_page_fault | load_page_fault;
  assign tlb_miss_v = N138 | commit_pkt_i[6];
  assign N138 = commit_pkt_i[9] | commit_pkt_i[7];
  assign walk_start = N89 & tlb_miss_v;
  assign walk_ready = N87 & ordered_i;
  assign walk_next = v_i & N140;
  assign N140 = ~N139;
  assign N139 = pte_is_leaf | page_fault_v;
  assign walk_done = v_i & N141;
  assign N141 = pte_is_leaf | page_fault_v;
  assign N48 = ~level_n[0];
  assign N49 = ~level_n[1];
  assign N50 = N48 & N49;
  assign N51 = N48 & level_n[1];
  assign N52 = level_n[0] & N49;
  assign N53 = ~walk_start;
  assign N54 = walk_start;
  assign N55 = ~walk_start;
  assign N56 = walk_start;
  assign walk_en = N142 | walk_done;
  assign N142 = walk_start | walk_next;
  assign N59 = ~walk_en;
  assign N60 = walk_en;
  assign v_o = N143 | walk_done;
  assign N143 = N84 | walk_next;
  assign walk_o = N84 | walk_next;
  assign itlb_fill_o = N144 & N145;
  assign N144 = walk_done & instr_r;
  assign N145 = ~page_fault_v;
  assign dtlb_fill_o = N147 & N145;
  assign N147 = walk_done & N146;
  assign N146 = ~instr_r;
  assign instr_page_fault_o = walk_done & instr_page_fault;
  assign load_page_fault_o = walk_done & load_page_fault;
  assign store_page_fault_o = walk_done & store_page_fault;
  assign N61 = ~walk_done;
  assign N64 = ~N63;
  assign N66 = ~N65;
  assign N68 = walk_start;
  assign N69 = ~walk_ready;
  assign N70 = walk_done | commit_pkt_i[4];
  assign N71 = ~N70;
  assign N74 = ~commit_pkt_i[4];
  assign N75 = walk_done & N74;

  always @(posedge clk_i) begin
    if(reset_i) begin
      state_r_1_sv2v_reg <= 1'b0;
      state_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      state_r_1_sv2v_reg <= state_n[1];
      state_r_0_sv2v_reg <= state_n[0];
    end 
  end


endmodule



module bsg_circular_ptr_slots_p128_max_add_p127
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [6:0] add_i;
  output [6:0] o;
  output [6:0] n_o;
  input clk;
  input reset_i;
  wire [6:0] o,n_o;
  reg o_6_sv2v_reg,o_5_sv2v_reg,o_4_sv2v_reg,o_3_sv2v_reg,o_2_sv2v_reg,o_1_sv2v_reg,
  o_0_sv2v_reg;
  assign o[6] = o_6_sv2v_reg;
  assign o[5] = o_5_sv2v_reg;
  assign o[4] = o_4_sv2v_reg;
  assign o[3] = o_3_sv2v_reg;
  assign o[2] = o_2_sv2v_reg;
  assign o[1] = o_1_sv2v_reg;
  assign o[0] = o_0_sv2v_reg;
  assign n_o = o + add_i;

  always @(posedge clk) begin
    if(reset_i) begin
      o_6_sv2v_reg <= 1'b0;
      o_5_sv2v_reg <= 1'b0;
      o_4_sv2v_reg <= 1'b0;
      o_3_sv2v_reg <= 1'b0;
      o_2_sv2v_reg <= 1'b0;
      o_1_sv2v_reg <= 1'b0;
      o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      o_6_sv2v_reg <= n_o[6];
      o_5_sv2v_reg <= n_o[5];
      o_4_sv2v_reg <= n_o[4];
      o_3_sv2v_reg <= n_o[3];
      o_2_sv2v_reg <= n_o[2];
      o_1_sv2v_reg <= n_o[1];
      o_0_sv2v_reg <= n_o[0];
    end 
  end


endmodule



module bsg_mem_1r1w_synth_00000050_00000008_0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [2:0] w_addr_i;
  input [79:0] w_data_i;
  input [2:0] r_addr_i;
  output [79:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [79:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45;
  wire [639:0] \nz.mem ;
  reg \nz.mem_639_sv2v_reg ,\nz.mem_638_sv2v_reg ,\nz.mem_637_sv2v_reg ,
  \nz.mem_636_sv2v_reg ,\nz.mem_635_sv2v_reg ,\nz.mem_634_sv2v_reg ,\nz.mem_633_sv2v_reg ,
  \nz.mem_632_sv2v_reg ,\nz.mem_631_sv2v_reg ,\nz.mem_630_sv2v_reg ,
  \nz.mem_629_sv2v_reg ,\nz.mem_628_sv2v_reg ,\nz.mem_627_sv2v_reg ,\nz.mem_626_sv2v_reg ,
  \nz.mem_625_sv2v_reg ,\nz.mem_624_sv2v_reg ,\nz.mem_623_sv2v_reg ,\nz.mem_622_sv2v_reg ,
  \nz.mem_621_sv2v_reg ,\nz.mem_620_sv2v_reg ,\nz.mem_619_sv2v_reg ,
  \nz.mem_618_sv2v_reg ,\nz.mem_617_sv2v_reg ,\nz.mem_616_sv2v_reg ,\nz.mem_615_sv2v_reg ,
  \nz.mem_614_sv2v_reg ,\nz.mem_613_sv2v_reg ,\nz.mem_612_sv2v_reg ,\nz.mem_611_sv2v_reg ,
  \nz.mem_610_sv2v_reg ,\nz.mem_609_sv2v_reg ,\nz.mem_608_sv2v_reg ,
  \nz.mem_607_sv2v_reg ,\nz.mem_606_sv2v_reg ,\nz.mem_605_sv2v_reg ,\nz.mem_604_sv2v_reg ,
  \nz.mem_603_sv2v_reg ,\nz.mem_602_sv2v_reg ,\nz.mem_601_sv2v_reg ,\nz.mem_600_sv2v_reg ,
  \nz.mem_599_sv2v_reg ,\nz.mem_598_sv2v_reg ,\nz.mem_597_sv2v_reg ,
  \nz.mem_596_sv2v_reg ,\nz.mem_595_sv2v_reg ,\nz.mem_594_sv2v_reg ,\nz.mem_593_sv2v_reg ,
  \nz.mem_592_sv2v_reg ,\nz.mem_591_sv2v_reg ,\nz.mem_590_sv2v_reg ,
  \nz.mem_589_sv2v_reg ,\nz.mem_588_sv2v_reg ,\nz.mem_587_sv2v_reg ,\nz.mem_586_sv2v_reg ,
  \nz.mem_585_sv2v_reg ,\nz.mem_584_sv2v_reg ,\nz.mem_583_sv2v_reg ,\nz.mem_582_sv2v_reg ,
  \nz.mem_581_sv2v_reg ,\nz.mem_580_sv2v_reg ,\nz.mem_579_sv2v_reg ,
  \nz.mem_578_sv2v_reg ,\nz.mem_577_sv2v_reg ,\nz.mem_576_sv2v_reg ,\nz.mem_575_sv2v_reg ,
  \nz.mem_574_sv2v_reg ,\nz.mem_573_sv2v_reg ,\nz.mem_572_sv2v_reg ,\nz.mem_571_sv2v_reg ,
  \nz.mem_570_sv2v_reg ,\nz.mem_569_sv2v_reg ,\nz.mem_568_sv2v_reg ,
  \nz.mem_567_sv2v_reg ,\nz.mem_566_sv2v_reg ,\nz.mem_565_sv2v_reg ,\nz.mem_564_sv2v_reg ,
  \nz.mem_563_sv2v_reg ,\nz.mem_562_sv2v_reg ,\nz.mem_561_sv2v_reg ,\nz.mem_560_sv2v_reg ,
  \nz.mem_559_sv2v_reg ,\nz.mem_558_sv2v_reg ,\nz.mem_557_sv2v_reg ,
  \nz.mem_556_sv2v_reg ,\nz.mem_555_sv2v_reg ,\nz.mem_554_sv2v_reg ,\nz.mem_553_sv2v_reg ,
  \nz.mem_552_sv2v_reg ,\nz.mem_551_sv2v_reg ,\nz.mem_550_sv2v_reg ,
  \nz.mem_549_sv2v_reg ,\nz.mem_548_sv2v_reg ,\nz.mem_547_sv2v_reg ,\nz.mem_546_sv2v_reg ,
  \nz.mem_545_sv2v_reg ,\nz.mem_544_sv2v_reg ,\nz.mem_543_sv2v_reg ,\nz.mem_542_sv2v_reg ,
  \nz.mem_541_sv2v_reg ,\nz.mem_540_sv2v_reg ,\nz.mem_539_sv2v_reg ,
  \nz.mem_538_sv2v_reg ,\nz.mem_537_sv2v_reg ,\nz.mem_536_sv2v_reg ,\nz.mem_535_sv2v_reg ,
  \nz.mem_534_sv2v_reg ,\nz.mem_533_sv2v_reg ,\nz.mem_532_sv2v_reg ,\nz.mem_531_sv2v_reg ,
  \nz.mem_530_sv2v_reg ,\nz.mem_529_sv2v_reg ,\nz.mem_528_sv2v_reg ,
  \nz.mem_527_sv2v_reg ,\nz.mem_526_sv2v_reg ,\nz.mem_525_sv2v_reg ,\nz.mem_524_sv2v_reg ,
  \nz.mem_523_sv2v_reg ,\nz.mem_522_sv2v_reg ,\nz.mem_521_sv2v_reg ,\nz.mem_520_sv2v_reg ,
  \nz.mem_519_sv2v_reg ,\nz.mem_518_sv2v_reg ,\nz.mem_517_sv2v_reg ,
  \nz.mem_516_sv2v_reg ,\nz.mem_515_sv2v_reg ,\nz.mem_514_sv2v_reg ,\nz.mem_513_sv2v_reg ,
  \nz.mem_512_sv2v_reg ,\nz.mem_511_sv2v_reg ,\nz.mem_510_sv2v_reg ,
  \nz.mem_509_sv2v_reg ,\nz.mem_508_sv2v_reg ,\nz.mem_507_sv2v_reg ,\nz.mem_506_sv2v_reg ,
  \nz.mem_505_sv2v_reg ,\nz.mem_504_sv2v_reg ,\nz.mem_503_sv2v_reg ,\nz.mem_502_sv2v_reg ,
  \nz.mem_501_sv2v_reg ,\nz.mem_500_sv2v_reg ,\nz.mem_499_sv2v_reg ,
  \nz.mem_498_sv2v_reg ,\nz.mem_497_sv2v_reg ,\nz.mem_496_sv2v_reg ,\nz.mem_495_sv2v_reg ,
  \nz.mem_494_sv2v_reg ,\nz.mem_493_sv2v_reg ,\nz.mem_492_sv2v_reg ,\nz.mem_491_sv2v_reg ,
  \nz.mem_490_sv2v_reg ,\nz.mem_489_sv2v_reg ,\nz.mem_488_sv2v_reg ,
  \nz.mem_487_sv2v_reg ,\nz.mem_486_sv2v_reg ,\nz.mem_485_sv2v_reg ,\nz.mem_484_sv2v_reg ,
  \nz.mem_483_sv2v_reg ,\nz.mem_482_sv2v_reg ,\nz.mem_481_sv2v_reg ,\nz.mem_480_sv2v_reg ,
  \nz.mem_479_sv2v_reg ,\nz.mem_478_sv2v_reg ,\nz.mem_477_sv2v_reg ,
  \nz.mem_476_sv2v_reg ,\nz.mem_475_sv2v_reg ,\nz.mem_474_sv2v_reg ,\nz.mem_473_sv2v_reg ,
  \nz.mem_472_sv2v_reg ,\nz.mem_471_sv2v_reg ,\nz.mem_470_sv2v_reg ,
  \nz.mem_469_sv2v_reg ,\nz.mem_468_sv2v_reg ,\nz.mem_467_sv2v_reg ,\nz.mem_466_sv2v_reg ,
  \nz.mem_465_sv2v_reg ,\nz.mem_464_sv2v_reg ,\nz.mem_463_sv2v_reg ,\nz.mem_462_sv2v_reg ,
  \nz.mem_461_sv2v_reg ,\nz.mem_460_sv2v_reg ,\nz.mem_459_sv2v_reg ,
  \nz.mem_458_sv2v_reg ,\nz.mem_457_sv2v_reg ,\nz.mem_456_sv2v_reg ,\nz.mem_455_sv2v_reg ,
  \nz.mem_454_sv2v_reg ,\nz.mem_453_sv2v_reg ,\nz.mem_452_sv2v_reg ,\nz.mem_451_sv2v_reg ,
  \nz.mem_450_sv2v_reg ,\nz.mem_449_sv2v_reg ,\nz.mem_448_sv2v_reg ,
  \nz.mem_447_sv2v_reg ,\nz.mem_446_sv2v_reg ,\nz.mem_445_sv2v_reg ,\nz.mem_444_sv2v_reg ,
  \nz.mem_443_sv2v_reg ,\nz.mem_442_sv2v_reg ,\nz.mem_441_sv2v_reg ,\nz.mem_440_sv2v_reg ,
  \nz.mem_439_sv2v_reg ,\nz.mem_438_sv2v_reg ,\nz.mem_437_sv2v_reg ,
  \nz.mem_436_sv2v_reg ,\nz.mem_435_sv2v_reg ,\nz.mem_434_sv2v_reg ,\nz.mem_433_sv2v_reg ,
  \nz.mem_432_sv2v_reg ,\nz.mem_431_sv2v_reg ,\nz.mem_430_sv2v_reg ,
  \nz.mem_429_sv2v_reg ,\nz.mem_428_sv2v_reg ,\nz.mem_427_sv2v_reg ,\nz.mem_426_sv2v_reg ,
  \nz.mem_425_sv2v_reg ,\nz.mem_424_sv2v_reg ,\nz.mem_423_sv2v_reg ,\nz.mem_422_sv2v_reg ,
  \nz.mem_421_sv2v_reg ,\nz.mem_420_sv2v_reg ,\nz.mem_419_sv2v_reg ,
  \nz.mem_418_sv2v_reg ,\nz.mem_417_sv2v_reg ,\nz.mem_416_sv2v_reg ,\nz.mem_415_sv2v_reg ,
  \nz.mem_414_sv2v_reg ,\nz.mem_413_sv2v_reg ,\nz.mem_412_sv2v_reg ,\nz.mem_411_sv2v_reg ,
  \nz.mem_410_sv2v_reg ,\nz.mem_409_sv2v_reg ,\nz.mem_408_sv2v_reg ,
  \nz.mem_407_sv2v_reg ,\nz.mem_406_sv2v_reg ,\nz.mem_405_sv2v_reg ,\nz.mem_404_sv2v_reg ,
  \nz.mem_403_sv2v_reg ,\nz.mem_402_sv2v_reg ,\nz.mem_401_sv2v_reg ,\nz.mem_400_sv2v_reg ,
  \nz.mem_399_sv2v_reg ,\nz.mem_398_sv2v_reg ,\nz.mem_397_sv2v_reg ,
  \nz.mem_396_sv2v_reg ,\nz.mem_395_sv2v_reg ,\nz.mem_394_sv2v_reg ,\nz.mem_393_sv2v_reg ,
  \nz.mem_392_sv2v_reg ,\nz.mem_391_sv2v_reg ,\nz.mem_390_sv2v_reg ,
  \nz.mem_389_sv2v_reg ,\nz.mem_388_sv2v_reg ,\nz.mem_387_sv2v_reg ,\nz.mem_386_sv2v_reg ,
  \nz.mem_385_sv2v_reg ,\nz.mem_384_sv2v_reg ,\nz.mem_383_sv2v_reg ,\nz.mem_382_sv2v_reg ,
  \nz.mem_381_sv2v_reg ,\nz.mem_380_sv2v_reg ,\nz.mem_379_sv2v_reg ,
  \nz.mem_378_sv2v_reg ,\nz.mem_377_sv2v_reg ,\nz.mem_376_sv2v_reg ,\nz.mem_375_sv2v_reg ,
  \nz.mem_374_sv2v_reg ,\nz.mem_373_sv2v_reg ,\nz.mem_372_sv2v_reg ,\nz.mem_371_sv2v_reg ,
  \nz.mem_370_sv2v_reg ,\nz.mem_369_sv2v_reg ,\nz.mem_368_sv2v_reg ,
  \nz.mem_367_sv2v_reg ,\nz.mem_366_sv2v_reg ,\nz.mem_365_sv2v_reg ,\nz.mem_364_sv2v_reg ,
  \nz.mem_363_sv2v_reg ,\nz.mem_362_sv2v_reg ,\nz.mem_361_sv2v_reg ,\nz.mem_360_sv2v_reg ,
  \nz.mem_359_sv2v_reg ,\nz.mem_358_sv2v_reg ,\nz.mem_357_sv2v_reg ,
  \nz.mem_356_sv2v_reg ,\nz.mem_355_sv2v_reg ,\nz.mem_354_sv2v_reg ,\nz.mem_353_sv2v_reg ,
  \nz.mem_352_sv2v_reg ,\nz.mem_351_sv2v_reg ,\nz.mem_350_sv2v_reg ,
  \nz.mem_349_sv2v_reg ,\nz.mem_348_sv2v_reg ,\nz.mem_347_sv2v_reg ,\nz.mem_346_sv2v_reg ,
  \nz.mem_345_sv2v_reg ,\nz.mem_344_sv2v_reg ,\nz.mem_343_sv2v_reg ,\nz.mem_342_sv2v_reg ,
  \nz.mem_341_sv2v_reg ,\nz.mem_340_sv2v_reg ,\nz.mem_339_sv2v_reg ,
  \nz.mem_338_sv2v_reg ,\nz.mem_337_sv2v_reg ,\nz.mem_336_sv2v_reg ,\nz.mem_335_sv2v_reg ,
  \nz.mem_334_sv2v_reg ,\nz.mem_333_sv2v_reg ,\nz.mem_332_sv2v_reg ,\nz.mem_331_sv2v_reg ,
  \nz.mem_330_sv2v_reg ,\nz.mem_329_sv2v_reg ,\nz.mem_328_sv2v_reg ,
  \nz.mem_327_sv2v_reg ,\nz.mem_326_sv2v_reg ,\nz.mem_325_sv2v_reg ,\nz.mem_324_sv2v_reg ,
  \nz.mem_323_sv2v_reg ,\nz.mem_322_sv2v_reg ,\nz.mem_321_sv2v_reg ,\nz.mem_320_sv2v_reg ,
  \nz.mem_319_sv2v_reg ,\nz.mem_318_sv2v_reg ,\nz.mem_317_sv2v_reg ,
  \nz.mem_316_sv2v_reg ,\nz.mem_315_sv2v_reg ,\nz.mem_314_sv2v_reg ,\nz.mem_313_sv2v_reg ,
  \nz.mem_312_sv2v_reg ,\nz.mem_311_sv2v_reg ,\nz.mem_310_sv2v_reg ,
  \nz.mem_309_sv2v_reg ,\nz.mem_308_sv2v_reg ,\nz.mem_307_sv2v_reg ,\nz.mem_306_sv2v_reg ,
  \nz.mem_305_sv2v_reg ,\nz.mem_304_sv2v_reg ,\nz.mem_303_sv2v_reg ,\nz.mem_302_sv2v_reg ,
  \nz.mem_301_sv2v_reg ,\nz.mem_300_sv2v_reg ,\nz.mem_299_sv2v_reg ,
  \nz.mem_298_sv2v_reg ,\nz.mem_297_sv2v_reg ,\nz.mem_296_sv2v_reg ,\nz.mem_295_sv2v_reg ,
  \nz.mem_294_sv2v_reg ,\nz.mem_293_sv2v_reg ,\nz.mem_292_sv2v_reg ,\nz.mem_291_sv2v_reg ,
  \nz.mem_290_sv2v_reg ,\nz.mem_289_sv2v_reg ,\nz.mem_288_sv2v_reg ,
  \nz.mem_287_sv2v_reg ,\nz.mem_286_sv2v_reg ,\nz.mem_285_sv2v_reg ,\nz.mem_284_sv2v_reg ,
  \nz.mem_283_sv2v_reg ,\nz.mem_282_sv2v_reg ,\nz.mem_281_sv2v_reg ,\nz.mem_280_sv2v_reg ,
  \nz.mem_279_sv2v_reg ,\nz.mem_278_sv2v_reg ,\nz.mem_277_sv2v_reg ,
  \nz.mem_276_sv2v_reg ,\nz.mem_275_sv2v_reg ,\nz.mem_274_sv2v_reg ,\nz.mem_273_sv2v_reg ,
  \nz.mem_272_sv2v_reg ,\nz.mem_271_sv2v_reg ,\nz.mem_270_sv2v_reg ,
  \nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,\nz.mem_267_sv2v_reg ,\nz.mem_266_sv2v_reg ,
  \nz.mem_265_sv2v_reg ,\nz.mem_264_sv2v_reg ,\nz.mem_263_sv2v_reg ,\nz.mem_262_sv2v_reg ,
  \nz.mem_261_sv2v_reg ,\nz.mem_260_sv2v_reg ,\nz.mem_259_sv2v_reg ,
  \nz.mem_258_sv2v_reg ,\nz.mem_257_sv2v_reg ,\nz.mem_256_sv2v_reg ,\nz.mem_255_sv2v_reg ,
  \nz.mem_254_sv2v_reg ,\nz.mem_253_sv2v_reg ,\nz.mem_252_sv2v_reg ,\nz.mem_251_sv2v_reg ,
  \nz.mem_250_sv2v_reg ,\nz.mem_249_sv2v_reg ,\nz.mem_248_sv2v_reg ,
  \nz.mem_247_sv2v_reg ,\nz.mem_246_sv2v_reg ,\nz.mem_245_sv2v_reg ,\nz.mem_244_sv2v_reg ,
  \nz.mem_243_sv2v_reg ,\nz.mem_242_sv2v_reg ,\nz.mem_241_sv2v_reg ,\nz.mem_240_sv2v_reg ,
  \nz.mem_239_sv2v_reg ,\nz.mem_238_sv2v_reg ,\nz.mem_237_sv2v_reg ,
  \nz.mem_236_sv2v_reg ,\nz.mem_235_sv2v_reg ,\nz.mem_234_sv2v_reg ,\nz.mem_233_sv2v_reg ,
  \nz.mem_232_sv2v_reg ,\nz.mem_231_sv2v_reg ,\nz.mem_230_sv2v_reg ,
  \nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,\nz.mem_227_sv2v_reg ,\nz.mem_226_sv2v_reg ,
  \nz.mem_225_sv2v_reg ,\nz.mem_224_sv2v_reg ,\nz.mem_223_sv2v_reg ,\nz.mem_222_sv2v_reg ,
  \nz.mem_221_sv2v_reg ,\nz.mem_220_sv2v_reg ,\nz.mem_219_sv2v_reg ,
  \nz.mem_218_sv2v_reg ,\nz.mem_217_sv2v_reg ,\nz.mem_216_sv2v_reg ,\nz.mem_215_sv2v_reg ,
  \nz.mem_214_sv2v_reg ,\nz.mem_213_sv2v_reg ,\nz.mem_212_sv2v_reg ,\nz.mem_211_sv2v_reg ,
  \nz.mem_210_sv2v_reg ,\nz.mem_209_sv2v_reg ,\nz.mem_208_sv2v_reg ,
  \nz.mem_207_sv2v_reg ,\nz.mem_206_sv2v_reg ,\nz.mem_205_sv2v_reg ,\nz.mem_204_sv2v_reg ,
  \nz.mem_203_sv2v_reg ,\nz.mem_202_sv2v_reg ,\nz.mem_201_sv2v_reg ,\nz.mem_200_sv2v_reg ,
  \nz.mem_199_sv2v_reg ,\nz.mem_198_sv2v_reg ,\nz.mem_197_sv2v_reg ,
  \nz.mem_196_sv2v_reg ,\nz.mem_195_sv2v_reg ,\nz.mem_194_sv2v_reg ,\nz.mem_193_sv2v_reg ,
  \nz.mem_192_sv2v_reg ,\nz.mem_191_sv2v_reg ,\nz.mem_190_sv2v_reg ,
  \nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,\nz.mem_187_sv2v_reg ,\nz.mem_186_sv2v_reg ,
  \nz.mem_185_sv2v_reg ,\nz.mem_184_sv2v_reg ,\nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,
  \nz.mem_181_sv2v_reg ,\nz.mem_180_sv2v_reg ,\nz.mem_179_sv2v_reg ,
  \nz.mem_178_sv2v_reg ,\nz.mem_177_sv2v_reg ,\nz.mem_176_sv2v_reg ,\nz.mem_175_sv2v_reg ,
  \nz.mem_174_sv2v_reg ,\nz.mem_173_sv2v_reg ,\nz.mem_172_sv2v_reg ,\nz.mem_171_sv2v_reg ,
  \nz.mem_170_sv2v_reg ,\nz.mem_169_sv2v_reg ,\nz.mem_168_sv2v_reg ,
  \nz.mem_167_sv2v_reg ,\nz.mem_166_sv2v_reg ,\nz.mem_165_sv2v_reg ,\nz.mem_164_sv2v_reg ,
  \nz.mem_163_sv2v_reg ,\nz.mem_162_sv2v_reg ,\nz.mem_161_sv2v_reg ,\nz.mem_160_sv2v_reg ,
  \nz.mem_159_sv2v_reg ,\nz.mem_158_sv2v_reg ,\nz.mem_157_sv2v_reg ,
  \nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,\nz.mem_154_sv2v_reg ,\nz.mem_153_sv2v_reg ,
  \nz.mem_152_sv2v_reg ,\nz.mem_151_sv2v_reg ,\nz.mem_150_sv2v_reg ,
  \nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,\nz.mem_147_sv2v_reg ,\nz.mem_146_sv2v_reg ,
  \nz.mem_145_sv2v_reg ,\nz.mem_144_sv2v_reg ,\nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,
  \nz.mem_141_sv2v_reg ,\nz.mem_140_sv2v_reg ,\nz.mem_139_sv2v_reg ,
  \nz.mem_138_sv2v_reg ,\nz.mem_137_sv2v_reg ,\nz.mem_136_sv2v_reg ,\nz.mem_135_sv2v_reg ,
  \nz.mem_134_sv2v_reg ,\nz.mem_133_sv2v_reg ,\nz.mem_132_sv2v_reg ,\nz.mem_131_sv2v_reg ,
  \nz.mem_130_sv2v_reg ,\nz.mem_129_sv2v_reg ,\nz.mem_128_sv2v_reg ,
  \nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,\nz.mem_125_sv2v_reg ,\nz.mem_124_sv2v_reg ,
  \nz.mem_123_sv2v_reg ,\nz.mem_122_sv2v_reg ,\nz.mem_121_sv2v_reg ,\nz.mem_120_sv2v_reg ,
  \nz.mem_119_sv2v_reg ,\nz.mem_118_sv2v_reg ,\nz.mem_117_sv2v_reg ,
  \nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,\nz.mem_114_sv2v_reg ,\nz.mem_113_sv2v_reg ,
  \nz.mem_112_sv2v_reg ,\nz.mem_111_sv2v_reg ,\nz.mem_110_sv2v_reg ,
  \nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,\nz.mem_107_sv2v_reg ,\nz.mem_106_sv2v_reg ,
  \nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,\nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,
  \nz.mem_101_sv2v_reg ,\nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,
  \nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,\nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,
  \nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,\nz.mem_92_sv2v_reg ,\nz.mem_91_sv2v_reg ,
  \nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,\nz.mem_88_sv2v_reg ,\nz.mem_87_sv2v_reg ,
  \nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,\nz.mem_83_sv2v_reg ,
  \nz.mem_82_sv2v_reg ,\nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,
  \nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,\nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,
  \nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,\nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,
  \nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,\nz.mem_69_sv2v_reg ,\nz.mem_68_sv2v_reg ,
  \nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,
  \nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,\nz.mem_60_sv2v_reg ,
  \nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,
  \nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,
  \nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,
  \nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,
  \nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,\nz.mem_41_sv2v_reg ,
  \nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,
  \nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,
  \nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,
  \nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,
  \nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,\nz.mem_22_sv2v_reg ,
  \nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,
  \nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,
  \nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,
  \nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,
  \nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,
  \nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.mem [639] = \nz.mem_639_sv2v_reg ;
  assign \nz.mem [638] = \nz.mem_638_sv2v_reg ;
  assign \nz.mem [637] = \nz.mem_637_sv2v_reg ;
  assign \nz.mem [636] = \nz.mem_636_sv2v_reg ;
  assign \nz.mem [635] = \nz.mem_635_sv2v_reg ;
  assign \nz.mem [634] = \nz.mem_634_sv2v_reg ;
  assign \nz.mem [633] = \nz.mem_633_sv2v_reg ;
  assign \nz.mem [632] = \nz.mem_632_sv2v_reg ;
  assign \nz.mem [631] = \nz.mem_631_sv2v_reg ;
  assign \nz.mem [630] = \nz.mem_630_sv2v_reg ;
  assign \nz.mem [629] = \nz.mem_629_sv2v_reg ;
  assign \nz.mem [628] = \nz.mem_628_sv2v_reg ;
  assign \nz.mem [627] = \nz.mem_627_sv2v_reg ;
  assign \nz.mem [626] = \nz.mem_626_sv2v_reg ;
  assign \nz.mem [625] = \nz.mem_625_sv2v_reg ;
  assign \nz.mem [624] = \nz.mem_624_sv2v_reg ;
  assign \nz.mem [623] = \nz.mem_623_sv2v_reg ;
  assign \nz.mem [622] = \nz.mem_622_sv2v_reg ;
  assign \nz.mem [621] = \nz.mem_621_sv2v_reg ;
  assign \nz.mem [620] = \nz.mem_620_sv2v_reg ;
  assign \nz.mem [619] = \nz.mem_619_sv2v_reg ;
  assign \nz.mem [618] = \nz.mem_618_sv2v_reg ;
  assign \nz.mem [617] = \nz.mem_617_sv2v_reg ;
  assign \nz.mem [616] = \nz.mem_616_sv2v_reg ;
  assign \nz.mem [615] = \nz.mem_615_sv2v_reg ;
  assign \nz.mem [614] = \nz.mem_614_sv2v_reg ;
  assign \nz.mem [613] = \nz.mem_613_sv2v_reg ;
  assign \nz.mem [612] = \nz.mem_612_sv2v_reg ;
  assign \nz.mem [611] = \nz.mem_611_sv2v_reg ;
  assign \nz.mem [610] = \nz.mem_610_sv2v_reg ;
  assign \nz.mem [609] = \nz.mem_609_sv2v_reg ;
  assign \nz.mem [608] = \nz.mem_608_sv2v_reg ;
  assign \nz.mem [607] = \nz.mem_607_sv2v_reg ;
  assign \nz.mem [606] = \nz.mem_606_sv2v_reg ;
  assign \nz.mem [605] = \nz.mem_605_sv2v_reg ;
  assign \nz.mem [604] = \nz.mem_604_sv2v_reg ;
  assign \nz.mem [603] = \nz.mem_603_sv2v_reg ;
  assign \nz.mem [602] = \nz.mem_602_sv2v_reg ;
  assign \nz.mem [601] = \nz.mem_601_sv2v_reg ;
  assign \nz.mem [600] = \nz.mem_600_sv2v_reg ;
  assign \nz.mem [599] = \nz.mem_599_sv2v_reg ;
  assign \nz.mem [598] = \nz.mem_598_sv2v_reg ;
  assign \nz.mem [597] = \nz.mem_597_sv2v_reg ;
  assign \nz.mem [596] = \nz.mem_596_sv2v_reg ;
  assign \nz.mem [595] = \nz.mem_595_sv2v_reg ;
  assign \nz.mem [594] = \nz.mem_594_sv2v_reg ;
  assign \nz.mem [593] = \nz.mem_593_sv2v_reg ;
  assign \nz.mem [592] = \nz.mem_592_sv2v_reg ;
  assign \nz.mem [591] = \nz.mem_591_sv2v_reg ;
  assign \nz.mem [590] = \nz.mem_590_sv2v_reg ;
  assign \nz.mem [589] = \nz.mem_589_sv2v_reg ;
  assign \nz.mem [588] = \nz.mem_588_sv2v_reg ;
  assign \nz.mem [587] = \nz.mem_587_sv2v_reg ;
  assign \nz.mem [586] = \nz.mem_586_sv2v_reg ;
  assign \nz.mem [585] = \nz.mem_585_sv2v_reg ;
  assign \nz.mem [584] = \nz.mem_584_sv2v_reg ;
  assign \nz.mem [583] = \nz.mem_583_sv2v_reg ;
  assign \nz.mem [582] = \nz.mem_582_sv2v_reg ;
  assign \nz.mem [581] = \nz.mem_581_sv2v_reg ;
  assign \nz.mem [580] = \nz.mem_580_sv2v_reg ;
  assign \nz.mem [579] = \nz.mem_579_sv2v_reg ;
  assign \nz.mem [578] = \nz.mem_578_sv2v_reg ;
  assign \nz.mem [577] = \nz.mem_577_sv2v_reg ;
  assign \nz.mem [576] = \nz.mem_576_sv2v_reg ;
  assign \nz.mem [575] = \nz.mem_575_sv2v_reg ;
  assign \nz.mem [574] = \nz.mem_574_sv2v_reg ;
  assign \nz.mem [573] = \nz.mem_573_sv2v_reg ;
  assign \nz.mem [572] = \nz.mem_572_sv2v_reg ;
  assign \nz.mem [571] = \nz.mem_571_sv2v_reg ;
  assign \nz.mem [570] = \nz.mem_570_sv2v_reg ;
  assign \nz.mem [569] = \nz.mem_569_sv2v_reg ;
  assign \nz.mem [568] = \nz.mem_568_sv2v_reg ;
  assign \nz.mem [567] = \nz.mem_567_sv2v_reg ;
  assign \nz.mem [566] = \nz.mem_566_sv2v_reg ;
  assign \nz.mem [565] = \nz.mem_565_sv2v_reg ;
  assign \nz.mem [564] = \nz.mem_564_sv2v_reg ;
  assign \nz.mem [563] = \nz.mem_563_sv2v_reg ;
  assign \nz.mem [562] = \nz.mem_562_sv2v_reg ;
  assign \nz.mem [561] = \nz.mem_561_sv2v_reg ;
  assign \nz.mem [560] = \nz.mem_560_sv2v_reg ;
  assign \nz.mem [559] = \nz.mem_559_sv2v_reg ;
  assign \nz.mem [558] = \nz.mem_558_sv2v_reg ;
  assign \nz.mem [557] = \nz.mem_557_sv2v_reg ;
  assign \nz.mem [556] = \nz.mem_556_sv2v_reg ;
  assign \nz.mem [555] = \nz.mem_555_sv2v_reg ;
  assign \nz.mem [554] = \nz.mem_554_sv2v_reg ;
  assign \nz.mem [553] = \nz.mem_553_sv2v_reg ;
  assign \nz.mem [552] = \nz.mem_552_sv2v_reg ;
  assign \nz.mem [551] = \nz.mem_551_sv2v_reg ;
  assign \nz.mem [550] = \nz.mem_550_sv2v_reg ;
  assign \nz.mem [549] = \nz.mem_549_sv2v_reg ;
  assign \nz.mem [548] = \nz.mem_548_sv2v_reg ;
  assign \nz.mem [547] = \nz.mem_547_sv2v_reg ;
  assign \nz.mem [546] = \nz.mem_546_sv2v_reg ;
  assign \nz.mem [545] = \nz.mem_545_sv2v_reg ;
  assign \nz.mem [544] = \nz.mem_544_sv2v_reg ;
  assign \nz.mem [543] = \nz.mem_543_sv2v_reg ;
  assign \nz.mem [542] = \nz.mem_542_sv2v_reg ;
  assign \nz.mem [541] = \nz.mem_541_sv2v_reg ;
  assign \nz.mem [540] = \nz.mem_540_sv2v_reg ;
  assign \nz.mem [539] = \nz.mem_539_sv2v_reg ;
  assign \nz.mem [538] = \nz.mem_538_sv2v_reg ;
  assign \nz.mem [537] = \nz.mem_537_sv2v_reg ;
  assign \nz.mem [536] = \nz.mem_536_sv2v_reg ;
  assign \nz.mem [535] = \nz.mem_535_sv2v_reg ;
  assign \nz.mem [534] = \nz.mem_534_sv2v_reg ;
  assign \nz.mem [533] = \nz.mem_533_sv2v_reg ;
  assign \nz.mem [532] = \nz.mem_532_sv2v_reg ;
  assign \nz.mem [531] = \nz.mem_531_sv2v_reg ;
  assign \nz.mem [530] = \nz.mem_530_sv2v_reg ;
  assign \nz.mem [529] = \nz.mem_529_sv2v_reg ;
  assign \nz.mem [528] = \nz.mem_528_sv2v_reg ;
  assign \nz.mem [527] = \nz.mem_527_sv2v_reg ;
  assign \nz.mem [526] = \nz.mem_526_sv2v_reg ;
  assign \nz.mem [525] = \nz.mem_525_sv2v_reg ;
  assign \nz.mem [524] = \nz.mem_524_sv2v_reg ;
  assign \nz.mem [523] = \nz.mem_523_sv2v_reg ;
  assign \nz.mem [522] = \nz.mem_522_sv2v_reg ;
  assign \nz.mem [521] = \nz.mem_521_sv2v_reg ;
  assign \nz.mem [520] = \nz.mem_520_sv2v_reg ;
  assign \nz.mem [519] = \nz.mem_519_sv2v_reg ;
  assign \nz.mem [518] = \nz.mem_518_sv2v_reg ;
  assign \nz.mem [517] = \nz.mem_517_sv2v_reg ;
  assign \nz.mem [516] = \nz.mem_516_sv2v_reg ;
  assign \nz.mem [515] = \nz.mem_515_sv2v_reg ;
  assign \nz.mem [514] = \nz.mem_514_sv2v_reg ;
  assign \nz.mem [513] = \nz.mem_513_sv2v_reg ;
  assign \nz.mem [512] = \nz.mem_512_sv2v_reg ;
  assign \nz.mem [511] = \nz.mem_511_sv2v_reg ;
  assign \nz.mem [510] = \nz.mem_510_sv2v_reg ;
  assign \nz.mem [509] = \nz.mem_509_sv2v_reg ;
  assign \nz.mem [508] = \nz.mem_508_sv2v_reg ;
  assign \nz.mem [507] = \nz.mem_507_sv2v_reg ;
  assign \nz.mem [506] = \nz.mem_506_sv2v_reg ;
  assign \nz.mem [505] = \nz.mem_505_sv2v_reg ;
  assign \nz.mem [504] = \nz.mem_504_sv2v_reg ;
  assign \nz.mem [503] = \nz.mem_503_sv2v_reg ;
  assign \nz.mem [502] = \nz.mem_502_sv2v_reg ;
  assign \nz.mem [501] = \nz.mem_501_sv2v_reg ;
  assign \nz.mem [500] = \nz.mem_500_sv2v_reg ;
  assign \nz.mem [499] = \nz.mem_499_sv2v_reg ;
  assign \nz.mem [498] = \nz.mem_498_sv2v_reg ;
  assign \nz.mem [497] = \nz.mem_497_sv2v_reg ;
  assign \nz.mem [496] = \nz.mem_496_sv2v_reg ;
  assign \nz.mem [495] = \nz.mem_495_sv2v_reg ;
  assign \nz.mem [494] = \nz.mem_494_sv2v_reg ;
  assign \nz.mem [493] = \nz.mem_493_sv2v_reg ;
  assign \nz.mem [492] = \nz.mem_492_sv2v_reg ;
  assign \nz.mem [491] = \nz.mem_491_sv2v_reg ;
  assign \nz.mem [490] = \nz.mem_490_sv2v_reg ;
  assign \nz.mem [489] = \nz.mem_489_sv2v_reg ;
  assign \nz.mem [488] = \nz.mem_488_sv2v_reg ;
  assign \nz.mem [487] = \nz.mem_487_sv2v_reg ;
  assign \nz.mem [486] = \nz.mem_486_sv2v_reg ;
  assign \nz.mem [485] = \nz.mem_485_sv2v_reg ;
  assign \nz.mem [484] = \nz.mem_484_sv2v_reg ;
  assign \nz.mem [483] = \nz.mem_483_sv2v_reg ;
  assign \nz.mem [482] = \nz.mem_482_sv2v_reg ;
  assign \nz.mem [481] = \nz.mem_481_sv2v_reg ;
  assign \nz.mem [480] = \nz.mem_480_sv2v_reg ;
  assign \nz.mem [479] = \nz.mem_479_sv2v_reg ;
  assign \nz.mem [478] = \nz.mem_478_sv2v_reg ;
  assign \nz.mem [477] = \nz.mem_477_sv2v_reg ;
  assign \nz.mem [476] = \nz.mem_476_sv2v_reg ;
  assign \nz.mem [475] = \nz.mem_475_sv2v_reg ;
  assign \nz.mem [474] = \nz.mem_474_sv2v_reg ;
  assign \nz.mem [473] = \nz.mem_473_sv2v_reg ;
  assign \nz.mem [472] = \nz.mem_472_sv2v_reg ;
  assign \nz.mem [471] = \nz.mem_471_sv2v_reg ;
  assign \nz.mem [470] = \nz.mem_470_sv2v_reg ;
  assign \nz.mem [469] = \nz.mem_469_sv2v_reg ;
  assign \nz.mem [468] = \nz.mem_468_sv2v_reg ;
  assign \nz.mem [467] = \nz.mem_467_sv2v_reg ;
  assign \nz.mem [466] = \nz.mem_466_sv2v_reg ;
  assign \nz.mem [465] = \nz.mem_465_sv2v_reg ;
  assign \nz.mem [464] = \nz.mem_464_sv2v_reg ;
  assign \nz.mem [463] = \nz.mem_463_sv2v_reg ;
  assign \nz.mem [462] = \nz.mem_462_sv2v_reg ;
  assign \nz.mem [461] = \nz.mem_461_sv2v_reg ;
  assign \nz.mem [460] = \nz.mem_460_sv2v_reg ;
  assign \nz.mem [459] = \nz.mem_459_sv2v_reg ;
  assign \nz.mem [458] = \nz.mem_458_sv2v_reg ;
  assign \nz.mem [457] = \nz.mem_457_sv2v_reg ;
  assign \nz.mem [456] = \nz.mem_456_sv2v_reg ;
  assign \nz.mem [455] = \nz.mem_455_sv2v_reg ;
  assign \nz.mem [454] = \nz.mem_454_sv2v_reg ;
  assign \nz.mem [453] = \nz.mem_453_sv2v_reg ;
  assign \nz.mem [452] = \nz.mem_452_sv2v_reg ;
  assign \nz.mem [451] = \nz.mem_451_sv2v_reg ;
  assign \nz.mem [450] = \nz.mem_450_sv2v_reg ;
  assign \nz.mem [449] = \nz.mem_449_sv2v_reg ;
  assign \nz.mem [448] = \nz.mem_448_sv2v_reg ;
  assign \nz.mem [447] = \nz.mem_447_sv2v_reg ;
  assign \nz.mem [446] = \nz.mem_446_sv2v_reg ;
  assign \nz.mem [445] = \nz.mem_445_sv2v_reg ;
  assign \nz.mem [444] = \nz.mem_444_sv2v_reg ;
  assign \nz.mem [443] = \nz.mem_443_sv2v_reg ;
  assign \nz.mem [442] = \nz.mem_442_sv2v_reg ;
  assign \nz.mem [441] = \nz.mem_441_sv2v_reg ;
  assign \nz.mem [440] = \nz.mem_440_sv2v_reg ;
  assign \nz.mem [439] = \nz.mem_439_sv2v_reg ;
  assign \nz.mem [438] = \nz.mem_438_sv2v_reg ;
  assign \nz.mem [437] = \nz.mem_437_sv2v_reg ;
  assign \nz.mem [436] = \nz.mem_436_sv2v_reg ;
  assign \nz.mem [435] = \nz.mem_435_sv2v_reg ;
  assign \nz.mem [434] = \nz.mem_434_sv2v_reg ;
  assign \nz.mem [433] = \nz.mem_433_sv2v_reg ;
  assign \nz.mem [432] = \nz.mem_432_sv2v_reg ;
  assign \nz.mem [431] = \nz.mem_431_sv2v_reg ;
  assign \nz.mem [430] = \nz.mem_430_sv2v_reg ;
  assign \nz.mem [429] = \nz.mem_429_sv2v_reg ;
  assign \nz.mem [428] = \nz.mem_428_sv2v_reg ;
  assign \nz.mem [427] = \nz.mem_427_sv2v_reg ;
  assign \nz.mem [426] = \nz.mem_426_sv2v_reg ;
  assign \nz.mem [425] = \nz.mem_425_sv2v_reg ;
  assign \nz.mem [424] = \nz.mem_424_sv2v_reg ;
  assign \nz.mem [423] = \nz.mem_423_sv2v_reg ;
  assign \nz.mem [422] = \nz.mem_422_sv2v_reg ;
  assign \nz.mem [421] = \nz.mem_421_sv2v_reg ;
  assign \nz.mem [420] = \nz.mem_420_sv2v_reg ;
  assign \nz.mem [419] = \nz.mem_419_sv2v_reg ;
  assign \nz.mem [418] = \nz.mem_418_sv2v_reg ;
  assign \nz.mem [417] = \nz.mem_417_sv2v_reg ;
  assign \nz.mem [416] = \nz.mem_416_sv2v_reg ;
  assign \nz.mem [415] = \nz.mem_415_sv2v_reg ;
  assign \nz.mem [414] = \nz.mem_414_sv2v_reg ;
  assign \nz.mem [413] = \nz.mem_413_sv2v_reg ;
  assign \nz.mem [412] = \nz.mem_412_sv2v_reg ;
  assign \nz.mem [411] = \nz.mem_411_sv2v_reg ;
  assign \nz.mem [410] = \nz.mem_410_sv2v_reg ;
  assign \nz.mem [409] = \nz.mem_409_sv2v_reg ;
  assign \nz.mem [408] = \nz.mem_408_sv2v_reg ;
  assign \nz.mem [407] = \nz.mem_407_sv2v_reg ;
  assign \nz.mem [406] = \nz.mem_406_sv2v_reg ;
  assign \nz.mem [405] = \nz.mem_405_sv2v_reg ;
  assign \nz.mem [404] = \nz.mem_404_sv2v_reg ;
  assign \nz.mem [403] = \nz.mem_403_sv2v_reg ;
  assign \nz.mem [402] = \nz.mem_402_sv2v_reg ;
  assign \nz.mem [401] = \nz.mem_401_sv2v_reg ;
  assign \nz.mem [400] = \nz.mem_400_sv2v_reg ;
  assign \nz.mem [399] = \nz.mem_399_sv2v_reg ;
  assign \nz.mem [398] = \nz.mem_398_sv2v_reg ;
  assign \nz.mem [397] = \nz.mem_397_sv2v_reg ;
  assign \nz.mem [396] = \nz.mem_396_sv2v_reg ;
  assign \nz.mem [395] = \nz.mem_395_sv2v_reg ;
  assign \nz.mem [394] = \nz.mem_394_sv2v_reg ;
  assign \nz.mem [393] = \nz.mem_393_sv2v_reg ;
  assign \nz.mem [392] = \nz.mem_392_sv2v_reg ;
  assign \nz.mem [391] = \nz.mem_391_sv2v_reg ;
  assign \nz.mem [390] = \nz.mem_390_sv2v_reg ;
  assign \nz.mem [389] = \nz.mem_389_sv2v_reg ;
  assign \nz.mem [388] = \nz.mem_388_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[79] = (N17)? \nz.mem [79] : 
                        (N19)? \nz.mem [159] : 
                        (N21)? \nz.mem [239] : 
                        (N23)? \nz.mem [319] : 
                        (N18)? \nz.mem [399] : 
                        (N20)? \nz.mem [479] : 
                        (N22)? \nz.mem [559] : 
                        (N24)? \nz.mem [639] : 1'b0;
  assign r_data_o[78] = (N17)? \nz.mem [78] : 
                        (N19)? \nz.mem [158] : 
                        (N21)? \nz.mem [238] : 
                        (N23)? \nz.mem [318] : 
                        (N18)? \nz.mem [398] : 
                        (N20)? \nz.mem [478] : 
                        (N22)? \nz.mem [558] : 
                        (N24)? \nz.mem [638] : 1'b0;
  assign r_data_o[77] = (N17)? \nz.mem [77] : 
                        (N19)? \nz.mem [157] : 
                        (N21)? \nz.mem [237] : 
                        (N23)? \nz.mem [317] : 
                        (N18)? \nz.mem [397] : 
                        (N20)? \nz.mem [477] : 
                        (N22)? \nz.mem [557] : 
                        (N24)? \nz.mem [637] : 1'b0;
  assign r_data_o[76] = (N17)? \nz.mem [76] : 
                        (N19)? \nz.mem [156] : 
                        (N21)? \nz.mem [236] : 
                        (N23)? \nz.mem [316] : 
                        (N18)? \nz.mem [396] : 
                        (N20)? \nz.mem [476] : 
                        (N22)? \nz.mem [556] : 
                        (N24)? \nz.mem [636] : 1'b0;
  assign r_data_o[75] = (N17)? \nz.mem [75] : 
                        (N19)? \nz.mem [155] : 
                        (N21)? \nz.mem [235] : 
                        (N23)? \nz.mem [315] : 
                        (N18)? \nz.mem [395] : 
                        (N20)? \nz.mem [475] : 
                        (N22)? \nz.mem [555] : 
                        (N24)? \nz.mem [635] : 1'b0;
  assign r_data_o[74] = (N17)? \nz.mem [74] : 
                        (N19)? \nz.mem [154] : 
                        (N21)? \nz.mem [234] : 
                        (N23)? \nz.mem [314] : 
                        (N18)? \nz.mem [394] : 
                        (N20)? \nz.mem [474] : 
                        (N22)? \nz.mem [554] : 
                        (N24)? \nz.mem [634] : 1'b0;
  assign r_data_o[73] = (N17)? \nz.mem [73] : 
                        (N19)? \nz.mem [153] : 
                        (N21)? \nz.mem [233] : 
                        (N23)? \nz.mem [313] : 
                        (N18)? \nz.mem [393] : 
                        (N20)? \nz.mem [473] : 
                        (N22)? \nz.mem [553] : 
                        (N24)? \nz.mem [633] : 1'b0;
  assign r_data_o[72] = (N17)? \nz.mem [72] : 
                        (N19)? \nz.mem [152] : 
                        (N21)? \nz.mem [232] : 
                        (N23)? \nz.mem [312] : 
                        (N18)? \nz.mem [392] : 
                        (N20)? \nz.mem [472] : 
                        (N22)? \nz.mem [552] : 
                        (N24)? \nz.mem [632] : 1'b0;
  assign r_data_o[71] = (N17)? \nz.mem [71] : 
                        (N19)? \nz.mem [151] : 
                        (N21)? \nz.mem [231] : 
                        (N23)? \nz.mem [311] : 
                        (N18)? \nz.mem [391] : 
                        (N20)? \nz.mem [471] : 
                        (N22)? \nz.mem [551] : 
                        (N24)? \nz.mem [631] : 1'b0;
  assign r_data_o[70] = (N17)? \nz.mem [70] : 
                        (N19)? \nz.mem [150] : 
                        (N21)? \nz.mem [230] : 
                        (N23)? \nz.mem [310] : 
                        (N18)? \nz.mem [390] : 
                        (N20)? \nz.mem [470] : 
                        (N22)? \nz.mem [550] : 
                        (N24)? \nz.mem [630] : 1'b0;
  assign r_data_o[69] = (N17)? \nz.mem [69] : 
                        (N19)? \nz.mem [149] : 
                        (N21)? \nz.mem [229] : 
                        (N23)? \nz.mem [309] : 
                        (N18)? \nz.mem [389] : 
                        (N20)? \nz.mem [469] : 
                        (N22)? \nz.mem [549] : 
                        (N24)? \nz.mem [629] : 1'b0;
  assign r_data_o[68] = (N17)? \nz.mem [68] : 
                        (N19)? \nz.mem [148] : 
                        (N21)? \nz.mem [228] : 
                        (N23)? \nz.mem [308] : 
                        (N18)? \nz.mem [388] : 
                        (N20)? \nz.mem [468] : 
                        (N22)? \nz.mem [548] : 
                        (N24)? \nz.mem [628] : 1'b0;
  assign r_data_o[67] = (N17)? \nz.mem [67] : 
                        (N19)? \nz.mem [147] : 
                        (N21)? \nz.mem [227] : 
                        (N23)? \nz.mem [307] : 
                        (N18)? \nz.mem [387] : 
                        (N20)? \nz.mem [467] : 
                        (N22)? \nz.mem [547] : 
                        (N24)? \nz.mem [627] : 1'b0;
  assign r_data_o[66] = (N17)? \nz.mem [66] : 
                        (N19)? \nz.mem [146] : 
                        (N21)? \nz.mem [226] : 
                        (N23)? \nz.mem [306] : 
                        (N18)? \nz.mem [386] : 
                        (N20)? \nz.mem [466] : 
                        (N22)? \nz.mem [546] : 
                        (N24)? \nz.mem [626] : 1'b0;
  assign r_data_o[65] = (N17)? \nz.mem [65] : 
                        (N19)? \nz.mem [145] : 
                        (N21)? \nz.mem [225] : 
                        (N23)? \nz.mem [305] : 
                        (N18)? \nz.mem [385] : 
                        (N20)? \nz.mem [465] : 
                        (N22)? \nz.mem [545] : 
                        (N24)? \nz.mem [625] : 1'b0;
  assign r_data_o[64] = (N17)? \nz.mem [64] : 
                        (N19)? \nz.mem [144] : 
                        (N21)? \nz.mem [224] : 
                        (N23)? \nz.mem [304] : 
                        (N18)? \nz.mem [384] : 
                        (N20)? \nz.mem [464] : 
                        (N22)? \nz.mem [544] : 
                        (N24)? \nz.mem [624] : 1'b0;
  assign r_data_o[63] = (N17)? \nz.mem [63] : 
                        (N19)? \nz.mem [143] : 
                        (N21)? \nz.mem [223] : 
                        (N23)? \nz.mem [303] : 
                        (N18)? \nz.mem [383] : 
                        (N20)? \nz.mem [463] : 
                        (N22)? \nz.mem [543] : 
                        (N24)? \nz.mem [623] : 1'b0;
  assign r_data_o[62] = (N17)? \nz.mem [62] : 
                        (N19)? \nz.mem [142] : 
                        (N21)? \nz.mem [222] : 
                        (N23)? \nz.mem [302] : 
                        (N18)? \nz.mem [382] : 
                        (N20)? \nz.mem [462] : 
                        (N22)? \nz.mem [542] : 
                        (N24)? \nz.mem [622] : 1'b0;
  assign r_data_o[61] = (N17)? \nz.mem [61] : 
                        (N19)? \nz.mem [141] : 
                        (N21)? \nz.mem [221] : 
                        (N23)? \nz.mem [301] : 
                        (N18)? \nz.mem [381] : 
                        (N20)? \nz.mem [461] : 
                        (N22)? \nz.mem [541] : 
                        (N24)? \nz.mem [621] : 1'b0;
  assign r_data_o[60] = (N17)? \nz.mem [60] : 
                        (N19)? \nz.mem [140] : 
                        (N21)? \nz.mem [220] : 
                        (N23)? \nz.mem [300] : 
                        (N18)? \nz.mem [380] : 
                        (N20)? \nz.mem [460] : 
                        (N22)? \nz.mem [540] : 
                        (N24)? \nz.mem [620] : 1'b0;
  assign r_data_o[59] = (N17)? \nz.mem [59] : 
                        (N19)? \nz.mem [139] : 
                        (N21)? \nz.mem [219] : 
                        (N23)? \nz.mem [299] : 
                        (N18)? \nz.mem [379] : 
                        (N20)? \nz.mem [459] : 
                        (N22)? \nz.mem [539] : 
                        (N24)? \nz.mem [619] : 1'b0;
  assign r_data_o[58] = (N17)? \nz.mem [58] : 
                        (N19)? \nz.mem [138] : 
                        (N21)? \nz.mem [218] : 
                        (N23)? \nz.mem [298] : 
                        (N18)? \nz.mem [378] : 
                        (N20)? \nz.mem [458] : 
                        (N22)? \nz.mem [538] : 
                        (N24)? \nz.mem [618] : 1'b0;
  assign r_data_o[57] = (N17)? \nz.mem [57] : 
                        (N19)? \nz.mem [137] : 
                        (N21)? \nz.mem [217] : 
                        (N23)? \nz.mem [297] : 
                        (N18)? \nz.mem [377] : 
                        (N20)? \nz.mem [457] : 
                        (N22)? \nz.mem [537] : 
                        (N24)? \nz.mem [617] : 1'b0;
  assign r_data_o[56] = (N17)? \nz.mem [56] : 
                        (N19)? \nz.mem [136] : 
                        (N21)? \nz.mem [216] : 
                        (N23)? \nz.mem [296] : 
                        (N18)? \nz.mem [376] : 
                        (N20)? \nz.mem [456] : 
                        (N22)? \nz.mem [536] : 
                        (N24)? \nz.mem [616] : 1'b0;
  assign r_data_o[55] = (N17)? \nz.mem [55] : 
                        (N19)? \nz.mem [135] : 
                        (N21)? \nz.mem [215] : 
                        (N23)? \nz.mem [295] : 
                        (N18)? \nz.mem [375] : 
                        (N20)? \nz.mem [455] : 
                        (N22)? \nz.mem [535] : 
                        (N24)? \nz.mem [615] : 1'b0;
  assign r_data_o[54] = (N17)? \nz.mem [54] : 
                        (N19)? \nz.mem [134] : 
                        (N21)? \nz.mem [214] : 
                        (N23)? \nz.mem [294] : 
                        (N18)? \nz.mem [374] : 
                        (N20)? \nz.mem [454] : 
                        (N22)? \nz.mem [534] : 
                        (N24)? \nz.mem [614] : 1'b0;
  assign r_data_o[53] = (N17)? \nz.mem [53] : 
                        (N19)? \nz.mem [133] : 
                        (N21)? \nz.mem [213] : 
                        (N23)? \nz.mem [293] : 
                        (N18)? \nz.mem [373] : 
                        (N20)? \nz.mem [453] : 
                        (N22)? \nz.mem [533] : 
                        (N24)? \nz.mem [613] : 1'b0;
  assign r_data_o[52] = (N17)? \nz.mem [52] : 
                        (N19)? \nz.mem [132] : 
                        (N21)? \nz.mem [212] : 
                        (N23)? \nz.mem [292] : 
                        (N18)? \nz.mem [372] : 
                        (N20)? \nz.mem [452] : 
                        (N22)? \nz.mem [532] : 
                        (N24)? \nz.mem [612] : 1'b0;
  assign r_data_o[51] = (N17)? \nz.mem [51] : 
                        (N19)? \nz.mem [131] : 
                        (N21)? \nz.mem [211] : 
                        (N23)? \nz.mem [291] : 
                        (N18)? \nz.mem [371] : 
                        (N20)? \nz.mem [451] : 
                        (N22)? \nz.mem [531] : 
                        (N24)? \nz.mem [611] : 1'b0;
  assign r_data_o[50] = (N17)? \nz.mem [50] : 
                        (N19)? \nz.mem [130] : 
                        (N21)? \nz.mem [210] : 
                        (N23)? \nz.mem [290] : 
                        (N18)? \nz.mem [370] : 
                        (N20)? \nz.mem [450] : 
                        (N22)? \nz.mem [530] : 
                        (N24)? \nz.mem [610] : 1'b0;
  assign r_data_o[49] = (N17)? \nz.mem [49] : 
                        (N19)? \nz.mem [129] : 
                        (N21)? \nz.mem [209] : 
                        (N23)? \nz.mem [289] : 
                        (N18)? \nz.mem [369] : 
                        (N20)? \nz.mem [449] : 
                        (N22)? \nz.mem [529] : 
                        (N24)? \nz.mem [609] : 1'b0;
  assign r_data_o[48] = (N17)? \nz.mem [48] : 
                        (N19)? \nz.mem [128] : 
                        (N21)? \nz.mem [208] : 
                        (N23)? \nz.mem [288] : 
                        (N18)? \nz.mem [368] : 
                        (N20)? \nz.mem [448] : 
                        (N22)? \nz.mem [528] : 
                        (N24)? \nz.mem [608] : 1'b0;
  assign r_data_o[47] = (N17)? \nz.mem [47] : 
                        (N19)? \nz.mem [127] : 
                        (N21)? \nz.mem [207] : 
                        (N23)? \nz.mem [287] : 
                        (N18)? \nz.mem [367] : 
                        (N20)? \nz.mem [447] : 
                        (N22)? \nz.mem [527] : 
                        (N24)? \nz.mem [607] : 1'b0;
  assign r_data_o[46] = (N17)? \nz.mem [46] : 
                        (N19)? \nz.mem [126] : 
                        (N21)? \nz.mem [206] : 
                        (N23)? \nz.mem [286] : 
                        (N18)? \nz.mem [366] : 
                        (N20)? \nz.mem [446] : 
                        (N22)? \nz.mem [526] : 
                        (N24)? \nz.mem [606] : 1'b0;
  assign r_data_o[45] = (N17)? \nz.mem [45] : 
                        (N19)? \nz.mem [125] : 
                        (N21)? \nz.mem [205] : 
                        (N23)? \nz.mem [285] : 
                        (N18)? \nz.mem [365] : 
                        (N20)? \nz.mem [445] : 
                        (N22)? \nz.mem [525] : 
                        (N24)? \nz.mem [605] : 1'b0;
  assign r_data_o[44] = (N17)? \nz.mem [44] : 
                        (N19)? \nz.mem [124] : 
                        (N21)? \nz.mem [204] : 
                        (N23)? \nz.mem [284] : 
                        (N18)? \nz.mem [364] : 
                        (N20)? \nz.mem [444] : 
                        (N22)? \nz.mem [524] : 
                        (N24)? \nz.mem [604] : 1'b0;
  assign r_data_o[43] = (N17)? \nz.mem [43] : 
                        (N19)? \nz.mem [123] : 
                        (N21)? \nz.mem [203] : 
                        (N23)? \nz.mem [283] : 
                        (N18)? \nz.mem [363] : 
                        (N20)? \nz.mem [443] : 
                        (N22)? \nz.mem [523] : 
                        (N24)? \nz.mem [603] : 1'b0;
  assign r_data_o[42] = (N17)? \nz.mem [42] : 
                        (N19)? \nz.mem [122] : 
                        (N21)? \nz.mem [202] : 
                        (N23)? \nz.mem [282] : 
                        (N18)? \nz.mem [362] : 
                        (N20)? \nz.mem [442] : 
                        (N22)? \nz.mem [522] : 
                        (N24)? \nz.mem [602] : 1'b0;
  assign r_data_o[41] = (N17)? \nz.mem [41] : 
                        (N19)? \nz.mem [121] : 
                        (N21)? \nz.mem [201] : 
                        (N23)? \nz.mem [281] : 
                        (N18)? \nz.mem [361] : 
                        (N20)? \nz.mem [441] : 
                        (N22)? \nz.mem [521] : 
                        (N24)? \nz.mem [601] : 1'b0;
  assign r_data_o[40] = (N17)? \nz.mem [40] : 
                        (N19)? \nz.mem [120] : 
                        (N21)? \nz.mem [200] : 
                        (N23)? \nz.mem [280] : 
                        (N18)? \nz.mem [360] : 
                        (N20)? \nz.mem [440] : 
                        (N22)? \nz.mem [520] : 
                        (N24)? \nz.mem [600] : 1'b0;
  assign r_data_o[39] = (N17)? \nz.mem [39] : 
                        (N19)? \nz.mem [119] : 
                        (N21)? \nz.mem [199] : 
                        (N23)? \nz.mem [279] : 
                        (N18)? \nz.mem [359] : 
                        (N20)? \nz.mem [439] : 
                        (N22)? \nz.mem [519] : 
                        (N24)? \nz.mem [599] : 1'b0;
  assign r_data_o[38] = (N17)? \nz.mem [38] : 
                        (N19)? \nz.mem [118] : 
                        (N21)? \nz.mem [198] : 
                        (N23)? \nz.mem [278] : 
                        (N18)? \nz.mem [358] : 
                        (N20)? \nz.mem [438] : 
                        (N22)? \nz.mem [518] : 
                        (N24)? \nz.mem [598] : 1'b0;
  assign r_data_o[37] = (N17)? \nz.mem [37] : 
                        (N19)? \nz.mem [117] : 
                        (N21)? \nz.mem [197] : 
                        (N23)? \nz.mem [277] : 
                        (N18)? \nz.mem [357] : 
                        (N20)? \nz.mem [437] : 
                        (N22)? \nz.mem [517] : 
                        (N24)? \nz.mem [597] : 1'b0;
  assign r_data_o[36] = (N17)? \nz.mem [36] : 
                        (N19)? \nz.mem [116] : 
                        (N21)? \nz.mem [196] : 
                        (N23)? \nz.mem [276] : 
                        (N18)? \nz.mem [356] : 
                        (N20)? \nz.mem [436] : 
                        (N22)? \nz.mem [516] : 
                        (N24)? \nz.mem [596] : 1'b0;
  assign r_data_o[35] = (N17)? \nz.mem [35] : 
                        (N19)? \nz.mem [115] : 
                        (N21)? \nz.mem [195] : 
                        (N23)? \nz.mem [275] : 
                        (N18)? \nz.mem [355] : 
                        (N20)? \nz.mem [435] : 
                        (N22)? \nz.mem [515] : 
                        (N24)? \nz.mem [595] : 1'b0;
  assign r_data_o[34] = (N17)? \nz.mem [34] : 
                        (N19)? \nz.mem [114] : 
                        (N21)? \nz.mem [194] : 
                        (N23)? \nz.mem [274] : 
                        (N18)? \nz.mem [354] : 
                        (N20)? \nz.mem [434] : 
                        (N22)? \nz.mem [514] : 
                        (N24)? \nz.mem [594] : 1'b0;
  assign r_data_o[33] = (N17)? \nz.mem [33] : 
                        (N19)? \nz.mem [113] : 
                        (N21)? \nz.mem [193] : 
                        (N23)? \nz.mem [273] : 
                        (N18)? \nz.mem [353] : 
                        (N20)? \nz.mem [433] : 
                        (N22)? \nz.mem [513] : 
                        (N24)? \nz.mem [593] : 1'b0;
  assign r_data_o[32] = (N17)? \nz.mem [32] : 
                        (N19)? \nz.mem [112] : 
                        (N21)? \nz.mem [192] : 
                        (N23)? \nz.mem [272] : 
                        (N18)? \nz.mem [352] : 
                        (N20)? \nz.mem [432] : 
                        (N22)? \nz.mem [512] : 
                        (N24)? \nz.mem [592] : 1'b0;
  assign r_data_o[31] = (N17)? \nz.mem [31] : 
                        (N19)? \nz.mem [111] : 
                        (N21)? \nz.mem [191] : 
                        (N23)? \nz.mem [271] : 
                        (N18)? \nz.mem [351] : 
                        (N20)? \nz.mem [431] : 
                        (N22)? \nz.mem [511] : 
                        (N24)? \nz.mem [591] : 1'b0;
  assign r_data_o[30] = (N17)? \nz.mem [30] : 
                        (N19)? \nz.mem [110] : 
                        (N21)? \nz.mem [190] : 
                        (N23)? \nz.mem [270] : 
                        (N18)? \nz.mem [350] : 
                        (N20)? \nz.mem [430] : 
                        (N22)? \nz.mem [510] : 
                        (N24)? \nz.mem [590] : 1'b0;
  assign r_data_o[29] = (N17)? \nz.mem [29] : 
                        (N19)? \nz.mem [109] : 
                        (N21)? \nz.mem [189] : 
                        (N23)? \nz.mem [269] : 
                        (N18)? \nz.mem [349] : 
                        (N20)? \nz.mem [429] : 
                        (N22)? \nz.mem [509] : 
                        (N24)? \nz.mem [589] : 1'b0;
  assign r_data_o[28] = (N17)? \nz.mem [28] : 
                        (N19)? \nz.mem [108] : 
                        (N21)? \nz.mem [188] : 
                        (N23)? \nz.mem [268] : 
                        (N18)? \nz.mem [348] : 
                        (N20)? \nz.mem [428] : 
                        (N22)? \nz.mem [508] : 
                        (N24)? \nz.mem [588] : 1'b0;
  assign r_data_o[27] = (N17)? \nz.mem [27] : 
                        (N19)? \nz.mem [107] : 
                        (N21)? \nz.mem [187] : 
                        (N23)? \nz.mem [267] : 
                        (N18)? \nz.mem [347] : 
                        (N20)? \nz.mem [427] : 
                        (N22)? \nz.mem [507] : 
                        (N24)? \nz.mem [587] : 1'b0;
  assign r_data_o[26] = (N17)? \nz.mem [26] : 
                        (N19)? \nz.mem [106] : 
                        (N21)? \nz.mem [186] : 
                        (N23)? \nz.mem [266] : 
                        (N18)? \nz.mem [346] : 
                        (N20)? \nz.mem [426] : 
                        (N22)? \nz.mem [506] : 
                        (N24)? \nz.mem [586] : 1'b0;
  assign r_data_o[25] = (N17)? \nz.mem [25] : 
                        (N19)? \nz.mem [105] : 
                        (N21)? \nz.mem [185] : 
                        (N23)? \nz.mem [265] : 
                        (N18)? \nz.mem [345] : 
                        (N20)? \nz.mem [425] : 
                        (N22)? \nz.mem [505] : 
                        (N24)? \nz.mem [585] : 1'b0;
  assign r_data_o[24] = (N17)? \nz.mem [24] : 
                        (N19)? \nz.mem [104] : 
                        (N21)? \nz.mem [184] : 
                        (N23)? \nz.mem [264] : 
                        (N18)? \nz.mem [344] : 
                        (N20)? \nz.mem [424] : 
                        (N22)? \nz.mem [504] : 
                        (N24)? \nz.mem [584] : 1'b0;
  assign r_data_o[23] = (N17)? \nz.mem [23] : 
                        (N19)? \nz.mem [103] : 
                        (N21)? \nz.mem [183] : 
                        (N23)? \nz.mem [263] : 
                        (N18)? \nz.mem [343] : 
                        (N20)? \nz.mem [423] : 
                        (N22)? \nz.mem [503] : 
                        (N24)? \nz.mem [583] : 1'b0;
  assign r_data_o[22] = (N17)? \nz.mem [22] : 
                        (N19)? \nz.mem [102] : 
                        (N21)? \nz.mem [182] : 
                        (N23)? \nz.mem [262] : 
                        (N18)? \nz.mem [342] : 
                        (N20)? \nz.mem [422] : 
                        (N22)? \nz.mem [502] : 
                        (N24)? \nz.mem [582] : 1'b0;
  assign r_data_o[21] = (N17)? \nz.mem [21] : 
                        (N19)? \nz.mem [101] : 
                        (N21)? \nz.mem [181] : 
                        (N23)? \nz.mem [261] : 
                        (N18)? \nz.mem [341] : 
                        (N20)? \nz.mem [421] : 
                        (N22)? \nz.mem [501] : 
                        (N24)? \nz.mem [581] : 1'b0;
  assign r_data_o[20] = (N17)? \nz.mem [20] : 
                        (N19)? \nz.mem [100] : 
                        (N21)? \nz.mem [180] : 
                        (N23)? \nz.mem [260] : 
                        (N18)? \nz.mem [340] : 
                        (N20)? \nz.mem [420] : 
                        (N22)? \nz.mem [500] : 
                        (N24)? \nz.mem [580] : 1'b0;
  assign r_data_o[19] = (N17)? \nz.mem [19] : 
                        (N19)? \nz.mem [99] : 
                        (N21)? \nz.mem [179] : 
                        (N23)? \nz.mem [259] : 
                        (N18)? \nz.mem [339] : 
                        (N20)? \nz.mem [419] : 
                        (N22)? \nz.mem [499] : 
                        (N24)? \nz.mem [579] : 1'b0;
  assign r_data_o[18] = (N17)? \nz.mem [18] : 
                        (N19)? \nz.mem [98] : 
                        (N21)? \nz.mem [178] : 
                        (N23)? \nz.mem [258] : 
                        (N18)? \nz.mem [338] : 
                        (N20)? \nz.mem [418] : 
                        (N22)? \nz.mem [498] : 
                        (N24)? \nz.mem [578] : 1'b0;
  assign r_data_o[17] = (N17)? \nz.mem [17] : 
                        (N19)? \nz.mem [97] : 
                        (N21)? \nz.mem [177] : 
                        (N23)? \nz.mem [257] : 
                        (N18)? \nz.mem [337] : 
                        (N20)? \nz.mem [417] : 
                        (N22)? \nz.mem [497] : 
                        (N24)? \nz.mem [577] : 1'b0;
  assign r_data_o[16] = (N17)? \nz.mem [16] : 
                        (N19)? \nz.mem [96] : 
                        (N21)? \nz.mem [176] : 
                        (N23)? \nz.mem [256] : 
                        (N18)? \nz.mem [336] : 
                        (N20)? \nz.mem [416] : 
                        (N22)? \nz.mem [496] : 
                        (N24)? \nz.mem [576] : 1'b0;
  assign r_data_o[15] = (N17)? \nz.mem [15] : 
                        (N19)? \nz.mem [95] : 
                        (N21)? \nz.mem [175] : 
                        (N23)? \nz.mem [255] : 
                        (N18)? \nz.mem [335] : 
                        (N20)? \nz.mem [415] : 
                        (N22)? \nz.mem [495] : 
                        (N24)? \nz.mem [575] : 1'b0;
  assign r_data_o[14] = (N17)? \nz.mem [14] : 
                        (N19)? \nz.mem [94] : 
                        (N21)? \nz.mem [174] : 
                        (N23)? \nz.mem [254] : 
                        (N18)? \nz.mem [334] : 
                        (N20)? \nz.mem [414] : 
                        (N22)? \nz.mem [494] : 
                        (N24)? \nz.mem [574] : 1'b0;
  assign r_data_o[13] = (N17)? \nz.mem [13] : 
                        (N19)? \nz.mem [93] : 
                        (N21)? \nz.mem [173] : 
                        (N23)? \nz.mem [253] : 
                        (N18)? \nz.mem [333] : 
                        (N20)? \nz.mem [413] : 
                        (N22)? \nz.mem [493] : 
                        (N24)? \nz.mem [573] : 1'b0;
  assign r_data_o[12] = (N17)? \nz.mem [12] : 
                        (N19)? \nz.mem [92] : 
                        (N21)? \nz.mem [172] : 
                        (N23)? \nz.mem [252] : 
                        (N18)? \nz.mem [332] : 
                        (N20)? \nz.mem [412] : 
                        (N22)? \nz.mem [492] : 
                        (N24)? \nz.mem [572] : 1'b0;
  assign r_data_o[11] = (N17)? \nz.mem [11] : 
                        (N19)? \nz.mem [91] : 
                        (N21)? \nz.mem [171] : 
                        (N23)? \nz.mem [251] : 
                        (N18)? \nz.mem [331] : 
                        (N20)? \nz.mem [411] : 
                        (N22)? \nz.mem [491] : 
                        (N24)? \nz.mem [571] : 1'b0;
  assign r_data_o[10] = (N17)? \nz.mem [10] : 
                        (N19)? \nz.mem [90] : 
                        (N21)? \nz.mem [170] : 
                        (N23)? \nz.mem [250] : 
                        (N18)? \nz.mem [330] : 
                        (N20)? \nz.mem [410] : 
                        (N22)? \nz.mem [490] : 
                        (N24)? \nz.mem [570] : 1'b0;
  assign r_data_o[9] = (N17)? \nz.mem [9] : 
                       (N19)? \nz.mem [89] : 
                       (N21)? \nz.mem [169] : 
                       (N23)? \nz.mem [249] : 
                       (N18)? \nz.mem [329] : 
                       (N20)? \nz.mem [409] : 
                       (N22)? \nz.mem [489] : 
                       (N24)? \nz.mem [569] : 1'b0;
  assign r_data_o[8] = (N17)? \nz.mem [8] : 
                       (N19)? \nz.mem [88] : 
                       (N21)? \nz.mem [168] : 
                       (N23)? \nz.mem [248] : 
                       (N18)? \nz.mem [328] : 
                       (N20)? \nz.mem [408] : 
                       (N22)? \nz.mem [488] : 
                       (N24)? \nz.mem [568] : 1'b0;
  assign r_data_o[7] = (N17)? \nz.mem [7] : 
                       (N19)? \nz.mem [87] : 
                       (N21)? \nz.mem [167] : 
                       (N23)? \nz.mem [247] : 
                       (N18)? \nz.mem [327] : 
                       (N20)? \nz.mem [407] : 
                       (N22)? \nz.mem [487] : 
                       (N24)? \nz.mem [567] : 1'b0;
  assign r_data_o[6] = (N17)? \nz.mem [6] : 
                       (N19)? \nz.mem [86] : 
                       (N21)? \nz.mem [166] : 
                       (N23)? \nz.mem [246] : 
                       (N18)? \nz.mem [326] : 
                       (N20)? \nz.mem [406] : 
                       (N22)? \nz.mem [486] : 
                       (N24)? \nz.mem [566] : 1'b0;
  assign r_data_o[5] = (N17)? \nz.mem [5] : 
                       (N19)? \nz.mem [85] : 
                       (N21)? \nz.mem [165] : 
                       (N23)? \nz.mem [245] : 
                       (N18)? \nz.mem [325] : 
                       (N20)? \nz.mem [405] : 
                       (N22)? \nz.mem [485] : 
                       (N24)? \nz.mem [565] : 1'b0;
  assign r_data_o[4] = (N17)? \nz.mem [4] : 
                       (N19)? \nz.mem [84] : 
                       (N21)? \nz.mem [164] : 
                       (N23)? \nz.mem [244] : 
                       (N18)? \nz.mem [324] : 
                       (N20)? \nz.mem [404] : 
                       (N22)? \nz.mem [484] : 
                       (N24)? \nz.mem [564] : 1'b0;
  assign r_data_o[3] = (N17)? \nz.mem [3] : 
                       (N19)? \nz.mem [83] : 
                       (N21)? \nz.mem [163] : 
                       (N23)? \nz.mem [243] : 
                       (N18)? \nz.mem [323] : 
                       (N20)? \nz.mem [403] : 
                       (N22)? \nz.mem [483] : 
                       (N24)? \nz.mem [563] : 1'b0;
  assign r_data_o[2] = (N17)? \nz.mem [2] : 
                       (N19)? \nz.mem [82] : 
                       (N21)? \nz.mem [162] : 
                       (N23)? \nz.mem [242] : 
                       (N18)? \nz.mem [322] : 
                       (N20)? \nz.mem [402] : 
                       (N22)? \nz.mem [482] : 
                       (N24)? \nz.mem [562] : 1'b0;
  assign r_data_o[1] = (N17)? \nz.mem [1] : 
                       (N19)? \nz.mem [81] : 
                       (N21)? \nz.mem [161] : 
                       (N23)? \nz.mem [241] : 
                       (N18)? \nz.mem [321] : 
                       (N20)? \nz.mem [401] : 
                       (N22)? \nz.mem [481] : 
                       (N24)? \nz.mem [561] : 1'b0;
  assign r_data_o[0] = (N17)? \nz.mem [0] : 
                       (N19)? \nz.mem [80] : 
                       (N21)? \nz.mem [160] : 
                       (N23)? \nz.mem [240] : 
                       (N18)? \nz.mem [320] : 
                       (N20)? \nz.mem [400] : 
                       (N22)? \nz.mem [480] : 
                       (N24)? \nz.mem [560] : 1'b0;
  assign N42 = w_addr_i[0] & w_addr_i[1];
  assign N33 = N42 & w_addr_i[2];
  assign N43 = N0 & w_addr_i[1];
  assign N0 = ~w_addr_i[0];
  assign N32 = N43 & w_addr_i[2];
  assign N44 = w_addr_i[0] & N1;
  assign N1 = ~w_addr_i[1];
  assign N31 = N44 & w_addr_i[2];
  assign N45 = N2 & N3;
  assign N2 = ~w_addr_i[0];
  assign N3 = ~w_addr_i[1];
  assign N30 = N45 & w_addr_i[2];
  assign N29 = N42 & N4;
  assign N4 = ~w_addr_i[2];
  assign N28 = N43 & N5;
  assign N5 = ~w_addr_i[2];
  assign N27 = N44 & N6;
  assign N6 = ~w_addr_i[2];
  assign N26 = N45 & N7;
  assign N7 = ~w_addr_i[2];
  assign { N41, N40, N39, N38, N37, N36, N35, N34 } = (N8)? { N33, N32, N31, N30, N29, N28, N27, N26 } : 
                                                      (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N25;
  assign N10 = ~r_addr_i[0];
  assign N11 = ~r_addr_i[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r_addr_i[1];
  assign N14 = r_addr_i[0] & N11;
  assign N15 = r_addr_i[0] & r_addr_i[1];
  assign N16 = ~r_addr_i[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r_addr_i[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r_addr_i[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r_addr_i[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r_addr_i[2];
  assign N25 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N41) begin
      \nz.mem_639_sv2v_reg  <= w_data_i[79];
      \nz.mem_638_sv2v_reg  <= w_data_i[78];
      \nz.mem_637_sv2v_reg  <= w_data_i[77];
      \nz.mem_636_sv2v_reg  <= w_data_i[76];
      \nz.mem_635_sv2v_reg  <= w_data_i[75];
      \nz.mem_634_sv2v_reg  <= w_data_i[74];
      \nz.mem_633_sv2v_reg  <= w_data_i[73];
      \nz.mem_632_sv2v_reg  <= w_data_i[72];
      \nz.mem_631_sv2v_reg  <= w_data_i[71];
      \nz.mem_630_sv2v_reg  <= w_data_i[70];
      \nz.mem_629_sv2v_reg  <= w_data_i[69];
      \nz.mem_628_sv2v_reg  <= w_data_i[68];
      \nz.mem_627_sv2v_reg  <= w_data_i[67];
      \nz.mem_626_sv2v_reg  <= w_data_i[66];
      \nz.mem_625_sv2v_reg  <= w_data_i[65];
      \nz.mem_624_sv2v_reg  <= w_data_i[64];
      \nz.mem_623_sv2v_reg  <= w_data_i[63];
      \nz.mem_622_sv2v_reg  <= w_data_i[62];
      \nz.mem_621_sv2v_reg  <= w_data_i[61];
      \nz.mem_620_sv2v_reg  <= w_data_i[60];
      \nz.mem_619_sv2v_reg  <= w_data_i[59];
      \nz.mem_618_sv2v_reg  <= w_data_i[58];
      \nz.mem_617_sv2v_reg  <= w_data_i[57];
      \nz.mem_616_sv2v_reg  <= w_data_i[56];
      \nz.mem_615_sv2v_reg  <= w_data_i[55];
      \nz.mem_614_sv2v_reg  <= w_data_i[54];
      \nz.mem_613_sv2v_reg  <= w_data_i[53];
      \nz.mem_612_sv2v_reg  <= w_data_i[52];
      \nz.mem_611_sv2v_reg  <= w_data_i[51];
      \nz.mem_610_sv2v_reg  <= w_data_i[50];
      \nz.mem_609_sv2v_reg  <= w_data_i[49];
      \nz.mem_608_sv2v_reg  <= w_data_i[48];
      \nz.mem_607_sv2v_reg  <= w_data_i[47];
      \nz.mem_606_sv2v_reg  <= w_data_i[46];
      \nz.mem_605_sv2v_reg  <= w_data_i[45];
      \nz.mem_604_sv2v_reg  <= w_data_i[44];
      \nz.mem_603_sv2v_reg  <= w_data_i[43];
      \nz.mem_602_sv2v_reg  <= w_data_i[42];
      \nz.mem_601_sv2v_reg  <= w_data_i[41];
      \nz.mem_600_sv2v_reg  <= w_data_i[40];
      \nz.mem_599_sv2v_reg  <= w_data_i[39];
      \nz.mem_598_sv2v_reg  <= w_data_i[38];
      \nz.mem_597_sv2v_reg  <= w_data_i[37];
      \nz.mem_596_sv2v_reg  <= w_data_i[36];
      \nz.mem_595_sv2v_reg  <= w_data_i[35];
      \nz.mem_594_sv2v_reg  <= w_data_i[34];
      \nz.mem_593_sv2v_reg  <= w_data_i[33];
      \nz.mem_592_sv2v_reg  <= w_data_i[32];
      \nz.mem_591_sv2v_reg  <= w_data_i[31];
      \nz.mem_590_sv2v_reg  <= w_data_i[30];
      \nz.mem_589_sv2v_reg  <= w_data_i[29];
      \nz.mem_588_sv2v_reg  <= w_data_i[28];
      \nz.mem_587_sv2v_reg  <= w_data_i[27];
      \nz.mem_586_sv2v_reg  <= w_data_i[26];
      \nz.mem_585_sv2v_reg  <= w_data_i[25];
      \nz.mem_584_sv2v_reg  <= w_data_i[24];
      \nz.mem_583_sv2v_reg  <= w_data_i[23];
      \nz.mem_582_sv2v_reg  <= w_data_i[22];
      \nz.mem_581_sv2v_reg  <= w_data_i[21];
      \nz.mem_580_sv2v_reg  <= w_data_i[20];
      \nz.mem_579_sv2v_reg  <= w_data_i[19];
      \nz.mem_578_sv2v_reg  <= w_data_i[18];
      \nz.mem_577_sv2v_reg  <= w_data_i[17];
      \nz.mem_576_sv2v_reg  <= w_data_i[16];
      \nz.mem_575_sv2v_reg  <= w_data_i[15];
      \nz.mem_574_sv2v_reg  <= w_data_i[14];
      \nz.mem_573_sv2v_reg  <= w_data_i[13];
      \nz.mem_572_sv2v_reg  <= w_data_i[12];
      \nz.mem_571_sv2v_reg  <= w_data_i[11];
      \nz.mem_570_sv2v_reg  <= w_data_i[10];
      \nz.mem_569_sv2v_reg  <= w_data_i[9];
      \nz.mem_568_sv2v_reg  <= w_data_i[8];
      \nz.mem_567_sv2v_reg  <= w_data_i[7];
      \nz.mem_566_sv2v_reg  <= w_data_i[6];
      \nz.mem_565_sv2v_reg  <= w_data_i[5];
      \nz.mem_564_sv2v_reg  <= w_data_i[4];
      \nz.mem_563_sv2v_reg  <= w_data_i[3];
      \nz.mem_562_sv2v_reg  <= w_data_i[2];
      \nz.mem_561_sv2v_reg  <= w_data_i[1];
      \nz.mem_560_sv2v_reg  <= w_data_i[0];
    end 
    if(N40) begin
      \nz.mem_559_sv2v_reg  <= w_data_i[79];
      \nz.mem_558_sv2v_reg  <= w_data_i[78];
      \nz.mem_557_sv2v_reg  <= w_data_i[77];
      \nz.mem_556_sv2v_reg  <= w_data_i[76];
      \nz.mem_555_sv2v_reg  <= w_data_i[75];
      \nz.mem_554_sv2v_reg  <= w_data_i[74];
      \nz.mem_553_sv2v_reg  <= w_data_i[73];
      \nz.mem_552_sv2v_reg  <= w_data_i[72];
      \nz.mem_551_sv2v_reg  <= w_data_i[71];
      \nz.mem_550_sv2v_reg  <= w_data_i[70];
      \nz.mem_549_sv2v_reg  <= w_data_i[69];
      \nz.mem_548_sv2v_reg  <= w_data_i[68];
      \nz.mem_547_sv2v_reg  <= w_data_i[67];
      \nz.mem_546_sv2v_reg  <= w_data_i[66];
      \nz.mem_545_sv2v_reg  <= w_data_i[65];
      \nz.mem_544_sv2v_reg  <= w_data_i[64];
      \nz.mem_543_sv2v_reg  <= w_data_i[63];
      \nz.mem_542_sv2v_reg  <= w_data_i[62];
      \nz.mem_541_sv2v_reg  <= w_data_i[61];
      \nz.mem_540_sv2v_reg  <= w_data_i[60];
      \nz.mem_539_sv2v_reg  <= w_data_i[59];
      \nz.mem_538_sv2v_reg  <= w_data_i[58];
      \nz.mem_537_sv2v_reg  <= w_data_i[57];
      \nz.mem_536_sv2v_reg  <= w_data_i[56];
      \nz.mem_535_sv2v_reg  <= w_data_i[55];
      \nz.mem_534_sv2v_reg  <= w_data_i[54];
      \nz.mem_533_sv2v_reg  <= w_data_i[53];
      \nz.mem_532_sv2v_reg  <= w_data_i[52];
      \nz.mem_531_sv2v_reg  <= w_data_i[51];
      \nz.mem_530_sv2v_reg  <= w_data_i[50];
      \nz.mem_529_sv2v_reg  <= w_data_i[49];
      \nz.mem_528_sv2v_reg  <= w_data_i[48];
      \nz.mem_527_sv2v_reg  <= w_data_i[47];
      \nz.mem_526_sv2v_reg  <= w_data_i[46];
      \nz.mem_525_sv2v_reg  <= w_data_i[45];
      \nz.mem_524_sv2v_reg  <= w_data_i[44];
      \nz.mem_523_sv2v_reg  <= w_data_i[43];
      \nz.mem_522_sv2v_reg  <= w_data_i[42];
      \nz.mem_521_sv2v_reg  <= w_data_i[41];
      \nz.mem_520_sv2v_reg  <= w_data_i[40];
      \nz.mem_519_sv2v_reg  <= w_data_i[39];
      \nz.mem_518_sv2v_reg  <= w_data_i[38];
      \nz.mem_517_sv2v_reg  <= w_data_i[37];
      \nz.mem_516_sv2v_reg  <= w_data_i[36];
      \nz.mem_515_sv2v_reg  <= w_data_i[35];
      \nz.mem_514_sv2v_reg  <= w_data_i[34];
      \nz.mem_513_sv2v_reg  <= w_data_i[33];
      \nz.mem_512_sv2v_reg  <= w_data_i[32];
      \nz.mem_511_sv2v_reg  <= w_data_i[31];
      \nz.mem_510_sv2v_reg  <= w_data_i[30];
      \nz.mem_509_sv2v_reg  <= w_data_i[29];
      \nz.mem_508_sv2v_reg  <= w_data_i[28];
      \nz.mem_507_sv2v_reg  <= w_data_i[27];
      \nz.mem_506_sv2v_reg  <= w_data_i[26];
      \nz.mem_505_sv2v_reg  <= w_data_i[25];
      \nz.mem_504_sv2v_reg  <= w_data_i[24];
      \nz.mem_503_sv2v_reg  <= w_data_i[23];
      \nz.mem_502_sv2v_reg  <= w_data_i[22];
      \nz.mem_501_sv2v_reg  <= w_data_i[21];
      \nz.mem_500_sv2v_reg  <= w_data_i[20];
      \nz.mem_499_sv2v_reg  <= w_data_i[19];
      \nz.mem_498_sv2v_reg  <= w_data_i[18];
      \nz.mem_497_sv2v_reg  <= w_data_i[17];
      \nz.mem_496_sv2v_reg  <= w_data_i[16];
      \nz.mem_495_sv2v_reg  <= w_data_i[15];
      \nz.mem_494_sv2v_reg  <= w_data_i[14];
      \nz.mem_493_sv2v_reg  <= w_data_i[13];
      \nz.mem_492_sv2v_reg  <= w_data_i[12];
      \nz.mem_491_sv2v_reg  <= w_data_i[11];
      \nz.mem_490_sv2v_reg  <= w_data_i[10];
      \nz.mem_489_sv2v_reg  <= w_data_i[9];
      \nz.mem_488_sv2v_reg  <= w_data_i[8];
      \nz.mem_487_sv2v_reg  <= w_data_i[7];
      \nz.mem_486_sv2v_reg  <= w_data_i[6];
      \nz.mem_485_sv2v_reg  <= w_data_i[5];
      \nz.mem_484_sv2v_reg  <= w_data_i[4];
      \nz.mem_483_sv2v_reg  <= w_data_i[3];
      \nz.mem_482_sv2v_reg  <= w_data_i[2];
      \nz.mem_481_sv2v_reg  <= w_data_i[1];
      \nz.mem_480_sv2v_reg  <= w_data_i[0];
    end 
    if(N39) begin
      \nz.mem_479_sv2v_reg  <= w_data_i[79];
      \nz.mem_478_sv2v_reg  <= w_data_i[78];
      \nz.mem_477_sv2v_reg  <= w_data_i[77];
      \nz.mem_476_sv2v_reg  <= w_data_i[76];
      \nz.mem_475_sv2v_reg  <= w_data_i[75];
      \nz.mem_474_sv2v_reg  <= w_data_i[74];
      \nz.mem_473_sv2v_reg  <= w_data_i[73];
      \nz.mem_472_sv2v_reg  <= w_data_i[72];
      \nz.mem_471_sv2v_reg  <= w_data_i[71];
      \nz.mem_470_sv2v_reg  <= w_data_i[70];
      \nz.mem_469_sv2v_reg  <= w_data_i[69];
      \nz.mem_468_sv2v_reg  <= w_data_i[68];
      \nz.mem_467_sv2v_reg  <= w_data_i[67];
      \nz.mem_466_sv2v_reg  <= w_data_i[66];
      \nz.mem_465_sv2v_reg  <= w_data_i[65];
      \nz.mem_464_sv2v_reg  <= w_data_i[64];
      \nz.mem_463_sv2v_reg  <= w_data_i[63];
      \nz.mem_462_sv2v_reg  <= w_data_i[62];
      \nz.mem_461_sv2v_reg  <= w_data_i[61];
      \nz.mem_460_sv2v_reg  <= w_data_i[60];
      \nz.mem_459_sv2v_reg  <= w_data_i[59];
      \nz.mem_458_sv2v_reg  <= w_data_i[58];
      \nz.mem_457_sv2v_reg  <= w_data_i[57];
      \nz.mem_456_sv2v_reg  <= w_data_i[56];
      \nz.mem_455_sv2v_reg  <= w_data_i[55];
      \nz.mem_454_sv2v_reg  <= w_data_i[54];
      \nz.mem_453_sv2v_reg  <= w_data_i[53];
      \nz.mem_452_sv2v_reg  <= w_data_i[52];
      \nz.mem_451_sv2v_reg  <= w_data_i[51];
      \nz.mem_450_sv2v_reg  <= w_data_i[50];
      \nz.mem_449_sv2v_reg  <= w_data_i[49];
      \nz.mem_448_sv2v_reg  <= w_data_i[48];
      \nz.mem_447_sv2v_reg  <= w_data_i[47];
      \nz.mem_446_sv2v_reg  <= w_data_i[46];
      \nz.mem_445_sv2v_reg  <= w_data_i[45];
      \nz.mem_444_sv2v_reg  <= w_data_i[44];
      \nz.mem_443_sv2v_reg  <= w_data_i[43];
      \nz.mem_442_sv2v_reg  <= w_data_i[42];
      \nz.mem_441_sv2v_reg  <= w_data_i[41];
      \nz.mem_440_sv2v_reg  <= w_data_i[40];
      \nz.mem_439_sv2v_reg  <= w_data_i[39];
      \nz.mem_438_sv2v_reg  <= w_data_i[38];
      \nz.mem_437_sv2v_reg  <= w_data_i[37];
      \nz.mem_436_sv2v_reg  <= w_data_i[36];
      \nz.mem_435_sv2v_reg  <= w_data_i[35];
      \nz.mem_434_sv2v_reg  <= w_data_i[34];
      \nz.mem_433_sv2v_reg  <= w_data_i[33];
      \nz.mem_432_sv2v_reg  <= w_data_i[32];
      \nz.mem_431_sv2v_reg  <= w_data_i[31];
      \nz.mem_430_sv2v_reg  <= w_data_i[30];
      \nz.mem_429_sv2v_reg  <= w_data_i[29];
      \nz.mem_428_sv2v_reg  <= w_data_i[28];
      \nz.mem_427_sv2v_reg  <= w_data_i[27];
      \nz.mem_426_sv2v_reg  <= w_data_i[26];
      \nz.mem_425_sv2v_reg  <= w_data_i[25];
      \nz.mem_424_sv2v_reg  <= w_data_i[24];
      \nz.mem_423_sv2v_reg  <= w_data_i[23];
      \nz.mem_422_sv2v_reg  <= w_data_i[22];
      \nz.mem_421_sv2v_reg  <= w_data_i[21];
      \nz.mem_420_sv2v_reg  <= w_data_i[20];
      \nz.mem_419_sv2v_reg  <= w_data_i[19];
      \nz.mem_418_sv2v_reg  <= w_data_i[18];
      \nz.mem_417_sv2v_reg  <= w_data_i[17];
      \nz.mem_416_sv2v_reg  <= w_data_i[16];
      \nz.mem_415_sv2v_reg  <= w_data_i[15];
      \nz.mem_414_sv2v_reg  <= w_data_i[14];
      \nz.mem_413_sv2v_reg  <= w_data_i[13];
      \nz.mem_412_sv2v_reg  <= w_data_i[12];
      \nz.mem_411_sv2v_reg  <= w_data_i[11];
      \nz.mem_410_sv2v_reg  <= w_data_i[10];
      \nz.mem_409_sv2v_reg  <= w_data_i[9];
      \nz.mem_408_sv2v_reg  <= w_data_i[8];
      \nz.mem_407_sv2v_reg  <= w_data_i[7];
      \nz.mem_406_sv2v_reg  <= w_data_i[6];
      \nz.mem_405_sv2v_reg  <= w_data_i[5];
      \nz.mem_404_sv2v_reg  <= w_data_i[4];
      \nz.mem_403_sv2v_reg  <= w_data_i[3];
      \nz.mem_402_sv2v_reg  <= w_data_i[2];
      \nz.mem_401_sv2v_reg  <= w_data_i[1];
      \nz.mem_400_sv2v_reg  <= w_data_i[0];
    end 
    if(N38) begin
      \nz.mem_399_sv2v_reg  <= w_data_i[79];
      \nz.mem_398_sv2v_reg  <= w_data_i[78];
      \nz.mem_397_sv2v_reg  <= w_data_i[77];
      \nz.mem_396_sv2v_reg  <= w_data_i[76];
      \nz.mem_395_sv2v_reg  <= w_data_i[75];
      \nz.mem_394_sv2v_reg  <= w_data_i[74];
      \nz.mem_393_sv2v_reg  <= w_data_i[73];
      \nz.mem_392_sv2v_reg  <= w_data_i[72];
      \nz.mem_391_sv2v_reg  <= w_data_i[71];
      \nz.mem_390_sv2v_reg  <= w_data_i[70];
      \nz.mem_389_sv2v_reg  <= w_data_i[69];
      \nz.mem_388_sv2v_reg  <= w_data_i[68];
      \nz.mem_387_sv2v_reg  <= w_data_i[67];
      \nz.mem_386_sv2v_reg  <= w_data_i[66];
      \nz.mem_385_sv2v_reg  <= w_data_i[65];
      \nz.mem_384_sv2v_reg  <= w_data_i[64];
      \nz.mem_383_sv2v_reg  <= w_data_i[63];
      \nz.mem_382_sv2v_reg  <= w_data_i[62];
      \nz.mem_381_sv2v_reg  <= w_data_i[61];
      \nz.mem_380_sv2v_reg  <= w_data_i[60];
      \nz.mem_379_sv2v_reg  <= w_data_i[59];
      \nz.mem_378_sv2v_reg  <= w_data_i[58];
      \nz.mem_377_sv2v_reg  <= w_data_i[57];
      \nz.mem_376_sv2v_reg  <= w_data_i[56];
      \nz.mem_375_sv2v_reg  <= w_data_i[55];
      \nz.mem_374_sv2v_reg  <= w_data_i[54];
      \nz.mem_373_sv2v_reg  <= w_data_i[53];
      \nz.mem_372_sv2v_reg  <= w_data_i[52];
      \nz.mem_371_sv2v_reg  <= w_data_i[51];
      \nz.mem_370_sv2v_reg  <= w_data_i[50];
      \nz.mem_369_sv2v_reg  <= w_data_i[49];
      \nz.mem_368_sv2v_reg  <= w_data_i[48];
      \nz.mem_367_sv2v_reg  <= w_data_i[47];
      \nz.mem_366_sv2v_reg  <= w_data_i[46];
      \nz.mem_365_sv2v_reg  <= w_data_i[45];
      \nz.mem_364_sv2v_reg  <= w_data_i[44];
      \nz.mem_363_sv2v_reg  <= w_data_i[43];
      \nz.mem_362_sv2v_reg  <= w_data_i[42];
      \nz.mem_361_sv2v_reg  <= w_data_i[41];
      \nz.mem_360_sv2v_reg  <= w_data_i[40];
      \nz.mem_359_sv2v_reg  <= w_data_i[39];
      \nz.mem_358_sv2v_reg  <= w_data_i[38];
      \nz.mem_357_sv2v_reg  <= w_data_i[37];
      \nz.mem_356_sv2v_reg  <= w_data_i[36];
      \nz.mem_355_sv2v_reg  <= w_data_i[35];
      \nz.mem_354_sv2v_reg  <= w_data_i[34];
      \nz.mem_353_sv2v_reg  <= w_data_i[33];
      \nz.mem_352_sv2v_reg  <= w_data_i[32];
      \nz.mem_351_sv2v_reg  <= w_data_i[31];
      \nz.mem_350_sv2v_reg  <= w_data_i[30];
      \nz.mem_349_sv2v_reg  <= w_data_i[29];
      \nz.mem_348_sv2v_reg  <= w_data_i[28];
      \nz.mem_347_sv2v_reg  <= w_data_i[27];
      \nz.mem_346_sv2v_reg  <= w_data_i[26];
      \nz.mem_345_sv2v_reg  <= w_data_i[25];
      \nz.mem_344_sv2v_reg  <= w_data_i[24];
      \nz.mem_343_sv2v_reg  <= w_data_i[23];
      \nz.mem_342_sv2v_reg  <= w_data_i[22];
      \nz.mem_341_sv2v_reg  <= w_data_i[21];
      \nz.mem_340_sv2v_reg  <= w_data_i[20];
      \nz.mem_339_sv2v_reg  <= w_data_i[19];
      \nz.mem_338_sv2v_reg  <= w_data_i[18];
      \nz.mem_337_sv2v_reg  <= w_data_i[17];
      \nz.mem_336_sv2v_reg  <= w_data_i[16];
      \nz.mem_335_sv2v_reg  <= w_data_i[15];
      \nz.mem_334_sv2v_reg  <= w_data_i[14];
      \nz.mem_333_sv2v_reg  <= w_data_i[13];
      \nz.mem_332_sv2v_reg  <= w_data_i[12];
      \nz.mem_331_sv2v_reg  <= w_data_i[11];
      \nz.mem_330_sv2v_reg  <= w_data_i[10];
      \nz.mem_329_sv2v_reg  <= w_data_i[9];
      \nz.mem_328_sv2v_reg  <= w_data_i[8];
      \nz.mem_327_sv2v_reg  <= w_data_i[7];
      \nz.mem_326_sv2v_reg  <= w_data_i[6];
      \nz.mem_325_sv2v_reg  <= w_data_i[5];
      \nz.mem_324_sv2v_reg  <= w_data_i[4];
      \nz.mem_323_sv2v_reg  <= w_data_i[3];
      \nz.mem_322_sv2v_reg  <= w_data_i[2];
      \nz.mem_321_sv2v_reg  <= w_data_i[1];
      \nz.mem_320_sv2v_reg  <= w_data_i[0];
    end 
    if(N37) begin
      \nz.mem_319_sv2v_reg  <= w_data_i[79];
      \nz.mem_318_sv2v_reg  <= w_data_i[78];
      \nz.mem_317_sv2v_reg  <= w_data_i[77];
      \nz.mem_316_sv2v_reg  <= w_data_i[76];
      \nz.mem_315_sv2v_reg  <= w_data_i[75];
      \nz.mem_314_sv2v_reg  <= w_data_i[74];
      \nz.mem_313_sv2v_reg  <= w_data_i[73];
      \nz.mem_312_sv2v_reg  <= w_data_i[72];
      \nz.mem_311_sv2v_reg  <= w_data_i[71];
      \nz.mem_310_sv2v_reg  <= w_data_i[70];
      \nz.mem_309_sv2v_reg  <= w_data_i[69];
      \nz.mem_308_sv2v_reg  <= w_data_i[68];
      \nz.mem_307_sv2v_reg  <= w_data_i[67];
      \nz.mem_306_sv2v_reg  <= w_data_i[66];
      \nz.mem_305_sv2v_reg  <= w_data_i[65];
      \nz.mem_304_sv2v_reg  <= w_data_i[64];
      \nz.mem_303_sv2v_reg  <= w_data_i[63];
      \nz.mem_302_sv2v_reg  <= w_data_i[62];
      \nz.mem_301_sv2v_reg  <= w_data_i[61];
      \nz.mem_300_sv2v_reg  <= w_data_i[60];
      \nz.mem_299_sv2v_reg  <= w_data_i[59];
      \nz.mem_298_sv2v_reg  <= w_data_i[58];
      \nz.mem_297_sv2v_reg  <= w_data_i[57];
      \nz.mem_296_sv2v_reg  <= w_data_i[56];
      \nz.mem_295_sv2v_reg  <= w_data_i[55];
      \nz.mem_294_sv2v_reg  <= w_data_i[54];
      \nz.mem_293_sv2v_reg  <= w_data_i[53];
      \nz.mem_292_sv2v_reg  <= w_data_i[52];
      \nz.mem_291_sv2v_reg  <= w_data_i[51];
      \nz.mem_290_sv2v_reg  <= w_data_i[50];
      \nz.mem_289_sv2v_reg  <= w_data_i[49];
      \nz.mem_288_sv2v_reg  <= w_data_i[48];
      \nz.mem_287_sv2v_reg  <= w_data_i[47];
      \nz.mem_286_sv2v_reg  <= w_data_i[46];
      \nz.mem_285_sv2v_reg  <= w_data_i[45];
      \nz.mem_284_sv2v_reg  <= w_data_i[44];
      \nz.mem_283_sv2v_reg  <= w_data_i[43];
      \nz.mem_282_sv2v_reg  <= w_data_i[42];
      \nz.mem_281_sv2v_reg  <= w_data_i[41];
      \nz.mem_280_sv2v_reg  <= w_data_i[40];
      \nz.mem_279_sv2v_reg  <= w_data_i[39];
      \nz.mem_278_sv2v_reg  <= w_data_i[38];
      \nz.mem_277_sv2v_reg  <= w_data_i[37];
      \nz.mem_276_sv2v_reg  <= w_data_i[36];
      \nz.mem_275_sv2v_reg  <= w_data_i[35];
      \nz.mem_274_sv2v_reg  <= w_data_i[34];
      \nz.mem_273_sv2v_reg  <= w_data_i[33];
      \nz.mem_272_sv2v_reg  <= w_data_i[32];
      \nz.mem_271_sv2v_reg  <= w_data_i[31];
      \nz.mem_270_sv2v_reg  <= w_data_i[30];
      \nz.mem_269_sv2v_reg  <= w_data_i[29];
      \nz.mem_268_sv2v_reg  <= w_data_i[28];
      \nz.mem_267_sv2v_reg  <= w_data_i[27];
      \nz.mem_266_sv2v_reg  <= w_data_i[26];
      \nz.mem_265_sv2v_reg  <= w_data_i[25];
      \nz.mem_264_sv2v_reg  <= w_data_i[24];
      \nz.mem_263_sv2v_reg  <= w_data_i[23];
      \nz.mem_262_sv2v_reg  <= w_data_i[22];
      \nz.mem_261_sv2v_reg  <= w_data_i[21];
      \nz.mem_260_sv2v_reg  <= w_data_i[20];
      \nz.mem_259_sv2v_reg  <= w_data_i[19];
      \nz.mem_258_sv2v_reg  <= w_data_i[18];
      \nz.mem_257_sv2v_reg  <= w_data_i[17];
      \nz.mem_256_sv2v_reg  <= w_data_i[16];
      \nz.mem_255_sv2v_reg  <= w_data_i[15];
      \nz.mem_254_sv2v_reg  <= w_data_i[14];
      \nz.mem_253_sv2v_reg  <= w_data_i[13];
      \nz.mem_252_sv2v_reg  <= w_data_i[12];
      \nz.mem_251_sv2v_reg  <= w_data_i[11];
      \nz.mem_250_sv2v_reg  <= w_data_i[10];
      \nz.mem_249_sv2v_reg  <= w_data_i[9];
      \nz.mem_248_sv2v_reg  <= w_data_i[8];
      \nz.mem_247_sv2v_reg  <= w_data_i[7];
      \nz.mem_246_sv2v_reg  <= w_data_i[6];
      \nz.mem_245_sv2v_reg  <= w_data_i[5];
      \nz.mem_244_sv2v_reg  <= w_data_i[4];
      \nz.mem_243_sv2v_reg  <= w_data_i[3];
      \nz.mem_242_sv2v_reg  <= w_data_i[2];
      \nz.mem_241_sv2v_reg  <= w_data_i[1];
      \nz.mem_240_sv2v_reg  <= w_data_i[0];
    end 
    if(N36) begin
      \nz.mem_239_sv2v_reg  <= w_data_i[79];
      \nz.mem_238_sv2v_reg  <= w_data_i[78];
      \nz.mem_237_sv2v_reg  <= w_data_i[77];
      \nz.mem_236_sv2v_reg  <= w_data_i[76];
      \nz.mem_235_sv2v_reg  <= w_data_i[75];
      \nz.mem_234_sv2v_reg  <= w_data_i[74];
      \nz.mem_233_sv2v_reg  <= w_data_i[73];
      \nz.mem_232_sv2v_reg  <= w_data_i[72];
      \nz.mem_231_sv2v_reg  <= w_data_i[71];
      \nz.mem_230_sv2v_reg  <= w_data_i[70];
      \nz.mem_229_sv2v_reg  <= w_data_i[69];
      \nz.mem_228_sv2v_reg  <= w_data_i[68];
      \nz.mem_227_sv2v_reg  <= w_data_i[67];
      \nz.mem_226_sv2v_reg  <= w_data_i[66];
      \nz.mem_225_sv2v_reg  <= w_data_i[65];
      \nz.mem_224_sv2v_reg  <= w_data_i[64];
      \nz.mem_223_sv2v_reg  <= w_data_i[63];
      \nz.mem_222_sv2v_reg  <= w_data_i[62];
      \nz.mem_221_sv2v_reg  <= w_data_i[61];
      \nz.mem_220_sv2v_reg  <= w_data_i[60];
      \nz.mem_219_sv2v_reg  <= w_data_i[59];
      \nz.mem_218_sv2v_reg  <= w_data_i[58];
      \nz.mem_217_sv2v_reg  <= w_data_i[57];
      \nz.mem_216_sv2v_reg  <= w_data_i[56];
      \nz.mem_215_sv2v_reg  <= w_data_i[55];
      \nz.mem_214_sv2v_reg  <= w_data_i[54];
      \nz.mem_213_sv2v_reg  <= w_data_i[53];
      \nz.mem_212_sv2v_reg  <= w_data_i[52];
      \nz.mem_211_sv2v_reg  <= w_data_i[51];
      \nz.mem_210_sv2v_reg  <= w_data_i[50];
      \nz.mem_209_sv2v_reg  <= w_data_i[49];
      \nz.mem_208_sv2v_reg  <= w_data_i[48];
      \nz.mem_207_sv2v_reg  <= w_data_i[47];
      \nz.mem_206_sv2v_reg  <= w_data_i[46];
      \nz.mem_205_sv2v_reg  <= w_data_i[45];
      \nz.mem_204_sv2v_reg  <= w_data_i[44];
      \nz.mem_203_sv2v_reg  <= w_data_i[43];
      \nz.mem_202_sv2v_reg  <= w_data_i[42];
      \nz.mem_201_sv2v_reg  <= w_data_i[41];
      \nz.mem_200_sv2v_reg  <= w_data_i[40];
      \nz.mem_199_sv2v_reg  <= w_data_i[39];
      \nz.mem_198_sv2v_reg  <= w_data_i[38];
      \nz.mem_197_sv2v_reg  <= w_data_i[37];
      \nz.mem_196_sv2v_reg  <= w_data_i[36];
      \nz.mem_195_sv2v_reg  <= w_data_i[35];
      \nz.mem_194_sv2v_reg  <= w_data_i[34];
      \nz.mem_193_sv2v_reg  <= w_data_i[33];
      \nz.mem_192_sv2v_reg  <= w_data_i[32];
      \nz.mem_191_sv2v_reg  <= w_data_i[31];
      \nz.mem_190_sv2v_reg  <= w_data_i[30];
      \nz.mem_189_sv2v_reg  <= w_data_i[29];
      \nz.mem_188_sv2v_reg  <= w_data_i[28];
      \nz.mem_187_sv2v_reg  <= w_data_i[27];
      \nz.mem_186_sv2v_reg  <= w_data_i[26];
      \nz.mem_185_sv2v_reg  <= w_data_i[25];
      \nz.mem_184_sv2v_reg  <= w_data_i[24];
      \nz.mem_183_sv2v_reg  <= w_data_i[23];
      \nz.mem_182_sv2v_reg  <= w_data_i[22];
      \nz.mem_181_sv2v_reg  <= w_data_i[21];
      \nz.mem_180_sv2v_reg  <= w_data_i[20];
      \nz.mem_179_sv2v_reg  <= w_data_i[19];
      \nz.mem_178_sv2v_reg  <= w_data_i[18];
      \nz.mem_177_sv2v_reg  <= w_data_i[17];
      \nz.mem_176_sv2v_reg  <= w_data_i[16];
      \nz.mem_175_sv2v_reg  <= w_data_i[15];
      \nz.mem_174_sv2v_reg  <= w_data_i[14];
      \nz.mem_173_sv2v_reg  <= w_data_i[13];
      \nz.mem_172_sv2v_reg  <= w_data_i[12];
      \nz.mem_171_sv2v_reg  <= w_data_i[11];
      \nz.mem_170_sv2v_reg  <= w_data_i[10];
      \nz.mem_169_sv2v_reg  <= w_data_i[9];
      \nz.mem_168_sv2v_reg  <= w_data_i[8];
      \nz.mem_167_sv2v_reg  <= w_data_i[7];
      \nz.mem_166_sv2v_reg  <= w_data_i[6];
      \nz.mem_165_sv2v_reg  <= w_data_i[5];
      \nz.mem_164_sv2v_reg  <= w_data_i[4];
      \nz.mem_163_sv2v_reg  <= w_data_i[3];
      \nz.mem_162_sv2v_reg  <= w_data_i[2];
      \nz.mem_161_sv2v_reg  <= w_data_i[1];
      \nz.mem_160_sv2v_reg  <= w_data_i[0];
    end 
    if(N35) begin
      \nz.mem_159_sv2v_reg  <= w_data_i[79];
      \nz.mem_158_sv2v_reg  <= w_data_i[78];
      \nz.mem_157_sv2v_reg  <= w_data_i[77];
      \nz.mem_156_sv2v_reg  <= w_data_i[76];
      \nz.mem_155_sv2v_reg  <= w_data_i[75];
      \nz.mem_154_sv2v_reg  <= w_data_i[74];
      \nz.mem_153_sv2v_reg  <= w_data_i[73];
      \nz.mem_152_sv2v_reg  <= w_data_i[72];
      \nz.mem_151_sv2v_reg  <= w_data_i[71];
      \nz.mem_150_sv2v_reg  <= w_data_i[70];
      \nz.mem_149_sv2v_reg  <= w_data_i[69];
      \nz.mem_148_sv2v_reg  <= w_data_i[68];
      \nz.mem_147_sv2v_reg  <= w_data_i[67];
      \nz.mem_146_sv2v_reg  <= w_data_i[66];
      \nz.mem_145_sv2v_reg  <= w_data_i[65];
      \nz.mem_144_sv2v_reg  <= w_data_i[64];
      \nz.mem_143_sv2v_reg  <= w_data_i[63];
      \nz.mem_142_sv2v_reg  <= w_data_i[62];
      \nz.mem_141_sv2v_reg  <= w_data_i[61];
      \nz.mem_140_sv2v_reg  <= w_data_i[60];
      \nz.mem_139_sv2v_reg  <= w_data_i[59];
      \nz.mem_138_sv2v_reg  <= w_data_i[58];
      \nz.mem_137_sv2v_reg  <= w_data_i[57];
      \nz.mem_136_sv2v_reg  <= w_data_i[56];
      \nz.mem_135_sv2v_reg  <= w_data_i[55];
      \nz.mem_134_sv2v_reg  <= w_data_i[54];
      \nz.mem_133_sv2v_reg  <= w_data_i[53];
      \nz.mem_132_sv2v_reg  <= w_data_i[52];
      \nz.mem_131_sv2v_reg  <= w_data_i[51];
      \nz.mem_130_sv2v_reg  <= w_data_i[50];
      \nz.mem_129_sv2v_reg  <= w_data_i[49];
      \nz.mem_128_sv2v_reg  <= w_data_i[48];
      \nz.mem_127_sv2v_reg  <= w_data_i[47];
      \nz.mem_126_sv2v_reg  <= w_data_i[46];
      \nz.mem_125_sv2v_reg  <= w_data_i[45];
      \nz.mem_124_sv2v_reg  <= w_data_i[44];
      \nz.mem_123_sv2v_reg  <= w_data_i[43];
      \nz.mem_122_sv2v_reg  <= w_data_i[42];
      \nz.mem_121_sv2v_reg  <= w_data_i[41];
      \nz.mem_120_sv2v_reg  <= w_data_i[40];
      \nz.mem_119_sv2v_reg  <= w_data_i[39];
      \nz.mem_118_sv2v_reg  <= w_data_i[38];
      \nz.mem_117_sv2v_reg  <= w_data_i[37];
      \nz.mem_116_sv2v_reg  <= w_data_i[36];
      \nz.mem_115_sv2v_reg  <= w_data_i[35];
      \nz.mem_114_sv2v_reg  <= w_data_i[34];
      \nz.mem_113_sv2v_reg  <= w_data_i[33];
      \nz.mem_112_sv2v_reg  <= w_data_i[32];
      \nz.mem_111_sv2v_reg  <= w_data_i[31];
      \nz.mem_110_sv2v_reg  <= w_data_i[30];
      \nz.mem_109_sv2v_reg  <= w_data_i[29];
      \nz.mem_108_sv2v_reg  <= w_data_i[28];
      \nz.mem_107_sv2v_reg  <= w_data_i[27];
      \nz.mem_106_sv2v_reg  <= w_data_i[26];
      \nz.mem_105_sv2v_reg  <= w_data_i[25];
      \nz.mem_104_sv2v_reg  <= w_data_i[24];
      \nz.mem_103_sv2v_reg  <= w_data_i[23];
      \nz.mem_102_sv2v_reg  <= w_data_i[22];
      \nz.mem_101_sv2v_reg  <= w_data_i[21];
      \nz.mem_100_sv2v_reg  <= w_data_i[20];
      \nz.mem_99_sv2v_reg  <= w_data_i[19];
      \nz.mem_98_sv2v_reg  <= w_data_i[18];
      \nz.mem_97_sv2v_reg  <= w_data_i[17];
      \nz.mem_96_sv2v_reg  <= w_data_i[16];
      \nz.mem_95_sv2v_reg  <= w_data_i[15];
      \nz.mem_94_sv2v_reg  <= w_data_i[14];
      \nz.mem_93_sv2v_reg  <= w_data_i[13];
      \nz.mem_92_sv2v_reg  <= w_data_i[12];
      \nz.mem_91_sv2v_reg  <= w_data_i[11];
      \nz.mem_90_sv2v_reg  <= w_data_i[10];
      \nz.mem_89_sv2v_reg  <= w_data_i[9];
      \nz.mem_88_sv2v_reg  <= w_data_i[8];
      \nz.mem_87_sv2v_reg  <= w_data_i[7];
      \nz.mem_86_sv2v_reg  <= w_data_i[6];
      \nz.mem_85_sv2v_reg  <= w_data_i[5];
      \nz.mem_84_sv2v_reg  <= w_data_i[4];
      \nz.mem_83_sv2v_reg  <= w_data_i[3];
      \nz.mem_82_sv2v_reg  <= w_data_i[2];
      \nz.mem_81_sv2v_reg  <= w_data_i[1];
      \nz.mem_80_sv2v_reg  <= w_data_i[0];
    end 
    if(N34) begin
      \nz.mem_79_sv2v_reg  <= w_data_i[79];
      \nz.mem_78_sv2v_reg  <= w_data_i[78];
      \nz.mem_77_sv2v_reg  <= w_data_i[77];
      \nz.mem_76_sv2v_reg  <= w_data_i[76];
      \nz.mem_75_sv2v_reg  <= w_data_i[75];
      \nz.mem_74_sv2v_reg  <= w_data_i[74];
      \nz.mem_73_sv2v_reg  <= w_data_i[73];
      \nz.mem_72_sv2v_reg  <= w_data_i[72];
      \nz.mem_71_sv2v_reg  <= w_data_i[71];
      \nz.mem_70_sv2v_reg  <= w_data_i[70];
      \nz.mem_69_sv2v_reg  <= w_data_i[69];
      \nz.mem_68_sv2v_reg  <= w_data_i[68];
      \nz.mem_67_sv2v_reg  <= w_data_i[67];
      \nz.mem_66_sv2v_reg  <= w_data_i[66];
      \nz.mem_65_sv2v_reg  <= w_data_i[65];
      \nz.mem_64_sv2v_reg  <= w_data_i[64];
      \nz.mem_63_sv2v_reg  <= w_data_i[63];
      \nz.mem_62_sv2v_reg  <= w_data_i[62];
      \nz.mem_61_sv2v_reg  <= w_data_i[61];
      \nz.mem_60_sv2v_reg  <= w_data_i[60];
      \nz.mem_59_sv2v_reg  <= w_data_i[59];
      \nz.mem_58_sv2v_reg  <= w_data_i[58];
      \nz.mem_57_sv2v_reg  <= w_data_i[57];
      \nz.mem_56_sv2v_reg  <= w_data_i[56];
      \nz.mem_55_sv2v_reg  <= w_data_i[55];
      \nz.mem_54_sv2v_reg  <= w_data_i[54];
      \nz.mem_53_sv2v_reg  <= w_data_i[53];
      \nz.mem_52_sv2v_reg  <= w_data_i[52];
      \nz.mem_51_sv2v_reg  <= w_data_i[51];
      \nz.mem_50_sv2v_reg  <= w_data_i[50];
      \nz.mem_49_sv2v_reg  <= w_data_i[49];
      \nz.mem_48_sv2v_reg  <= w_data_i[48];
      \nz.mem_47_sv2v_reg  <= w_data_i[47];
      \nz.mem_46_sv2v_reg  <= w_data_i[46];
      \nz.mem_45_sv2v_reg  <= w_data_i[45];
      \nz.mem_44_sv2v_reg  <= w_data_i[44];
      \nz.mem_43_sv2v_reg  <= w_data_i[43];
      \nz.mem_42_sv2v_reg  <= w_data_i[42];
      \nz.mem_41_sv2v_reg  <= w_data_i[41];
      \nz.mem_40_sv2v_reg  <= w_data_i[40];
      \nz.mem_39_sv2v_reg  <= w_data_i[39];
      \nz.mem_38_sv2v_reg  <= w_data_i[38];
      \nz.mem_37_sv2v_reg  <= w_data_i[37];
      \nz.mem_36_sv2v_reg  <= w_data_i[36];
      \nz.mem_35_sv2v_reg  <= w_data_i[35];
      \nz.mem_34_sv2v_reg  <= w_data_i[34];
      \nz.mem_33_sv2v_reg  <= w_data_i[33];
      \nz.mem_32_sv2v_reg  <= w_data_i[32];
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_00000050_00000008
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [2:0] w_addr_i;
  input [79:0] w_data_i;
  input [2:0] r_addr_i;
  output [79:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [79:0] r_data_o;

  bsg_mem_1r1w_synth_00000050_00000008_0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bp_be_expander
(
  cinstr_i,
  instr_o
);

  input [15:0] cinstr_i;
  output [31:0] instr_o;
  wire [31:0] instr_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511;
  wire [4:3] rs1,rs2;
  wire [4:0] rd;
  wire [63:0] imm;
  assign N9 = cinstr_i[1] & N209;
  assign N10 = N212 & cinstr_i[0];
  assign N11 = N210 & N191;
  assign N12 = N11 & cinstr_i[0];
  assign N13 = N190 & N211;
  assign N14 = N13 & cinstr_i[0];
  assign N16 = cinstr_i[1] | N209;
  assign N18 = N198 & N209;
  assign N20 = N210 & N185;
  assign N21 = N20 & N209;
  assign N23 = N40 & N182;
  assign N24 = N23 & N209;
  assign N25 = N140 & N185;
  assign N26 = N25 & N209;
  assign N27 = N40 & N185;
  assign N28 = N27 & N209;
  assign N30 = N13 & N209;
  assign N31 = N41 & N209;
  assign N33 = N11 & N209;
  assign N34 = N192 & N209;
  assign N35 = N38 & N209;
  assign N36 = N43 & N209;
  assign N38 = N140 & N191;
  assign N39 = N38 & cinstr_i[0];
  assign N40 = cinstr_i[15] & cinstr_i[14];
  assign N41 = N40 & N211;
  assign N42 = N41 & cinstr_i[0];
  assign N43 = N40 & N191;
  assign N44 = N43 & cinstr_i[0];
  assign N46 = cinstr_i[15] | cinstr_i[14];
  assign N47 = cinstr_i[13] | cinstr_i[12];
  assign N48 = cinstr_i[11] | cinstr_i[10];
  assign N49 = cinstr_i[9] | cinstr_i[8];
  assign N50 = cinstr_i[7] | cinstr_i[6];
  assign N51 = cinstr_i[5] | cinstr_i[4];
  assign N52 = cinstr_i[3] | cinstr_i[2];
  assign N53 = N46 | N47;
  assign N54 = N48 | N49;
  assign N55 = N50 | N51;
  assign N56 = N52 | N16;
  assign N57 = N53 | N54;
  assign N58 = N55 | N56;
  assign N59 = N57 | N58;
  assign N60 = N74 & N65;
  assign N62 = N210 & N182;
  assign N63 = N62 & N209;
  assign N64 = N195 & N198;
  assign N65 = N64 & cinstr_i[0];
  assign N66 = N70 & N65;
  assign N68 = N208 & N194;
  assign N69 = cinstr_i[10] & N198;
  assign N70 = N140 & N68;
  assign N71 = N69 & cinstr_i[0];
  assign N72 = N70 & N71;
  assign N73 = N208 & cinstr_i[11];
  assign N74 = N140 & N73;
  assign N75 = N74 & cinstr_i[10];
  assign N76 = N208 & N209;
  assign N77 = N140 & N76;
  assign N80 = N194 & N195;
  assign N81 = N196 & N79;
  assign N82 = N197 & N133;
  assign N83 = N134 & N103;
  assign N84 = N104 & N105;
  assign N85 = N210 & N125;
  assign N86 = N80 & N81;
  assign N87 = N82 & N83;
  assign N88 = N84 & N18;
  assign N89 = N85 & N86;
  assign N90 = N87 & N88;
  assign N91 = N89 & N90;
  assign N92 = N189 | cinstr_i[14];
  assign N93 = cinstr_i[13] | N124;
  assign N94 = N198 | cinstr_i[0];
  assign N95 = N92 | N93;
  assign N96 = N52 | N94;
  assign N97 = N95 | N54;
  assign N98 = N55 | N96;
  assign N99 = N97 | N98;
  assign N101 = N126 & N108;
  assign N102 = N101 & N109;
  assign N106 = N103 & N104;
  assign N107 = N105 & cinstr_i[1];
  assign N108 = N135 & N106;
  assign N109 = N107 & N209;
  assign N110 = N144 & N108;
  assign N111 = N110 & N109;
  assign N112 = N126 & N9;
  assign N113 = N144 & N9;
  assign N114 = cinstr_i[6] & cinstr_i[5];
  assign N115 = N142 & N114;
  assign N116 = N126 & N115;
  assign N117 = N116 & N202;
  assign N118 = cinstr_i[6] & N134;
  assign N119 = N142 & N118;
  assign N120 = N126 & N119;
  assign N121 = N120 & N202;
  assign N122 = N126 & N130;
  assign N123 = N122 & N202;
  assign N125 = N208 & N124;
  assign N126 = N140 & N125;
  assign N127 = N126 & N136;
  assign N128 = N127 & N202;
  assign N129 = N133 & cinstr_i[5];
  assign N130 = N142 & N129;
  assign N131 = N144 & N130;
  assign N132 = N131 & N202;
  assign N135 = N133 & N134;
  assign N136 = N142 & N135;
  assign N137 = N144 & N136;
  assign N138 = N137 & N202;
  assign N139 = cinstr_i[1] & cinstr_i[0];
  assign N140 = cinstr_i[15] & N207;
  assign N141 = N208 & cinstr_i[12];
  assign N142 = cinstr_i[11] & cinstr_i[10];
  assign N143 = cinstr_i[6] & cinstr_i[0];
  assign N144 = N140 & N141;
  assign N145 = N142 & N143;
  assign N146 = N144 & N145;
  assign N147 = N140 & N211;
  assign N148 = N147 & N209;
  assign N182 = N208 & cinstr_i[1];
  assign N183 = N190 & N182;
  assign N184 = N183 & N209;
  assign N185 = cinstr_i[13] & cinstr_i[1];
  assign N186 = N190 & N185;
  assign N187 = N186 & N209;
  assign N190 = N189 & cinstr_i[14];
  assign N191 = cinstr_i[13] & N198;
  assign N192 = N190 & N191;
  assign N193 = N192 & cinstr_i[0];
  assign N199 = cinstr_i[13] & N194;
  assign N200 = N195 & N196;
  assign N201 = cinstr_i[8] & N197;
  assign N202 = N198 & cinstr_i[0];
  assign N203 = N190 & N199;
  assign N204 = N200 & N201;
  assign N205 = N203 & N204;
  assign N206 = N205 & N202;
  assign N210 = N189 & N207;
  assign N211 = N208 & N198;
  assign N212 = N210 & N211;
  assign N213 = N212 & N209;
  assign rs1 = (N0)? cinstr_i[11:10] : 
               (N284)? { 1'b0, 1'b1 } : 
               (N286)? { 1'b0, 1'b1 } : 1'b0;
  assign N0 = N15;
  assign rs2 = (N0)? cinstr_i[6:5] : 
               (N284)? { 1'b0, 1'b1 } : 
               (N286)? { 1'b0, 1'b1 } : 1'b0;
  assign rd = (N0)? cinstr_i[11:7] : 
              (N284)? { 1'b0, 1'b1, cinstr_i[9:7] } : 
              (N286)? { 1'b0, 1'b1, cinstr_i[4:2] } : 1'b0;
  assign imm = (N1)? { cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[4:3], cinstr_i[5:5], cinstr_i[2:2], cinstr_i[6:6], 1'b0, 1'b0, 1'b0, 1'b0 } : 
               (N288)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[10:7], cinstr_i[12:11], cinstr_i[5:5], cinstr_i[6:6], 1'b0, 1'b0 } : 
               (N291)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[3:2], cinstr_i[12:12], cinstr_i[6:4], 1'b0, 1'b0 } : 
               (N294)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[4:2], cinstr_i[12:12], cinstr_i[6:5], 1'b0, 1'b0, 1'b0 } : 
               (N297)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[8:7], cinstr_i[12:9], 1'b0, 1'b0 } : 
               (N300)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[9:7], cinstr_i[12:10], 1'b0, 1'b0, 1'b0 } : 
               (N303)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[5:5], cinstr_i[12:10], cinstr_i[6:6], 1'b0, 1'b0 } : 
               (N306)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[6:5], cinstr_i[12:10], 1'b0, 1'b0, 1'b0 } : 
               (N309)? { cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[8:8], cinstr_i[10:9], cinstr_i[6:6], cinstr_i[7:7], cinstr_i[2:2], cinstr_i[11:11], cinstr_i[5:3], 1'b0 } : 
               (N312)? { cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[6:5], cinstr_i[2:2], cinstr_i[11:10], cinstr_i[4:3], 1'b0 } : 
               (N315)? { cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[6:2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
               (N318)? { cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[6:2] } : 
               (N321)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[12:12], cinstr_i[6:2] } : 
               (N324)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[12:12], cinstr_i[6:2] } : 
               (N327)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = N206;
  assign { N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150 } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N329)? { imm[11:0], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N331)? { imm[11:0], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N333)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N335)? { imm[11:0], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, rd, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N337)? { imm[11:0], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, rd, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N340)? { imm[11:5], rs2, cinstr_i[4:2], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, imm[4:0], 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N342)? { imm[11:5], rs2, cinstr_i[4:2], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, imm[4:0], 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N345)? { imm[11:0], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, rd, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N348)? { imm[11:5], rs2, cinstr_i[4:2], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, imm[4:0], 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N351)? { imm[11:0], rs1, cinstr_i[9:7], 1'b0, 1'b1, 1'b0, rd, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N354)? { imm[11:0], rs1, cinstr_i[9:7], 1'b0, 1'b1, 1'b1, rd, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N357)? { imm[11:5], rs2, cinstr_i[4:2], rs1, cinstr_i[9:7], 1'b0, 1'b1, 1'b0, imm[4:0], 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N360)? { imm[11:5], rs2, cinstr_i[4:2], rs1, cinstr_i[9:7], 1'b0, 1'b1, 1'b1, imm[4:0], 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N363)? { imm[11:0], rs1, cinstr_i[9:7], 1'b0, 1'b1, 1'b1, rd, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N366)? { imm[11:5], rs2, cinstr_i[4:2], rs1, cinstr_i[9:7], 1'b0, 1'b1, 1'b1, imm[4:0], 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N369)? { imm[20:20], imm[10:1], imm[11:11], imm[19:12], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N371)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs1, cinstr_i[9:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N374)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs1, cinstr_i[9:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N377)? { imm[12:12], imm[10:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs1, cinstr_i[9:7], 1'b0, 1'b0, 1'b0, imm[4:1], imm[11:11], 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N380)? { imm[12:12], imm[10:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs1, cinstr_i[9:7], 1'b0, 1'b0, 1'b1, imm[4:1], imm[11:11], 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N383)? { imm[11:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N386)? { imm[31:12], rd, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N388)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N390)? { imm[11:0], rd, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N393)? { imm[11:0], rd, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N396)? { imm[11:0], rd, 1'b0, 1'b0, 1'b1, rd, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N399)? { imm[11:0], rd, 1'b1, 1'b0, 1'b1, rd, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N402)? { imm[11:0], rd, 1'b1, 1'b0, 1'b1, rd, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N404)? { imm[11:0], rd, 1'b1, 1'b1, 1'b1, rd, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N407)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs2, cinstr_i[4:2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N410)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs2, cinstr_i[4:2], rd, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N413)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs2, cinstr_i[4:2], rd, 1'b1, 1'b1, 1'b1, rd, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N416)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs2, cinstr_i[4:2], rd, 1'b1, 1'b1, 1'b0, rd, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N419)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs2, cinstr_i[4:2], rd, 1'b1, 1'b0, 1'b0, rd, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N422)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs2, cinstr_i[4:2], rd, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N425)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs2, cinstr_i[4:2], rd, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N428)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs2, cinstr_i[4:2], rd, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N431)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i } : 1'b0;
  assign N2 = N91;
  assign { N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218 } = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N4)? { N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150 } : 1'b0;
  assign N3 = N217;
  assign N4 = N448;
  assign { N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N6)? { N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150 } : 1'b0;
  assign N5 = N250;
  assign N6 = N511;
  assign instr_o = (N7)? { N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218 } : 
                   (N8)? { N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251 } : 
                   (N216)? { N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150 } : 1'b0;
  assign N7 = N188;
  assign N8 = N214;
  assign N15 = N435 | N193;
  assign N435 = N434 | N206;
  assign N434 = N433 | N14;
  assign N433 = N432 | N12;
  assign N432 = N9 | N10;
  assign N17 = ~N16;
  assign N19 = N139 | N18;
  assign N22 = N21 | N187;
  assign N29 = N26 | N28;
  assign N32 = N30 | N31;
  assign N37 = N437 | N36;
  assign N437 = N436 | N35;
  assign N436 = N33 | N34;
  assign N45 = N42 | N44;
  assign N61 = N441 | N60;
  assign N441 = N440 | N14;
  assign N440 = N439 | N12;
  assign N439 = N438 | N10;
  assign N438 = ~N59;
  assign N67 = N63 | N66;
  assign N78 = N139 | N442;
  assign N442 = N75 | N77;
  assign N79 = ~cinstr_i[8];
  assign N100 = ~N99;
  assign N103 = ~cinstr_i[4];
  assign N104 = ~cinstr_i[3];
  assign N105 = ~cinstr_i[2];
  assign N124 = ~cinstr_i[12];
  assign N133 = ~cinstr_i[6];
  assign N134 = ~cinstr_i[5];
  assign N149 = N139 | N443;
  assign N443 = N146 | N148;
  assign N188 = N184 | N187;
  assign N189 = ~cinstr_i[15];
  assign N194 = ~cinstr_i[11];
  assign N195 = ~cinstr_i[10];
  assign N196 = ~cinstr_i[9];
  assign N197 = ~cinstr_i[7];
  assign N198 = ~cinstr_i[1];
  assign N207 = ~cinstr_i[14];
  assign N208 = ~cinstr_i[13];
  assign N209 = ~cinstr_i[0];
  assign N214 = N444 | N213;
  assign N444 = N193 | N206;
  assign N215 = N214 | N188;
  assign N216 = ~N215;
  assign N217 = ~N448;
  assign N448 = N447 | cinstr_i[7];
  assign N447 = N446 | cinstr_i[8];
  assign N446 = N445 | cinstr_i[9];
  assign N445 = cinstr_i[11] | cinstr_i[10];
  assign N250 = ~N511;
  assign N511 = N510 | imm[0];
  assign N510 = N509 | imm[1];
  assign N509 = N508 | imm[2];
  assign N508 = N507 | imm[3];
  assign N507 = N506 | imm[4];
  assign N506 = N505 | imm[5];
  assign N505 = N504 | imm[6];
  assign N504 = N503 | imm[7];
  assign N503 = N502 | imm[8];
  assign N502 = N501 | imm[9];
  assign N501 = N500 | imm[10];
  assign N500 = N499 | imm[11];
  assign N499 = N498 | imm[12];
  assign N498 = N497 | imm[13];
  assign N497 = N496 | imm[14];
  assign N496 = N495 | imm[15];
  assign N495 = N494 | imm[16];
  assign N494 = N493 | imm[17];
  assign N493 = N492 | imm[18];
  assign N492 = N491 | imm[19];
  assign N491 = N490 | imm[20];
  assign N490 = N489 | imm[21];
  assign N489 = N488 | imm[22];
  assign N488 = N487 | imm[23];
  assign N487 = N486 | imm[24];
  assign N486 = N485 | imm[25];
  assign N485 = N484 | imm[26];
  assign N484 = N483 | imm[27];
  assign N483 = N482 | imm[28];
  assign N482 = N481 | imm[29];
  assign N481 = N480 | imm[30];
  assign N480 = N479 | imm[31];
  assign N479 = N478 | imm[32];
  assign N478 = N477 | imm[33];
  assign N477 = N476 | imm[34];
  assign N476 = N475 | imm[35];
  assign N475 = N474 | imm[36];
  assign N474 = N473 | imm[37];
  assign N473 = N472 | imm[38];
  assign N472 = N471 | imm[39];
  assign N471 = N470 | imm[40];
  assign N470 = N469 | imm[41];
  assign N469 = N468 | imm[42];
  assign N468 = N467 | imm[43];
  assign N467 = N466 | imm[44];
  assign N466 = N465 | imm[45];
  assign N465 = N464 | imm[46];
  assign N464 = N463 | imm[47];
  assign N463 = N462 | imm[48];
  assign N462 = N461 | imm[49];
  assign N461 = N460 | imm[50];
  assign N460 = N459 | imm[51];
  assign N459 = N458 | imm[52];
  assign N458 = N457 | imm[53];
  assign N457 = N456 | imm[54];
  assign N456 = N455 | imm[55];
  assign N455 = N454 | imm[56];
  assign N454 = N453 | imm[57];
  assign N453 = N452 | imm[58];
  assign N452 = N451 | imm[59];
  assign N451 = N450 | imm[60];
  assign N450 = N449 | imm[61];
  assign N449 = imm[63] | imm[62];
  assign N283 = ~N15;
  assign N284 = N17 & N283;
  assign N285 = N283 & N16;
  assign N286 = N19 & N285;
  assign N287 = ~N206;
  assign N288 = N213 & N287;
  assign N289 = ~N213;
  assign N290 = N287 & N289;
  assign N291 = N184 & N290;
  assign N292 = ~N184;
  assign N293 = N290 & N292;
  assign N294 = N22 & N293;
  assign N295 = ~N22;
  assign N296 = N293 & N295;
  assign N297 = N24 & N296;
  assign N298 = ~N24;
  assign N299 = N296 & N298;
  assign N300 = N29 & N299;
  assign N301 = ~N29;
  assign N302 = N299 & N301;
  assign N303 = N32 & N302;
  assign N304 = ~N32;
  assign N305 = N302 & N304;
  assign N306 = N37 & N305;
  assign N307 = ~N37;
  assign N308 = N305 & N307;
  assign N309 = N39 & N308;
  assign N310 = ~N39;
  assign N311 = N308 & N310;
  assign N312 = N45 & N311;
  assign N313 = ~N45;
  assign N314 = N311 & N313;
  assign N315 = N193 & N314;
  assign N316 = ~N193;
  assign N317 = N314 & N316;
  assign N318 = N61 & N317;
  assign N319 = ~N61;
  assign N320 = N317 & N319;
  assign N321 = N67 & N320;
  assign N322 = ~N67;
  assign N323 = N320 & N322;
  assign N324 = N72 & N323;
  assign N325 = ~N72;
  assign N326 = N323 & N325;
  assign N327 = N78 & N326;
  assign N328 = ~N91;
  assign N329 = N213 & N328;
  assign N330 = N328 & N289;
  assign N331 = N206 & N330;
  assign N332 = N330 & N287;
  assign N333 = N100 & N332;
  assign N334 = N332 & N99;
  assign N335 = N184 & N334;
  assign N336 = N334 & N292;
  assign N337 = N187 & N336;
  assign N338 = ~N187;
  assign N339 = N336 & N338;
  assign N340 = N24 & N339;
  assign N341 = N339 & N298;
  assign N342 = N28 & N341;
  assign N343 = ~N28;
  assign N344 = N341 & N343;
  assign N345 = N21 & N344;
  assign N346 = ~N21;
  assign N347 = N344 & N346;
  assign N348 = N26 & N347;
  assign N349 = ~N26;
  assign N350 = N347 & N349;
  assign N351 = N30 & N350;
  assign N352 = ~N30;
  assign N353 = N350 & N352;
  assign N354 = N34 & N353;
  assign N355 = ~N34;
  assign N356 = N353 & N355;
  assign N357 = N31 & N356;
  assign N358 = ~N31;
  assign N359 = N356 & N358;
  assign N360 = N36 & N359;
  assign N361 = ~N36;
  assign N362 = N359 & N361;
  assign N363 = N33 & N362;
  assign N364 = ~N33;
  assign N365 = N362 & N364;
  assign N366 = N35 & N365;
  assign N367 = ~N35;
  assign N368 = N365 & N367;
  assign N369 = N39 & N368;
  assign N370 = N368 & N310;
  assign N371 = N102 & N370;
  assign N372 = ~N102;
  assign N373 = N370 & N372;
  assign N374 = N111 & N373;
  assign N375 = ~N111;
  assign N376 = N373 & N375;
  assign N377 = N42 & N376;
  assign N378 = ~N42;
  assign N379 = N376 & N378;
  assign N380 = N44 & N379;
  assign N381 = ~N44;
  assign N382 = N379 & N381;
  assign N383 = N14 & N382;
  assign N384 = ~N14;
  assign N385 = N382 & N384;
  assign N386 = N193 & N385;
  assign N387 = N385 & N316;
  assign N388 = N438 & N387;
  assign N389 = N387 & N59;
  assign N390 = N10 & N389;
  assign N391 = ~N10;
  assign N392 = N389 & N391;
  assign N393 = N12 & N392;
  assign N394 = ~N12;
  assign N395 = N392 & N394;
  assign N396 = N63 & N395;
  assign N397 = ~N63;
  assign N398 = N395 & N397;
  assign N399 = N66 & N398;
  assign N400 = ~N66;
  assign N401 = N398 & N400;
  assign N402 = N72 & N401;
  assign N403 = N401 & N325;
  assign N404 = N60 & N403;
  assign N405 = ~N60;
  assign N406 = N403 & N405;
  assign N407 = N112 & N406;
  assign N408 = ~N112;
  assign N409 = N406 & N408;
  assign N410 = N113 & N409;
  assign N411 = ~N113;
  assign N412 = N409 & N411;
  assign N413 = N117 & N412;
  assign N414 = ~N117;
  assign N415 = N412 & N414;
  assign N416 = N121 & N415;
  assign N417 = ~N121;
  assign N418 = N415 & N417;
  assign N419 = N123 & N418;
  assign N420 = ~N123;
  assign N421 = N418 & N420;
  assign N422 = N128 & N421;
  assign N423 = ~N128;
  assign N424 = N421 & N423;
  assign N425 = N132 & N424;
  assign N426 = ~N132;
  assign N427 = N424 & N426;
  assign N428 = N138 & N427;
  assign N429 = ~N138;
  assign N430 = N427 & N429;
  assign N431 = N149 & N430;

endmodule



module bsg_dff_reset_en_width_p39
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [38:0] data_i;
  output [38:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [38:0] data_o;
  wire N0,N1,N2;
  reg data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,
  data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,
  data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,
  data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,
  data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,
  data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_synth_000000ae_00000008_0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [2:0] w_addr_i;
  input [173:0] w_data_i;
  input [2:0] r_addr_i;
  output [173:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [173:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53;
  wire [1391:0] \nz.mem ;
  reg \nz.mem_1391_sv2v_reg ,\nz.mem_1390_sv2v_reg ,\nz.mem_1389_sv2v_reg ,
  \nz.mem_1388_sv2v_reg ,\nz.mem_1387_sv2v_reg ,\nz.mem_1386_sv2v_reg ,
  \nz.mem_1385_sv2v_reg ,\nz.mem_1384_sv2v_reg ,\nz.mem_1383_sv2v_reg ,\nz.mem_1382_sv2v_reg ,
  \nz.mem_1381_sv2v_reg ,\nz.mem_1380_sv2v_reg ,\nz.mem_1379_sv2v_reg ,
  \nz.mem_1378_sv2v_reg ,\nz.mem_1377_sv2v_reg ,\nz.mem_1376_sv2v_reg ,\nz.mem_1375_sv2v_reg ,
  \nz.mem_1374_sv2v_reg ,\nz.mem_1373_sv2v_reg ,\nz.mem_1372_sv2v_reg ,
  \nz.mem_1371_sv2v_reg ,\nz.mem_1370_sv2v_reg ,\nz.mem_1369_sv2v_reg ,\nz.mem_1368_sv2v_reg ,
  \nz.mem_1367_sv2v_reg ,\nz.mem_1366_sv2v_reg ,\nz.mem_1365_sv2v_reg ,
  \nz.mem_1364_sv2v_reg ,\nz.mem_1363_sv2v_reg ,\nz.mem_1362_sv2v_reg ,\nz.mem_1361_sv2v_reg ,
  \nz.mem_1360_sv2v_reg ,\nz.mem_1359_sv2v_reg ,\nz.mem_1358_sv2v_reg ,
  \nz.mem_1357_sv2v_reg ,\nz.mem_1356_sv2v_reg ,\nz.mem_1355_sv2v_reg ,\nz.mem_1354_sv2v_reg ,
  \nz.mem_1353_sv2v_reg ,\nz.mem_1352_sv2v_reg ,\nz.mem_1351_sv2v_reg ,
  \nz.mem_1350_sv2v_reg ,\nz.mem_1349_sv2v_reg ,\nz.mem_1348_sv2v_reg ,\nz.mem_1347_sv2v_reg ,
  \nz.mem_1346_sv2v_reg ,\nz.mem_1345_sv2v_reg ,\nz.mem_1344_sv2v_reg ,
  \nz.mem_1343_sv2v_reg ,\nz.mem_1342_sv2v_reg ,\nz.mem_1341_sv2v_reg ,\nz.mem_1340_sv2v_reg ,
  \nz.mem_1339_sv2v_reg ,\nz.mem_1338_sv2v_reg ,\nz.mem_1337_sv2v_reg ,
  \nz.mem_1336_sv2v_reg ,\nz.mem_1335_sv2v_reg ,\nz.mem_1334_sv2v_reg ,\nz.mem_1333_sv2v_reg ,
  \nz.mem_1332_sv2v_reg ,\nz.mem_1331_sv2v_reg ,\nz.mem_1330_sv2v_reg ,
  \nz.mem_1329_sv2v_reg ,\nz.mem_1328_sv2v_reg ,\nz.mem_1327_sv2v_reg ,\nz.mem_1326_sv2v_reg ,
  \nz.mem_1325_sv2v_reg ,\nz.mem_1324_sv2v_reg ,\nz.mem_1323_sv2v_reg ,
  \nz.mem_1322_sv2v_reg ,\nz.mem_1321_sv2v_reg ,\nz.mem_1320_sv2v_reg ,\nz.mem_1319_sv2v_reg ,
  \nz.mem_1318_sv2v_reg ,\nz.mem_1317_sv2v_reg ,\nz.mem_1316_sv2v_reg ,
  \nz.mem_1315_sv2v_reg ,\nz.mem_1314_sv2v_reg ,\nz.mem_1313_sv2v_reg ,\nz.mem_1312_sv2v_reg ,
  \nz.mem_1311_sv2v_reg ,\nz.mem_1310_sv2v_reg ,\nz.mem_1309_sv2v_reg ,
  \nz.mem_1308_sv2v_reg ,\nz.mem_1307_sv2v_reg ,\nz.mem_1306_sv2v_reg ,
  \nz.mem_1305_sv2v_reg ,\nz.mem_1304_sv2v_reg ,\nz.mem_1303_sv2v_reg ,\nz.mem_1302_sv2v_reg ,
  \nz.mem_1301_sv2v_reg ,\nz.mem_1300_sv2v_reg ,\nz.mem_1299_sv2v_reg ,
  \nz.mem_1298_sv2v_reg ,\nz.mem_1297_sv2v_reg ,\nz.mem_1296_sv2v_reg ,\nz.mem_1295_sv2v_reg ,
  \nz.mem_1294_sv2v_reg ,\nz.mem_1293_sv2v_reg ,\nz.mem_1292_sv2v_reg ,
  \nz.mem_1291_sv2v_reg ,\nz.mem_1290_sv2v_reg ,\nz.mem_1289_sv2v_reg ,\nz.mem_1288_sv2v_reg ,
  \nz.mem_1287_sv2v_reg ,\nz.mem_1286_sv2v_reg ,\nz.mem_1285_sv2v_reg ,
  \nz.mem_1284_sv2v_reg ,\nz.mem_1283_sv2v_reg ,\nz.mem_1282_sv2v_reg ,\nz.mem_1281_sv2v_reg ,
  \nz.mem_1280_sv2v_reg ,\nz.mem_1279_sv2v_reg ,\nz.mem_1278_sv2v_reg ,
  \nz.mem_1277_sv2v_reg ,\nz.mem_1276_sv2v_reg ,\nz.mem_1275_sv2v_reg ,\nz.mem_1274_sv2v_reg ,
  \nz.mem_1273_sv2v_reg ,\nz.mem_1272_sv2v_reg ,\nz.mem_1271_sv2v_reg ,
  \nz.mem_1270_sv2v_reg ,\nz.mem_1269_sv2v_reg ,\nz.mem_1268_sv2v_reg ,\nz.mem_1267_sv2v_reg ,
  \nz.mem_1266_sv2v_reg ,\nz.mem_1265_sv2v_reg ,\nz.mem_1264_sv2v_reg ,
  \nz.mem_1263_sv2v_reg ,\nz.mem_1262_sv2v_reg ,\nz.mem_1261_sv2v_reg ,\nz.mem_1260_sv2v_reg ,
  \nz.mem_1259_sv2v_reg ,\nz.mem_1258_sv2v_reg ,\nz.mem_1257_sv2v_reg ,
  \nz.mem_1256_sv2v_reg ,\nz.mem_1255_sv2v_reg ,\nz.mem_1254_sv2v_reg ,\nz.mem_1253_sv2v_reg ,
  \nz.mem_1252_sv2v_reg ,\nz.mem_1251_sv2v_reg ,\nz.mem_1250_sv2v_reg ,
  \nz.mem_1249_sv2v_reg ,\nz.mem_1248_sv2v_reg ,\nz.mem_1247_sv2v_reg ,\nz.mem_1246_sv2v_reg ,
  \nz.mem_1245_sv2v_reg ,\nz.mem_1244_sv2v_reg ,\nz.mem_1243_sv2v_reg ,
  \nz.mem_1242_sv2v_reg ,\nz.mem_1241_sv2v_reg ,\nz.mem_1240_sv2v_reg ,\nz.mem_1239_sv2v_reg ,
  \nz.mem_1238_sv2v_reg ,\nz.mem_1237_sv2v_reg ,\nz.mem_1236_sv2v_reg ,
  \nz.mem_1235_sv2v_reg ,\nz.mem_1234_sv2v_reg ,\nz.mem_1233_sv2v_reg ,\nz.mem_1232_sv2v_reg ,
  \nz.mem_1231_sv2v_reg ,\nz.mem_1230_sv2v_reg ,\nz.mem_1229_sv2v_reg ,
  \nz.mem_1228_sv2v_reg ,\nz.mem_1227_sv2v_reg ,\nz.mem_1226_sv2v_reg ,
  \nz.mem_1225_sv2v_reg ,\nz.mem_1224_sv2v_reg ,\nz.mem_1223_sv2v_reg ,\nz.mem_1222_sv2v_reg ,
  \nz.mem_1221_sv2v_reg ,\nz.mem_1220_sv2v_reg ,\nz.mem_1219_sv2v_reg ,
  \nz.mem_1218_sv2v_reg ,\nz.mem_1217_sv2v_reg ,\nz.mem_1216_sv2v_reg ,\nz.mem_1215_sv2v_reg ,
  \nz.mem_1214_sv2v_reg ,\nz.mem_1213_sv2v_reg ,\nz.mem_1212_sv2v_reg ,
  \nz.mem_1211_sv2v_reg ,\nz.mem_1210_sv2v_reg ,\nz.mem_1209_sv2v_reg ,\nz.mem_1208_sv2v_reg ,
  \nz.mem_1207_sv2v_reg ,\nz.mem_1206_sv2v_reg ,\nz.mem_1205_sv2v_reg ,
  \nz.mem_1204_sv2v_reg ,\nz.mem_1203_sv2v_reg ,\nz.mem_1202_sv2v_reg ,\nz.mem_1201_sv2v_reg ,
  \nz.mem_1200_sv2v_reg ,\nz.mem_1199_sv2v_reg ,\nz.mem_1198_sv2v_reg ,
  \nz.mem_1197_sv2v_reg ,\nz.mem_1196_sv2v_reg ,\nz.mem_1195_sv2v_reg ,\nz.mem_1194_sv2v_reg ,
  \nz.mem_1193_sv2v_reg ,\nz.mem_1192_sv2v_reg ,\nz.mem_1191_sv2v_reg ,
  \nz.mem_1190_sv2v_reg ,\nz.mem_1189_sv2v_reg ,\nz.mem_1188_sv2v_reg ,\nz.mem_1187_sv2v_reg ,
  \nz.mem_1186_sv2v_reg ,\nz.mem_1185_sv2v_reg ,\nz.mem_1184_sv2v_reg ,
  \nz.mem_1183_sv2v_reg ,\nz.mem_1182_sv2v_reg ,\nz.mem_1181_sv2v_reg ,\nz.mem_1180_sv2v_reg ,
  \nz.mem_1179_sv2v_reg ,\nz.mem_1178_sv2v_reg ,\nz.mem_1177_sv2v_reg ,
  \nz.mem_1176_sv2v_reg ,\nz.mem_1175_sv2v_reg ,\nz.mem_1174_sv2v_reg ,\nz.mem_1173_sv2v_reg ,
  \nz.mem_1172_sv2v_reg ,\nz.mem_1171_sv2v_reg ,\nz.mem_1170_sv2v_reg ,
  \nz.mem_1169_sv2v_reg ,\nz.mem_1168_sv2v_reg ,\nz.mem_1167_sv2v_reg ,\nz.mem_1166_sv2v_reg ,
  \nz.mem_1165_sv2v_reg ,\nz.mem_1164_sv2v_reg ,\nz.mem_1163_sv2v_reg ,
  \nz.mem_1162_sv2v_reg ,\nz.mem_1161_sv2v_reg ,\nz.mem_1160_sv2v_reg ,\nz.mem_1159_sv2v_reg ,
  \nz.mem_1158_sv2v_reg ,\nz.mem_1157_sv2v_reg ,\nz.mem_1156_sv2v_reg ,
  \nz.mem_1155_sv2v_reg ,\nz.mem_1154_sv2v_reg ,\nz.mem_1153_sv2v_reg ,\nz.mem_1152_sv2v_reg ,
  \nz.mem_1151_sv2v_reg ,\nz.mem_1150_sv2v_reg ,\nz.mem_1149_sv2v_reg ,
  \nz.mem_1148_sv2v_reg ,\nz.mem_1147_sv2v_reg ,\nz.mem_1146_sv2v_reg ,
  \nz.mem_1145_sv2v_reg ,\nz.mem_1144_sv2v_reg ,\nz.mem_1143_sv2v_reg ,\nz.mem_1142_sv2v_reg ,
  \nz.mem_1141_sv2v_reg ,\nz.mem_1140_sv2v_reg ,\nz.mem_1139_sv2v_reg ,
  \nz.mem_1138_sv2v_reg ,\nz.mem_1137_sv2v_reg ,\nz.mem_1136_sv2v_reg ,\nz.mem_1135_sv2v_reg ,
  \nz.mem_1134_sv2v_reg ,\nz.mem_1133_sv2v_reg ,\nz.mem_1132_sv2v_reg ,
  \nz.mem_1131_sv2v_reg ,\nz.mem_1130_sv2v_reg ,\nz.mem_1129_sv2v_reg ,\nz.mem_1128_sv2v_reg ,
  \nz.mem_1127_sv2v_reg ,\nz.mem_1126_sv2v_reg ,\nz.mem_1125_sv2v_reg ,
  \nz.mem_1124_sv2v_reg ,\nz.mem_1123_sv2v_reg ,\nz.mem_1122_sv2v_reg ,\nz.mem_1121_sv2v_reg ,
  \nz.mem_1120_sv2v_reg ,\nz.mem_1119_sv2v_reg ,\nz.mem_1118_sv2v_reg ,
  \nz.mem_1117_sv2v_reg ,\nz.mem_1116_sv2v_reg ,\nz.mem_1115_sv2v_reg ,\nz.mem_1114_sv2v_reg ,
  \nz.mem_1113_sv2v_reg ,\nz.mem_1112_sv2v_reg ,\nz.mem_1111_sv2v_reg ,
  \nz.mem_1110_sv2v_reg ,\nz.mem_1109_sv2v_reg ,\nz.mem_1108_sv2v_reg ,\nz.mem_1107_sv2v_reg ,
  \nz.mem_1106_sv2v_reg ,\nz.mem_1105_sv2v_reg ,\nz.mem_1104_sv2v_reg ,
  \nz.mem_1103_sv2v_reg ,\nz.mem_1102_sv2v_reg ,\nz.mem_1101_sv2v_reg ,\nz.mem_1100_sv2v_reg ,
  \nz.mem_1099_sv2v_reg ,\nz.mem_1098_sv2v_reg ,\nz.mem_1097_sv2v_reg ,
  \nz.mem_1096_sv2v_reg ,\nz.mem_1095_sv2v_reg ,\nz.mem_1094_sv2v_reg ,\nz.mem_1093_sv2v_reg ,
  \nz.mem_1092_sv2v_reg ,\nz.mem_1091_sv2v_reg ,\nz.mem_1090_sv2v_reg ,
  \nz.mem_1089_sv2v_reg ,\nz.mem_1088_sv2v_reg ,\nz.mem_1087_sv2v_reg ,\nz.mem_1086_sv2v_reg ,
  \nz.mem_1085_sv2v_reg ,\nz.mem_1084_sv2v_reg ,\nz.mem_1083_sv2v_reg ,
  \nz.mem_1082_sv2v_reg ,\nz.mem_1081_sv2v_reg ,\nz.mem_1080_sv2v_reg ,\nz.mem_1079_sv2v_reg ,
  \nz.mem_1078_sv2v_reg ,\nz.mem_1077_sv2v_reg ,\nz.mem_1076_sv2v_reg ,
  \nz.mem_1075_sv2v_reg ,\nz.mem_1074_sv2v_reg ,\nz.mem_1073_sv2v_reg ,\nz.mem_1072_sv2v_reg ,
  \nz.mem_1071_sv2v_reg ,\nz.mem_1070_sv2v_reg ,\nz.mem_1069_sv2v_reg ,
  \nz.mem_1068_sv2v_reg ,\nz.mem_1067_sv2v_reg ,\nz.mem_1066_sv2v_reg ,
  \nz.mem_1065_sv2v_reg ,\nz.mem_1064_sv2v_reg ,\nz.mem_1063_sv2v_reg ,\nz.mem_1062_sv2v_reg ,
  \nz.mem_1061_sv2v_reg ,\nz.mem_1060_sv2v_reg ,\nz.mem_1059_sv2v_reg ,
  \nz.mem_1058_sv2v_reg ,\nz.mem_1057_sv2v_reg ,\nz.mem_1056_sv2v_reg ,\nz.mem_1055_sv2v_reg ,
  \nz.mem_1054_sv2v_reg ,\nz.mem_1053_sv2v_reg ,\nz.mem_1052_sv2v_reg ,
  \nz.mem_1051_sv2v_reg ,\nz.mem_1050_sv2v_reg ,\nz.mem_1049_sv2v_reg ,\nz.mem_1048_sv2v_reg ,
  \nz.mem_1047_sv2v_reg ,\nz.mem_1046_sv2v_reg ,\nz.mem_1045_sv2v_reg ,
  \nz.mem_1044_sv2v_reg ,\nz.mem_1043_sv2v_reg ,\nz.mem_1042_sv2v_reg ,\nz.mem_1041_sv2v_reg ,
  \nz.mem_1040_sv2v_reg ,\nz.mem_1039_sv2v_reg ,\nz.mem_1038_sv2v_reg ,
  \nz.mem_1037_sv2v_reg ,\nz.mem_1036_sv2v_reg ,\nz.mem_1035_sv2v_reg ,\nz.mem_1034_sv2v_reg ,
  \nz.mem_1033_sv2v_reg ,\nz.mem_1032_sv2v_reg ,\nz.mem_1031_sv2v_reg ,
  \nz.mem_1030_sv2v_reg ,\nz.mem_1029_sv2v_reg ,\nz.mem_1028_sv2v_reg ,\nz.mem_1027_sv2v_reg ,
  \nz.mem_1026_sv2v_reg ,\nz.mem_1025_sv2v_reg ,\nz.mem_1024_sv2v_reg ,
  \nz.mem_1023_sv2v_reg ,\nz.mem_1022_sv2v_reg ,\nz.mem_1021_sv2v_reg ,\nz.mem_1020_sv2v_reg ,
  \nz.mem_1019_sv2v_reg ,\nz.mem_1018_sv2v_reg ,\nz.mem_1017_sv2v_reg ,
  \nz.mem_1016_sv2v_reg ,\nz.mem_1015_sv2v_reg ,\nz.mem_1014_sv2v_reg ,\nz.mem_1013_sv2v_reg ,
  \nz.mem_1012_sv2v_reg ,\nz.mem_1011_sv2v_reg ,\nz.mem_1010_sv2v_reg ,
  \nz.mem_1009_sv2v_reg ,\nz.mem_1008_sv2v_reg ,\nz.mem_1007_sv2v_reg ,\nz.mem_1006_sv2v_reg ,
  \nz.mem_1005_sv2v_reg ,\nz.mem_1004_sv2v_reg ,\nz.mem_1003_sv2v_reg ,
  \nz.mem_1002_sv2v_reg ,\nz.mem_1001_sv2v_reg ,\nz.mem_1000_sv2v_reg ,\nz.mem_999_sv2v_reg ,
  \nz.mem_998_sv2v_reg ,\nz.mem_997_sv2v_reg ,\nz.mem_996_sv2v_reg ,
  \nz.mem_995_sv2v_reg ,\nz.mem_994_sv2v_reg ,\nz.mem_993_sv2v_reg ,\nz.mem_992_sv2v_reg ,
  \nz.mem_991_sv2v_reg ,\nz.mem_990_sv2v_reg ,\nz.mem_989_sv2v_reg ,\nz.mem_988_sv2v_reg ,
  \nz.mem_987_sv2v_reg ,\nz.mem_986_sv2v_reg ,\nz.mem_985_sv2v_reg ,
  \nz.mem_984_sv2v_reg ,\nz.mem_983_sv2v_reg ,\nz.mem_982_sv2v_reg ,\nz.mem_981_sv2v_reg ,
  \nz.mem_980_sv2v_reg ,\nz.mem_979_sv2v_reg ,\nz.mem_978_sv2v_reg ,
  \nz.mem_977_sv2v_reg ,\nz.mem_976_sv2v_reg ,\nz.mem_975_sv2v_reg ,\nz.mem_974_sv2v_reg ,
  \nz.mem_973_sv2v_reg ,\nz.mem_972_sv2v_reg ,\nz.mem_971_sv2v_reg ,\nz.mem_970_sv2v_reg ,
  \nz.mem_969_sv2v_reg ,\nz.mem_968_sv2v_reg ,\nz.mem_967_sv2v_reg ,
  \nz.mem_966_sv2v_reg ,\nz.mem_965_sv2v_reg ,\nz.mem_964_sv2v_reg ,\nz.mem_963_sv2v_reg ,
  \nz.mem_962_sv2v_reg ,\nz.mem_961_sv2v_reg ,\nz.mem_960_sv2v_reg ,\nz.mem_959_sv2v_reg ,
  \nz.mem_958_sv2v_reg ,\nz.mem_957_sv2v_reg ,\nz.mem_956_sv2v_reg ,
  \nz.mem_955_sv2v_reg ,\nz.mem_954_sv2v_reg ,\nz.mem_953_sv2v_reg ,\nz.mem_952_sv2v_reg ,
  \nz.mem_951_sv2v_reg ,\nz.mem_950_sv2v_reg ,\nz.mem_949_sv2v_reg ,\nz.mem_948_sv2v_reg ,
  \nz.mem_947_sv2v_reg ,\nz.mem_946_sv2v_reg ,\nz.mem_945_sv2v_reg ,
  \nz.mem_944_sv2v_reg ,\nz.mem_943_sv2v_reg ,\nz.mem_942_sv2v_reg ,\nz.mem_941_sv2v_reg ,
  \nz.mem_940_sv2v_reg ,\nz.mem_939_sv2v_reg ,\nz.mem_938_sv2v_reg ,
  \nz.mem_937_sv2v_reg ,\nz.mem_936_sv2v_reg ,\nz.mem_935_sv2v_reg ,\nz.mem_934_sv2v_reg ,
  \nz.mem_933_sv2v_reg ,\nz.mem_932_sv2v_reg ,\nz.mem_931_sv2v_reg ,\nz.mem_930_sv2v_reg ,
  \nz.mem_929_sv2v_reg ,\nz.mem_928_sv2v_reg ,\nz.mem_927_sv2v_reg ,
  \nz.mem_926_sv2v_reg ,\nz.mem_925_sv2v_reg ,\nz.mem_924_sv2v_reg ,\nz.mem_923_sv2v_reg ,
  \nz.mem_922_sv2v_reg ,\nz.mem_921_sv2v_reg ,\nz.mem_920_sv2v_reg ,\nz.mem_919_sv2v_reg ,
  \nz.mem_918_sv2v_reg ,\nz.mem_917_sv2v_reg ,\nz.mem_916_sv2v_reg ,
  \nz.mem_915_sv2v_reg ,\nz.mem_914_sv2v_reg ,\nz.mem_913_sv2v_reg ,\nz.mem_912_sv2v_reg ,
  \nz.mem_911_sv2v_reg ,\nz.mem_910_sv2v_reg ,\nz.mem_909_sv2v_reg ,\nz.mem_908_sv2v_reg ,
  \nz.mem_907_sv2v_reg ,\nz.mem_906_sv2v_reg ,\nz.mem_905_sv2v_reg ,
  \nz.mem_904_sv2v_reg ,\nz.mem_903_sv2v_reg ,\nz.mem_902_sv2v_reg ,\nz.mem_901_sv2v_reg ,
  \nz.mem_900_sv2v_reg ,\nz.mem_899_sv2v_reg ,\nz.mem_898_sv2v_reg ,
  \nz.mem_897_sv2v_reg ,\nz.mem_896_sv2v_reg ,\nz.mem_895_sv2v_reg ,\nz.mem_894_sv2v_reg ,
  \nz.mem_893_sv2v_reg ,\nz.mem_892_sv2v_reg ,\nz.mem_891_sv2v_reg ,\nz.mem_890_sv2v_reg ,
  \nz.mem_889_sv2v_reg ,\nz.mem_888_sv2v_reg ,\nz.mem_887_sv2v_reg ,
  \nz.mem_886_sv2v_reg ,\nz.mem_885_sv2v_reg ,\nz.mem_884_sv2v_reg ,\nz.mem_883_sv2v_reg ,
  \nz.mem_882_sv2v_reg ,\nz.mem_881_sv2v_reg ,\nz.mem_880_sv2v_reg ,\nz.mem_879_sv2v_reg ,
  \nz.mem_878_sv2v_reg ,\nz.mem_877_sv2v_reg ,\nz.mem_876_sv2v_reg ,
  \nz.mem_875_sv2v_reg ,\nz.mem_874_sv2v_reg ,\nz.mem_873_sv2v_reg ,\nz.mem_872_sv2v_reg ,
  \nz.mem_871_sv2v_reg ,\nz.mem_870_sv2v_reg ,\nz.mem_869_sv2v_reg ,\nz.mem_868_sv2v_reg ,
  \nz.mem_867_sv2v_reg ,\nz.mem_866_sv2v_reg ,\nz.mem_865_sv2v_reg ,
  \nz.mem_864_sv2v_reg ,\nz.mem_863_sv2v_reg ,\nz.mem_862_sv2v_reg ,\nz.mem_861_sv2v_reg ,
  \nz.mem_860_sv2v_reg ,\nz.mem_859_sv2v_reg ,\nz.mem_858_sv2v_reg ,
  \nz.mem_857_sv2v_reg ,\nz.mem_856_sv2v_reg ,\nz.mem_855_sv2v_reg ,\nz.mem_854_sv2v_reg ,
  \nz.mem_853_sv2v_reg ,\nz.mem_852_sv2v_reg ,\nz.mem_851_sv2v_reg ,\nz.mem_850_sv2v_reg ,
  \nz.mem_849_sv2v_reg ,\nz.mem_848_sv2v_reg ,\nz.mem_847_sv2v_reg ,
  \nz.mem_846_sv2v_reg ,\nz.mem_845_sv2v_reg ,\nz.mem_844_sv2v_reg ,\nz.mem_843_sv2v_reg ,
  \nz.mem_842_sv2v_reg ,\nz.mem_841_sv2v_reg ,\nz.mem_840_sv2v_reg ,\nz.mem_839_sv2v_reg ,
  \nz.mem_838_sv2v_reg ,\nz.mem_837_sv2v_reg ,\nz.mem_836_sv2v_reg ,
  \nz.mem_835_sv2v_reg ,\nz.mem_834_sv2v_reg ,\nz.mem_833_sv2v_reg ,\nz.mem_832_sv2v_reg ,
  \nz.mem_831_sv2v_reg ,\nz.mem_830_sv2v_reg ,\nz.mem_829_sv2v_reg ,\nz.mem_828_sv2v_reg ,
  \nz.mem_827_sv2v_reg ,\nz.mem_826_sv2v_reg ,\nz.mem_825_sv2v_reg ,
  \nz.mem_824_sv2v_reg ,\nz.mem_823_sv2v_reg ,\nz.mem_822_sv2v_reg ,\nz.mem_821_sv2v_reg ,
  \nz.mem_820_sv2v_reg ,\nz.mem_819_sv2v_reg ,\nz.mem_818_sv2v_reg ,
  \nz.mem_817_sv2v_reg ,\nz.mem_816_sv2v_reg ,\nz.mem_815_sv2v_reg ,\nz.mem_814_sv2v_reg ,
  \nz.mem_813_sv2v_reg ,\nz.mem_812_sv2v_reg ,\nz.mem_811_sv2v_reg ,\nz.mem_810_sv2v_reg ,
  \nz.mem_809_sv2v_reg ,\nz.mem_808_sv2v_reg ,\nz.mem_807_sv2v_reg ,
  \nz.mem_806_sv2v_reg ,\nz.mem_805_sv2v_reg ,\nz.mem_804_sv2v_reg ,\nz.mem_803_sv2v_reg ,
  \nz.mem_802_sv2v_reg ,\nz.mem_801_sv2v_reg ,\nz.mem_800_sv2v_reg ,\nz.mem_799_sv2v_reg ,
  \nz.mem_798_sv2v_reg ,\nz.mem_797_sv2v_reg ,\nz.mem_796_sv2v_reg ,
  \nz.mem_795_sv2v_reg ,\nz.mem_794_sv2v_reg ,\nz.mem_793_sv2v_reg ,\nz.mem_792_sv2v_reg ,
  \nz.mem_791_sv2v_reg ,\nz.mem_790_sv2v_reg ,\nz.mem_789_sv2v_reg ,\nz.mem_788_sv2v_reg ,
  \nz.mem_787_sv2v_reg ,\nz.mem_786_sv2v_reg ,\nz.mem_785_sv2v_reg ,
  \nz.mem_784_sv2v_reg ,\nz.mem_783_sv2v_reg ,\nz.mem_782_sv2v_reg ,\nz.mem_781_sv2v_reg ,
  \nz.mem_780_sv2v_reg ,\nz.mem_779_sv2v_reg ,\nz.mem_778_sv2v_reg ,
  \nz.mem_777_sv2v_reg ,\nz.mem_776_sv2v_reg ,\nz.mem_775_sv2v_reg ,\nz.mem_774_sv2v_reg ,
  \nz.mem_773_sv2v_reg ,\nz.mem_772_sv2v_reg ,\nz.mem_771_sv2v_reg ,\nz.mem_770_sv2v_reg ,
  \nz.mem_769_sv2v_reg ,\nz.mem_768_sv2v_reg ,\nz.mem_767_sv2v_reg ,
  \nz.mem_766_sv2v_reg ,\nz.mem_765_sv2v_reg ,\nz.mem_764_sv2v_reg ,\nz.mem_763_sv2v_reg ,
  \nz.mem_762_sv2v_reg ,\nz.mem_761_sv2v_reg ,\nz.mem_760_sv2v_reg ,\nz.mem_759_sv2v_reg ,
  \nz.mem_758_sv2v_reg ,\nz.mem_757_sv2v_reg ,\nz.mem_756_sv2v_reg ,
  \nz.mem_755_sv2v_reg ,\nz.mem_754_sv2v_reg ,\nz.mem_753_sv2v_reg ,\nz.mem_752_sv2v_reg ,
  \nz.mem_751_sv2v_reg ,\nz.mem_750_sv2v_reg ,\nz.mem_749_sv2v_reg ,\nz.mem_748_sv2v_reg ,
  \nz.mem_747_sv2v_reg ,\nz.mem_746_sv2v_reg ,\nz.mem_745_sv2v_reg ,
  \nz.mem_744_sv2v_reg ,\nz.mem_743_sv2v_reg ,\nz.mem_742_sv2v_reg ,\nz.mem_741_sv2v_reg ,
  \nz.mem_740_sv2v_reg ,\nz.mem_739_sv2v_reg ,\nz.mem_738_sv2v_reg ,
  \nz.mem_737_sv2v_reg ,\nz.mem_736_sv2v_reg ,\nz.mem_735_sv2v_reg ,\nz.mem_734_sv2v_reg ,
  \nz.mem_733_sv2v_reg ,\nz.mem_732_sv2v_reg ,\nz.mem_731_sv2v_reg ,\nz.mem_730_sv2v_reg ,
  \nz.mem_729_sv2v_reg ,\nz.mem_728_sv2v_reg ,\nz.mem_727_sv2v_reg ,
  \nz.mem_726_sv2v_reg ,\nz.mem_725_sv2v_reg ,\nz.mem_724_sv2v_reg ,\nz.mem_723_sv2v_reg ,
  \nz.mem_722_sv2v_reg ,\nz.mem_721_sv2v_reg ,\nz.mem_720_sv2v_reg ,\nz.mem_719_sv2v_reg ,
  \nz.mem_718_sv2v_reg ,\nz.mem_717_sv2v_reg ,\nz.mem_716_sv2v_reg ,
  \nz.mem_715_sv2v_reg ,\nz.mem_714_sv2v_reg ,\nz.mem_713_sv2v_reg ,\nz.mem_712_sv2v_reg ,
  \nz.mem_711_sv2v_reg ,\nz.mem_710_sv2v_reg ,\nz.mem_709_sv2v_reg ,\nz.mem_708_sv2v_reg ,
  \nz.mem_707_sv2v_reg ,\nz.mem_706_sv2v_reg ,\nz.mem_705_sv2v_reg ,
  \nz.mem_704_sv2v_reg ,\nz.mem_703_sv2v_reg ,\nz.mem_702_sv2v_reg ,\nz.mem_701_sv2v_reg ,
  \nz.mem_700_sv2v_reg ,\nz.mem_699_sv2v_reg ,\nz.mem_698_sv2v_reg ,
  \nz.mem_697_sv2v_reg ,\nz.mem_696_sv2v_reg ,\nz.mem_695_sv2v_reg ,\nz.mem_694_sv2v_reg ,
  \nz.mem_693_sv2v_reg ,\nz.mem_692_sv2v_reg ,\nz.mem_691_sv2v_reg ,\nz.mem_690_sv2v_reg ,
  \nz.mem_689_sv2v_reg ,\nz.mem_688_sv2v_reg ,\nz.mem_687_sv2v_reg ,
  \nz.mem_686_sv2v_reg ,\nz.mem_685_sv2v_reg ,\nz.mem_684_sv2v_reg ,\nz.mem_683_sv2v_reg ,
  \nz.mem_682_sv2v_reg ,\nz.mem_681_sv2v_reg ,\nz.mem_680_sv2v_reg ,\nz.mem_679_sv2v_reg ,
  \nz.mem_678_sv2v_reg ,\nz.mem_677_sv2v_reg ,\nz.mem_676_sv2v_reg ,
  \nz.mem_675_sv2v_reg ,\nz.mem_674_sv2v_reg ,\nz.mem_673_sv2v_reg ,\nz.mem_672_sv2v_reg ,
  \nz.mem_671_sv2v_reg ,\nz.mem_670_sv2v_reg ,\nz.mem_669_sv2v_reg ,\nz.mem_668_sv2v_reg ,
  \nz.mem_667_sv2v_reg ,\nz.mem_666_sv2v_reg ,\nz.mem_665_sv2v_reg ,
  \nz.mem_664_sv2v_reg ,\nz.mem_663_sv2v_reg ,\nz.mem_662_sv2v_reg ,\nz.mem_661_sv2v_reg ,
  \nz.mem_660_sv2v_reg ,\nz.mem_659_sv2v_reg ,\nz.mem_658_sv2v_reg ,
  \nz.mem_657_sv2v_reg ,\nz.mem_656_sv2v_reg ,\nz.mem_655_sv2v_reg ,\nz.mem_654_sv2v_reg ,
  \nz.mem_653_sv2v_reg ,\nz.mem_652_sv2v_reg ,\nz.mem_651_sv2v_reg ,\nz.mem_650_sv2v_reg ,
  \nz.mem_649_sv2v_reg ,\nz.mem_648_sv2v_reg ,\nz.mem_647_sv2v_reg ,
  \nz.mem_646_sv2v_reg ,\nz.mem_645_sv2v_reg ,\nz.mem_644_sv2v_reg ,\nz.mem_643_sv2v_reg ,
  \nz.mem_642_sv2v_reg ,\nz.mem_641_sv2v_reg ,\nz.mem_640_sv2v_reg ,\nz.mem_639_sv2v_reg ,
  \nz.mem_638_sv2v_reg ,\nz.mem_637_sv2v_reg ,\nz.mem_636_sv2v_reg ,
  \nz.mem_635_sv2v_reg ,\nz.mem_634_sv2v_reg ,\nz.mem_633_sv2v_reg ,\nz.mem_632_sv2v_reg ,
  \nz.mem_631_sv2v_reg ,\nz.mem_630_sv2v_reg ,\nz.mem_629_sv2v_reg ,\nz.mem_628_sv2v_reg ,
  \nz.mem_627_sv2v_reg ,\nz.mem_626_sv2v_reg ,\nz.mem_625_sv2v_reg ,
  \nz.mem_624_sv2v_reg ,\nz.mem_623_sv2v_reg ,\nz.mem_622_sv2v_reg ,\nz.mem_621_sv2v_reg ,
  \nz.mem_620_sv2v_reg ,\nz.mem_619_sv2v_reg ,\nz.mem_618_sv2v_reg ,
  \nz.mem_617_sv2v_reg ,\nz.mem_616_sv2v_reg ,\nz.mem_615_sv2v_reg ,\nz.mem_614_sv2v_reg ,
  \nz.mem_613_sv2v_reg ,\nz.mem_612_sv2v_reg ,\nz.mem_611_sv2v_reg ,\nz.mem_610_sv2v_reg ,
  \nz.mem_609_sv2v_reg ,\nz.mem_608_sv2v_reg ,\nz.mem_607_sv2v_reg ,
  \nz.mem_606_sv2v_reg ,\nz.mem_605_sv2v_reg ,\nz.mem_604_sv2v_reg ,\nz.mem_603_sv2v_reg ,
  \nz.mem_602_sv2v_reg ,\nz.mem_601_sv2v_reg ,\nz.mem_600_sv2v_reg ,\nz.mem_599_sv2v_reg ,
  \nz.mem_598_sv2v_reg ,\nz.mem_597_sv2v_reg ,\nz.mem_596_sv2v_reg ,
  \nz.mem_595_sv2v_reg ,\nz.mem_594_sv2v_reg ,\nz.mem_593_sv2v_reg ,\nz.mem_592_sv2v_reg ,
  \nz.mem_591_sv2v_reg ,\nz.mem_590_sv2v_reg ,\nz.mem_589_sv2v_reg ,\nz.mem_588_sv2v_reg ,
  \nz.mem_587_sv2v_reg ,\nz.mem_586_sv2v_reg ,\nz.mem_585_sv2v_reg ,
  \nz.mem_584_sv2v_reg ,\nz.mem_583_sv2v_reg ,\nz.mem_582_sv2v_reg ,\nz.mem_581_sv2v_reg ,
  \nz.mem_580_sv2v_reg ,\nz.mem_579_sv2v_reg ,\nz.mem_578_sv2v_reg ,
  \nz.mem_577_sv2v_reg ,\nz.mem_576_sv2v_reg ,\nz.mem_575_sv2v_reg ,\nz.mem_574_sv2v_reg ,
  \nz.mem_573_sv2v_reg ,\nz.mem_572_sv2v_reg ,\nz.mem_571_sv2v_reg ,\nz.mem_570_sv2v_reg ,
  \nz.mem_569_sv2v_reg ,\nz.mem_568_sv2v_reg ,\nz.mem_567_sv2v_reg ,
  \nz.mem_566_sv2v_reg ,\nz.mem_565_sv2v_reg ,\nz.mem_564_sv2v_reg ,\nz.mem_563_sv2v_reg ,
  \nz.mem_562_sv2v_reg ,\nz.mem_561_sv2v_reg ,\nz.mem_560_sv2v_reg ,\nz.mem_559_sv2v_reg ,
  \nz.mem_558_sv2v_reg ,\nz.mem_557_sv2v_reg ,\nz.mem_556_sv2v_reg ,
  \nz.mem_555_sv2v_reg ,\nz.mem_554_sv2v_reg ,\nz.mem_553_sv2v_reg ,\nz.mem_552_sv2v_reg ,
  \nz.mem_551_sv2v_reg ,\nz.mem_550_sv2v_reg ,\nz.mem_549_sv2v_reg ,\nz.mem_548_sv2v_reg ,
  \nz.mem_547_sv2v_reg ,\nz.mem_546_sv2v_reg ,\nz.mem_545_sv2v_reg ,
  \nz.mem_544_sv2v_reg ,\nz.mem_543_sv2v_reg ,\nz.mem_542_sv2v_reg ,\nz.mem_541_sv2v_reg ,
  \nz.mem_540_sv2v_reg ,\nz.mem_539_sv2v_reg ,\nz.mem_538_sv2v_reg ,
  \nz.mem_537_sv2v_reg ,\nz.mem_536_sv2v_reg ,\nz.mem_535_sv2v_reg ,\nz.mem_534_sv2v_reg ,
  \nz.mem_533_sv2v_reg ,\nz.mem_532_sv2v_reg ,\nz.mem_531_sv2v_reg ,\nz.mem_530_sv2v_reg ,
  \nz.mem_529_sv2v_reg ,\nz.mem_528_sv2v_reg ,\nz.mem_527_sv2v_reg ,
  \nz.mem_526_sv2v_reg ,\nz.mem_525_sv2v_reg ,\nz.mem_524_sv2v_reg ,\nz.mem_523_sv2v_reg ,
  \nz.mem_522_sv2v_reg ,\nz.mem_521_sv2v_reg ,\nz.mem_520_sv2v_reg ,\nz.mem_519_sv2v_reg ,
  \nz.mem_518_sv2v_reg ,\nz.mem_517_sv2v_reg ,\nz.mem_516_sv2v_reg ,
  \nz.mem_515_sv2v_reg ,\nz.mem_514_sv2v_reg ,\nz.mem_513_sv2v_reg ,\nz.mem_512_sv2v_reg ,
  \nz.mem_511_sv2v_reg ,\nz.mem_510_sv2v_reg ,\nz.mem_509_sv2v_reg ,\nz.mem_508_sv2v_reg ,
  \nz.mem_507_sv2v_reg ,\nz.mem_506_sv2v_reg ,\nz.mem_505_sv2v_reg ,
  \nz.mem_504_sv2v_reg ,\nz.mem_503_sv2v_reg ,\nz.mem_502_sv2v_reg ,\nz.mem_501_sv2v_reg ,
  \nz.mem_500_sv2v_reg ,\nz.mem_499_sv2v_reg ,\nz.mem_498_sv2v_reg ,
  \nz.mem_497_sv2v_reg ,\nz.mem_496_sv2v_reg ,\nz.mem_495_sv2v_reg ,\nz.mem_494_sv2v_reg ,
  \nz.mem_493_sv2v_reg ,\nz.mem_492_sv2v_reg ,\nz.mem_491_sv2v_reg ,\nz.mem_490_sv2v_reg ,
  \nz.mem_489_sv2v_reg ,\nz.mem_488_sv2v_reg ,\nz.mem_487_sv2v_reg ,
  \nz.mem_486_sv2v_reg ,\nz.mem_485_sv2v_reg ,\nz.mem_484_sv2v_reg ,\nz.mem_483_sv2v_reg ,
  \nz.mem_482_sv2v_reg ,\nz.mem_481_sv2v_reg ,\nz.mem_480_sv2v_reg ,\nz.mem_479_sv2v_reg ,
  \nz.mem_478_sv2v_reg ,\nz.mem_477_sv2v_reg ,\nz.mem_476_sv2v_reg ,
  \nz.mem_475_sv2v_reg ,\nz.mem_474_sv2v_reg ,\nz.mem_473_sv2v_reg ,\nz.mem_472_sv2v_reg ,
  \nz.mem_471_sv2v_reg ,\nz.mem_470_sv2v_reg ,\nz.mem_469_sv2v_reg ,\nz.mem_468_sv2v_reg ,
  \nz.mem_467_sv2v_reg ,\nz.mem_466_sv2v_reg ,\nz.mem_465_sv2v_reg ,
  \nz.mem_464_sv2v_reg ,\nz.mem_463_sv2v_reg ,\nz.mem_462_sv2v_reg ,\nz.mem_461_sv2v_reg ,
  \nz.mem_460_sv2v_reg ,\nz.mem_459_sv2v_reg ,\nz.mem_458_sv2v_reg ,
  \nz.mem_457_sv2v_reg ,\nz.mem_456_sv2v_reg ,\nz.mem_455_sv2v_reg ,\nz.mem_454_sv2v_reg ,
  \nz.mem_453_sv2v_reg ,\nz.mem_452_sv2v_reg ,\nz.mem_451_sv2v_reg ,\nz.mem_450_sv2v_reg ,
  \nz.mem_449_sv2v_reg ,\nz.mem_448_sv2v_reg ,\nz.mem_447_sv2v_reg ,
  \nz.mem_446_sv2v_reg ,\nz.mem_445_sv2v_reg ,\nz.mem_444_sv2v_reg ,\nz.mem_443_sv2v_reg ,
  \nz.mem_442_sv2v_reg ,\nz.mem_441_sv2v_reg ,\nz.mem_440_sv2v_reg ,\nz.mem_439_sv2v_reg ,
  \nz.mem_438_sv2v_reg ,\nz.mem_437_sv2v_reg ,\nz.mem_436_sv2v_reg ,
  \nz.mem_435_sv2v_reg ,\nz.mem_434_sv2v_reg ,\nz.mem_433_sv2v_reg ,\nz.mem_432_sv2v_reg ,
  \nz.mem_431_sv2v_reg ,\nz.mem_430_sv2v_reg ,\nz.mem_429_sv2v_reg ,\nz.mem_428_sv2v_reg ,
  \nz.mem_427_sv2v_reg ,\nz.mem_426_sv2v_reg ,\nz.mem_425_sv2v_reg ,
  \nz.mem_424_sv2v_reg ,\nz.mem_423_sv2v_reg ,\nz.mem_422_sv2v_reg ,\nz.mem_421_sv2v_reg ,
  \nz.mem_420_sv2v_reg ,\nz.mem_419_sv2v_reg ,\nz.mem_418_sv2v_reg ,
  \nz.mem_417_sv2v_reg ,\nz.mem_416_sv2v_reg ,\nz.mem_415_sv2v_reg ,\nz.mem_414_sv2v_reg ,
  \nz.mem_413_sv2v_reg ,\nz.mem_412_sv2v_reg ,\nz.mem_411_sv2v_reg ,\nz.mem_410_sv2v_reg ,
  \nz.mem_409_sv2v_reg ,\nz.mem_408_sv2v_reg ,\nz.mem_407_sv2v_reg ,
  \nz.mem_406_sv2v_reg ,\nz.mem_405_sv2v_reg ,\nz.mem_404_sv2v_reg ,\nz.mem_403_sv2v_reg ,
  \nz.mem_402_sv2v_reg ,\nz.mem_401_sv2v_reg ,\nz.mem_400_sv2v_reg ,\nz.mem_399_sv2v_reg ,
  \nz.mem_398_sv2v_reg ,\nz.mem_397_sv2v_reg ,\nz.mem_396_sv2v_reg ,
  \nz.mem_395_sv2v_reg ,\nz.mem_394_sv2v_reg ,\nz.mem_393_sv2v_reg ,\nz.mem_392_sv2v_reg ,
  \nz.mem_391_sv2v_reg ,\nz.mem_390_sv2v_reg ,\nz.mem_389_sv2v_reg ,\nz.mem_388_sv2v_reg ,
  \nz.mem_387_sv2v_reg ,\nz.mem_386_sv2v_reg ,\nz.mem_385_sv2v_reg ,
  \nz.mem_384_sv2v_reg ,\nz.mem_383_sv2v_reg ,\nz.mem_382_sv2v_reg ,\nz.mem_381_sv2v_reg ,
  \nz.mem_380_sv2v_reg ,\nz.mem_379_sv2v_reg ,\nz.mem_378_sv2v_reg ,
  \nz.mem_377_sv2v_reg ,\nz.mem_376_sv2v_reg ,\nz.mem_375_sv2v_reg ,\nz.mem_374_sv2v_reg ,
  \nz.mem_373_sv2v_reg ,\nz.mem_372_sv2v_reg ,\nz.mem_371_sv2v_reg ,\nz.mem_370_sv2v_reg ,
  \nz.mem_369_sv2v_reg ,\nz.mem_368_sv2v_reg ,\nz.mem_367_sv2v_reg ,
  \nz.mem_366_sv2v_reg ,\nz.mem_365_sv2v_reg ,\nz.mem_364_sv2v_reg ,\nz.mem_363_sv2v_reg ,
  \nz.mem_362_sv2v_reg ,\nz.mem_361_sv2v_reg ,\nz.mem_360_sv2v_reg ,\nz.mem_359_sv2v_reg ,
  \nz.mem_358_sv2v_reg ,\nz.mem_357_sv2v_reg ,\nz.mem_356_sv2v_reg ,
  \nz.mem_355_sv2v_reg ,\nz.mem_354_sv2v_reg ,\nz.mem_353_sv2v_reg ,\nz.mem_352_sv2v_reg ,
  \nz.mem_351_sv2v_reg ,\nz.mem_350_sv2v_reg ,\nz.mem_349_sv2v_reg ,\nz.mem_348_sv2v_reg ,
  \nz.mem_347_sv2v_reg ,\nz.mem_346_sv2v_reg ,\nz.mem_345_sv2v_reg ,
  \nz.mem_344_sv2v_reg ,\nz.mem_343_sv2v_reg ,\nz.mem_342_sv2v_reg ,\nz.mem_341_sv2v_reg ,
  \nz.mem_340_sv2v_reg ,\nz.mem_339_sv2v_reg ,\nz.mem_338_sv2v_reg ,
  \nz.mem_337_sv2v_reg ,\nz.mem_336_sv2v_reg ,\nz.mem_335_sv2v_reg ,\nz.mem_334_sv2v_reg ,
  \nz.mem_333_sv2v_reg ,\nz.mem_332_sv2v_reg ,\nz.mem_331_sv2v_reg ,\nz.mem_330_sv2v_reg ,
  \nz.mem_329_sv2v_reg ,\nz.mem_328_sv2v_reg ,\nz.mem_327_sv2v_reg ,
  \nz.mem_326_sv2v_reg ,\nz.mem_325_sv2v_reg ,\nz.mem_324_sv2v_reg ,\nz.mem_323_sv2v_reg ,
  \nz.mem_322_sv2v_reg ,\nz.mem_321_sv2v_reg ,\nz.mem_320_sv2v_reg ,\nz.mem_319_sv2v_reg ,
  \nz.mem_318_sv2v_reg ,\nz.mem_317_sv2v_reg ,\nz.mem_316_sv2v_reg ,
  \nz.mem_315_sv2v_reg ,\nz.mem_314_sv2v_reg ,\nz.mem_313_sv2v_reg ,\nz.mem_312_sv2v_reg ,
  \nz.mem_311_sv2v_reg ,\nz.mem_310_sv2v_reg ,\nz.mem_309_sv2v_reg ,\nz.mem_308_sv2v_reg ,
  \nz.mem_307_sv2v_reg ,\nz.mem_306_sv2v_reg ,\nz.mem_305_sv2v_reg ,
  \nz.mem_304_sv2v_reg ,\nz.mem_303_sv2v_reg ,\nz.mem_302_sv2v_reg ,\nz.mem_301_sv2v_reg ,
  \nz.mem_300_sv2v_reg ,\nz.mem_299_sv2v_reg ,\nz.mem_298_sv2v_reg ,
  \nz.mem_297_sv2v_reg ,\nz.mem_296_sv2v_reg ,\nz.mem_295_sv2v_reg ,\nz.mem_294_sv2v_reg ,
  \nz.mem_293_sv2v_reg ,\nz.mem_292_sv2v_reg ,\nz.mem_291_sv2v_reg ,\nz.mem_290_sv2v_reg ,
  \nz.mem_289_sv2v_reg ,\nz.mem_288_sv2v_reg ,\nz.mem_287_sv2v_reg ,
  \nz.mem_286_sv2v_reg ,\nz.mem_285_sv2v_reg ,\nz.mem_284_sv2v_reg ,\nz.mem_283_sv2v_reg ,
  \nz.mem_282_sv2v_reg ,\nz.mem_281_sv2v_reg ,\nz.mem_280_sv2v_reg ,\nz.mem_279_sv2v_reg ,
  \nz.mem_278_sv2v_reg ,\nz.mem_277_sv2v_reg ,\nz.mem_276_sv2v_reg ,
  \nz.mem_275_sv2v_reg ,\nz.mem_274_sv2v_reg ,\nz.mem_273_sv2v_reg ,\nz.mem_272_sv2v_reg ,
  \nz.mem_271_sv2v_reg ,\nz.mem_270_sv2v_reg ,\nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,
  \nz.mem_267_sv2v_reg ,\nz.mem_266_sv2v_reg ,\nz.mem_265_sv2v_reg ,
  \nz.mem_264_sv2v_reg ,\nz.mem_263_sv2v_reg ,\nz.mem_262_sv2v_reg ,\nz.mem_261_sv2v_reg ,
  \nz.mem_260_sv2v_reg ,\nz.mem_259_sv2v_reg ,\nz.mem_258_sv2v_reg ,
  \nz.mem_257_sv2v_reg ,\nz.mem_256_sv2v_reg ,\nz.mem_255_sv2v_reg ,\nz.mem_254_sv2v_reg ,
  \nz.mem_253_sv2v_reg ,\nz.mem_252_sv2v_reg ,\nz.mem_251_sv2v_reg ,\nz.mem_250_sv2v_reg ,
  \nz.mem_249_sv2v_reg ,\nz.mem_248_sv2v_reg ,\nz.mem_247_sv2v_reg ,
  \nz.mem_246_sv2v_reg ,\nz.mem_245_sv2v_reg ,\nz.mem_244_sv2v_reg ,\nz.mem_243_sv2v_reg ,
  \nz.mem_242_sv2v_reg ,\nz.mem_241_sv2v_reg ,\nz.mem_240_sv2v_reg ,\nz.mem_239_sv2v_reg ,
  \nz.mem_238_sv2v_reg ,\nz.mem_237_sv2v_reg ,\nz.mem_236_sv2v_reg ,
  \nz.mem_235_sv2v_reg ,\nz.mem_234_sv2v_reg ,\nz.mem_233_sv2v_reg ,\nz.mem_232_sv2v_reg ,
  \nz.mem_231_sv2v_reg ,\nz.mem_230_sv2v_reg ,\nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,
  \nz.mem_227_sv2v_reg ,\nz.mem_226_sv2v_reg ,\nz.mem_225_sv2v_reg ,
  \nz.mem_224_sv2v_reg ,\nz.mem_223_sv2v_reg ,\nz.mem_222_sv2v_reg ,\nz.mem_221_sv2v_reg ,
  \nz.mem_220_sv2v_reg ,\nz.mem_219_sv2v_reg ,\nz.mem_218_sv2v_reg ,
  \nz.mem_217_sv2v_reg ,\nz.mem_216_sv2v_reg ,\nz.mem_215_sv2v_reg ,\nz.mem_214_sv2v_reg ,
  \nz.mem_213_sv2v_reg ,\nz.mem_212_sv2v_reg ,\nz.mem_211_sv2v_reg ,\nz.mem_210_sv2v_reg ,
  \nz.mem_209_sv2v_reg ,\nz.mem_208_sv2v_reg ,\nz.mem_207_sv2v_reg ,
  \nz.mem_206_sv2v_reg ,\nz.mem_205_sv2v_reg ,\nz.mem_204_sv2v_reg ,\nz.mem_203_sv2v_reg ,
  \nz.mem_202_sv2v_reg ,\nz.mem_201_sv2v_reg ,\nz.mem_200_sv2v_reg ,\nz.mem_199_sv2v_reg ,
  \nz.mem_198_sv2v_reg ,\nz.mem_197_sv2v_reg ,\nz.mem_196_sv2v_reg ,
  \nz.mem_195_sv2v_reg ,\nz.mem_194_sv2v_reg ,\nz.mem_193_sv2v_reg ,\nz.mem_192_sv2v_reg ,
  \nz.mem_191_sv2v_reg ,\nz.mem_190_sv2v_reg ,\nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,
  \nz.mem_187_sv2v_reg ,\nz.mem_186_sv2v_reg ,\nz.mem_185_sv2v_reg ,
  \nz.mem_184_sv2v_reg ,\nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,\nz.mem_181_sv2v_reg ,
  \nz.mem_180_sv2v_reg ,\nz.mem_179_sv2v_reg ,\nz.mem_178_sv2v_reg ,
  \nz.mem_177_sv2v_reg ,\nz.mem_176_sv2v_reg ,\nz.mem_175_sv2v_reg ,\nz.mem_174_sv2v_reg ,
  \nz.mem_173_sv2v_reg ,\nz.mem_172_sv2v_reg ,\nz.mem_171_sv2v_reg ,\nz.mem_170_sv2v_reg ,
  \nz.mem_169_sv2v_reg ,\nz.mem_168_sv2v_reg ,\nz.mem_167_sv2v_reg ,
  \nz.mem_166_sv2v_reg ,\nz.mem_165_sv2v_reg ,\nz.mem_164_sv2v_reg ,\nz.mem_163_sv2v_reg ,
  \nz.mem_162_sv2v_reg ,\nz.mem_161_sv2v_reg ,\nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,
  \nz.mem_158_sv2v_reg ,\nz.mem_157_sv2v_reg ,\nz.mem_156_sv2v_reg ,
  \nz.mem_155_sv2v_reg ,\nz.mem_154_sv2v_reg ,\nz.mem_153_sv2v_reg ,\nz.mem_152_sv2v_reg ,
  \nz.mem_151_sv2v_reg ,\nz.mem_150_sv2v_reg ,\nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,
  \nz.mem_147_sv2v_reg ,\nz.mem_146_sv2v_reg ,\nz.mem_145_sv2v_reg ,
  \nz.mem_144_sv2v_reg ,\nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,\nz.mem_141_sv2v_reg ,
  \nz.mem_140_sv2v_reg ,\nz.mem_139_sv2v_reg ,\nz.mem_138_sv2v_reg ,
  \nz.mem_137_sv2v_reg ,\nz.mem_136_sv2v_reg ,\nz.mem_135_sv2v_reg ,\nz.mem_134_sv2v_reg ,
  \nz.mem_133_sv2v_reg ,\nz.mem_132_sv2v_reg ,\nz.mem_131_sv2v_reg ,\nz.mem_130_sv2v_reg ,
  \nz.mem_129_sv2v_reg ,\nz.mem_128_sv2v_reg ,\nz.mem_127_sv2v_reg ,
  \nz.mem_126_sv2v_reg ,\nz.mem_125_sv2v_reg ,\nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,
  \nz.mem_122_sv2v_reg ,\nz.mem_121_sv2v_reg ,\nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,
  \nz.mem_118_sv2v_reg ,\nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,
  \nz.mem_115_sv2v_reg ,\nz.mem_114_sv2v_reg ,\nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,
  \nz.mem_111_sv2v_reg ,\nz.mem_110_sv2v_reg ,\nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,
  \nz.mem_107_sv2v_reg ,\nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,
  \nz.mem_104_sv2v_reg ,\nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,
  \nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,\nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,
  \nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,
  \nz.mem_93_sv2v_reg ,\nz.mem_92_sv2v_reg ,\nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,
  \nz.mem_89_sv2v_reg ,\nz.mem_88_sv2v_reg ,\nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,
  \nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,\nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,
  \nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,\nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,
  \nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,\nz.mem_75_sv2v_reg ,
  \nz.mem_74_sv2v_reg ,\nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,
  \nz.mem_70_sv2v_reg ,\nz.mem_69_sv2v_reg ,\nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,
  \nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,
  \nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,\nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,
  \nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,\nz.mem_56_sv2v_reg ,
  \nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,
  \nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,
  \nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,
  \nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,\nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,
  \nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,\nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,
  \nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,
  \nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,
  \nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,
  \nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,\nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,
  \nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,\nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,
  \nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,
  \nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,
  \nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,
  \nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,
  \nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.mem [1391] = \nz.mem_1391_sv2v_reg ;
  assign \nz.mem [1390] = \nz.mem_1390_sv2v_reg ;
  assign \nz.mem [1389] = \nz.mem_1389_sv2v_reg ;
  assign \nz.mem [1388] = \nz.mem_1388_sv2v_reg ;
  assign \nz.mem [1387] = \nz.mem_1387_sv2v_reg ;
  assign \nz.mem [1386] = \nz.mem_1386_sv2v_reg ;
  assign \nz.mem [1385] = \nz.mem_1385_sv2v_reg ;
  assign \nz.mem [1384] = \nz.mem_1384_sv2v_reg ;
  assign \nz.mem [1383] = \nz.mem_1383_sv2v_reg ;
  assign \nz.mem [1382] = \nz.mem_1382_sv2v_reg ;
  assign \nz.mem [1381] = \nz.mem_1381_sv2v_reg ;
  assign \nz.mem [1380] = \nz.mem_1380_sv2v_reg ;
  assign \nz.mem [1379] = \nz.mem_1379_sv2v_reg ;
  assign \nz.mem [1378] = \nz.mem_1378_sv2v_reg ;
  assign \nz.mem [1377] = \nz.mem_1377_sv2v_reg ;
  assign \nz.mem [1376] = \nz.mem_1376_sv2v_reg ;
  assign \nz.mem [1375] = \nz.mem_1375_sv2v_reg ;
  assign \nz.mem [1374] = \nz.mem_1374_sv2v_reg ;
  assign \nz.mem [1373] = \nz.mem_1373_sv2v_reg ;
  assign \nz.mem [1372] = \nz.mem_1372_sv2v_reg ;
  assign \nz.mem [1371] = \nz.mem_1371_sv2v_reg ;
  assign \nz.mem [1370] = \nz.mem_1370_sv2v_reg ;
  assign \nz.mem [1369] = \nz.mem_1369_sv2v_reg ;
  assign \nz.mem [1368] = \nz.mem_1368_sv2v_reg ;
  assign \nz.mem [1367] = \nz.mem_1367_sv2v_reg ;
  assign \nz.mem [1366] = \nz.mem_1366_sv2v_reg ;
  assign \nz.mem [1365] = \nz.mem_1365_sv2v_reg ;
  assign \nz.mem [1364] = \nz.mem_1364_sv2v_reg ;
  assign \nz.mem [1363] = \nz.mem_1363_sv2v_reg ;
  assign \nz.mem [1362] = \nz.mem_1362_sv2v_reg ;
  assign \nz.mem [1361] = \nz.mem_1361_sv2v_reg ;
  assign \nz.mem [1360] = \nz.mem_1360_sv2v_reg ;
  assign \nz.mem [1359] = \nz.mem_1359_sv2v_reg ;
  assign \nz.mem [1358] = \nz.mem_1358_sv2v_reg ;
  assign \nz.mem [1357] = \nz.mem_1357_sv2v_reg ;
  assign \nz.mem [1356] = \nz.mem_1356_sv2v_reg ;
  assign \nz.mem [1355] = \nz.mem_1355_sv2v_reg ;
  assign \nz.mem [1354] = \nz.mem_1354_sv2v_reg ;
  assign \nz.mem [1353] = \nz.mem_1353_sv2v_reg ;
  assign \nz.mem [1352] = \nz.mem_1352_sv2v_reg ;
  assign \nz.mem [1351] = \nz.mem_1351_sv2v_reg ;
  assign \nz.mem [1350] = \nz.mem_1350_sv2v_reg ;
  assign \nz.mem [1349] = \nz.mem_1349_sv2v_reg ;
  assign \nz.mem [1348] = \nz.mem_1348_sv2v_reg ;
  assign \nz.mem [1347] = \nz.mem_1347_sv2v_reg ;
  assign \nz.mem [1346] = \nz.mem_1346_sv2v_reg ;
  assign \nz.mem [1345] = \nz.mem_1345_sv2v_reg ;
  assign \nz.mem [1344] = \nz.mem_1344_sv2v_reg ;
  assign \nz.mem [1343] = \nz.mem_1343_sv2v_reg ;
  assign \nz.mem [1342] = \nz.mem_1342_sv2v_reg ;
  assign \nz.mem [1341] = \nz.mem_1341_sv2v_reg ;
  assign \nz.mem [1340] = \nz.mem_1340_sv2v_reg ;
  assign \nz.mem [1339] = \nz.mem_1339_sv2v_reg ;
  assign \nz.mem [1338] = \nz.mem_1338_sv2v_reg ;
  assign \nz.mem [1337] = \nz.mem_1337_sv2v_reg ;
  assign \nz.mem [1336] = \nz.mem_1336_sv2v_reg ;
  assign \nz.mem [1335] = \nz.mem_1335_sv2v_reg ;
  assign \nz.mem [1334] = \nz.mem_1334_sv2v_reg ;
  assign \nz.mem [1333] = \nz.mem_1333_sv2v_reg ;
  assign \nz.mem [1332] = \nz.mem_1332_sv2v_reg ;
  assign \nz.mem [1331] = \nz.mem_1331_sv2v_reg ;
  assign \nz.mem [1330] = \nz.mem_1330_sv2v_reg ;
  assign \nz.mem [1329] = \nz.mem_1329_sv2v_reg ;
  assign \nz.mem [1328] = \nz.mem_1328_sv2v_reg ;
  assign \nz.mem [1327] = \nz.mem_1327_sv2v_reg ;
  assign \nz.mem [1326] = \nz.mem_1326_sv2v_reg ;
  assign \nz.mem [1325] = \nz.mem_1325_sv2v_reg ;
  assign \nz.mem [1324] = \nz.mem_1324_sv2v_reg ;
  assign \nz.mem [1323] = \nz.mem_1323_sv2v_reg ;
  assign \nz.mem [1322] = \nz.mem_1322_sv2v_reg ;
  assign \nz.mem [1321] = \nz.mem_1321_sv2v_reg ;
  assign \nz.mem [1320] = \nz.mem_1320_sv2v_reg ;
  assign \nz.mem [1319] = \nz.mem_1319_sv2v_reg ;
  assign \nz.mem [1318] = \nz.mem_1318_sv2v_reg ;
  assign \nz.mem [1317] = \nz.mem_1317_sv2v_reg ;
  assign \nz.mem [1316] = \nz.mem_1316_sv2v_reg ;
  assign \nz.mem [1315] = \nz.mem_1315_sv2v_reg ;
  assign \nz.mem [1314] = \nz.mem_1314_sv2v_reg ;
  assign \nz.mem [1313] = \nz.mem_1313_sv2v_reg ;
  assign \nz.mem [1312] = \nz.mem_1312_sv2v_reg ;
  assign \nz.mem [1311] = \nz.mem_1311_sv2v_reg ;
  assign \nz.mem [1310] = \nz.mem_1310_sv2v_reg ;
  assign \nz.mem [1309] = \nz.mem_1309_sv2v_reg ;
  assign \nz.mem [1308] = \nz.mem_1308_sv2v_reg ;
  assign \nz.mem [1307] = \nz.mem_1307_sv2v_reg ;
  assign \nz.mem [1306] = \nz.mem_1306_sv2v_reg ;
  assign \nz.mem [1305] = \nz.mem_1305_sv2v_reg ;
  assign \nz.mem [1304] = \nz.mem_1304_sv2v_reg ;
  assign \nz.mem [1303] = \nz.mem_1303_sv2v_reg ;
  assign \nz.mem [1302] = \nz.mem_1302_sv2v_reg ;
  assign \nz.mem [1301] = \nz.mem_1301_sv2v_reg ;
  assign \nz.mem [1300] = \nz.mem_1300_sv2v_reg ;
  assign \nz.mem [1299] = \nz.mem_1299_sv2v_reg ;
  assign \nz.mem [1298] = \nz.mem_1298_sv2v_reg ;
  assign \nz.mem [1297] = \nz.mem_1297_sv2v_reg ;
  assign \nz.mem [1296] = \nz.mem_1296_sv2v_reg ;
  assign \nz.mem [1295] = \nz.mem_1295_sv2v_reg ;
  assign \nz.mem [1294] = \nz.mem_1294_sv2v_reg ;
  assign \nz.mem [1293] = \nz.mem_1293_sv2v_reg ;
  assign \nz.mem [1292] = \nz.mem_1292_sv2v_reg ;
  assign \nz.mem [1291] = \nz.mem_1291_sv2v_reg ;
  assign \nz.mem [1290] = \nz.mem_1290_sv2v_reg ;
  assign \nz.mem [1289] = \nz.mem_1289_sv2v_reg ;
  assign \nz.mem [1288] = \nz.mem_1288_sv2v_reg ;
  assign \nz.mem [1287] = \nz.mem_1287_sv2v_reg ;
  assign \nz.mem [1286] = \nz.mem_1286_sv2v_reg ;
  assign \nz.mem [1285] = \nz.mem_1285_sv2v_reg ;
  assign \nz.mem [1284] = \nz.mem_1284_sv2v_reg ;
  assign \nz.mem [1283] = \nz.mem_1283_sv2v_reg ;
  assign \nz.mem [1282] = \nz.mem_1282_sv2v_reg ;
  assign \nz.mem [1281] = \nz.mem_1281_sv2v_reg ;
  assign \nz.mem [1280] = \nz.mem_1280_sv2v_reg ;
  assign \nz.mem [1279] = \nz.mem_1279_sv2v_reg ;
  assign \nz.mem [1278] = \nz.mem_1278_sv2v_reg ;
  assign \nz.mem [1277] = \nz.mem_1277_sv2v_reg ;
  assign \nz.mem [1276] = \nz.mem_1276_sv2v_reg ;
  assign \nz.mem [1275] = \nz.mem_1275_sv2v_reg ;
  assign \nz.mem [1274] = \nz.mem_1274_sv2v_reg ;
  assign \nz.mem [1273] = \nz.mem_1273_sv2v_reg ;
  assign \nz.mem [1272] = \nz.mem_1272_sv2v_reg ;
  assign \nz.mem [1271] = \nz.mem_1271_sv2v_reg ;
  assign \nz.mem [1270] = \nz.mem_1270_sv2v_reg ;
  assign \nz.mem [1269] = \nz.mem_1269_sv2v_reg ;
  assign \nz.mem [1268] = \nz.mem_1268_sv2v_reg ;
  assign \nz.mem [1267] = \nz.mem_1267_sv2v_reg ;
  assign \nz.mem [1266] = \nz.mem_1266_sv2v_reg ;
  assign \nz.mem [1265] = \nz.mem_1265_sv2v_reg ;
  assign \nz.mem [1264] = \nz.mem_1264_sv2v_reg ;
  assign \nz.mem [1263] = \nz.mem_1263_sv2v_reg ;
  assign \nz.mem [1262] = \nz.mem_1262_sv2v_reg ;
  assign \nz.mem [1261] = \nz.mem_1261_sv2v_reg ;
  assign \nz.mem [1260] = \nz.mem_1260_sv2v_reg ;
  assign \nz.mem [1259] = \nz.mem_1259_sv2v_reg ;
  assign \nz.mem [1258] = \nz.mem_1258_sv2v_reg ;
  assign \nz.mem [1257] = \nz.mem_1257_sv2v_reg ;
  assign \nz.mem [1256] = \nz.mem_1256_sv2v_reg ;
  assign \nz.mem [1255] = \nz.mem_1255_sv2v_reg ;
  assign \nz.mem [1254] = \nz.mem_1254_sv2v_reg ;
  assign \nz.mem [1253] = \nz.mem_1253_sv2v_reg ;
  assign \nz.mem [1252] = \nz.mem_1252_sv2v_reg ;
  assign \nz.mem [1251] = \nz.mem_1251_sv2v_reg ;
  assign \nz.mem [1250] = \nz.mem_1250_sv2v_reg ;
  assign \nz.mem [1249] = \nz.mem_1249_sv2v_reg ;
  assign \nz.mem [1248] = \nz.mem_1248_sv2v_reg ;
  assign \nz.mem [1247] = \nz.mem_1247_sv2v_reg ;
  assign \nz.mem [1246] = \nz.mem_1246_sv2v_reg ;
  assign \nz.mem [1245] = \nz.mem_1245_sv2v_reg ;
  assign \nz.mem [1244] = \nz.mem_1244_sv2v_reg ;
  assign \nz.mem [1243] = \nz.mem_1243_sv2v_reg ;
  assign \nz.mem [1242] = \nz.mem_1242_sv2v_reg ;
  assign \nz.mem [1241] = \nz.mem_1241_sv2v_reg ;
  assign \nz.mem [1240] = \nz.mem_1240_sv2v_reg ;
  assign \nz.mem [1239] = \nz.mem_1239_sv2v_reg ;
  assign \nz.mem [1238] = \nz.mem_1238_sv2v_reg ;
  assign \nz.mem [1237] = \nz.mem_1237_sv2v_reg ;
  assign \nz.mem [1236] = \nz.mem_1236_sv2v_reg ;
  assign \nz.mem [1235] = \nz.mem_1235_sv2v_reg ;
  assign \nz.mem [1234] = \nz.mem_1234_sv2v_reg ;
  assign \nz.mem [1233] = \nz.mem_1233_sv2v_reg ;
  assign \nz.mem [1232] = \nz.mem_1232_sv2v_reg ;
  assign \nz.mem [1231] = \nz.mem_1231_sv2v_reg ;
  assign \nz.mem [1230] = \nz.mem_1230_sv2v_reg ;
  assign \nz.mem [1229] = \nz.mem_1229_sv2v_reg ;
  assign \nz.mem [1228] = \nz.mem_1228_sv2v_reg ;
  assign \nz.mem [1227] = \nz.mem_1227_sv2v_reg ;
  assign \nz.mem [1226] = \nz.mem_1226_sv2v_reg ;
  assign \nz.mem [1225] = \nz.mem_1225_sv2v_reg ;
  assign \nz.mem [1224] = \nz.mem_1224_sv2v_reg ;
  assign \nz.mem [1223] = \nz.mem_1223_sv2v_reg ;
  assign \nz.mem [1222] = \nz.mem_1222_sv2v_reg ;
  assign \nz.mem [1221] = \nz.mem_1221_sv2v_reg ;
  assign \nz.mem [1220] = \nz.mem_1220_sv2v_reg ;
  assign \nz.mem [1219] = \nz.mem_1219_sv2v_reg ;
  assign \nz.mem [1218] = \nz.mem_1218_sv2v_reg ;
  assign \nz.mem [1217] = \nz.mem_1217_sv2v_reg ;
  assign \nz.mem [1216] = \nz.mem_1216_sv2v_reg ;
  assign \nz.mem [1215] = \nz.mem_1215_sv2v_reg ;
  assign \nz.mem [1214] = \nz.mem_1214_sv2v_reg ;
  assign \nz.mem [1213] = \nz.mem_1213_sv2v_reg ;
  assign \nz.mem [1212] = \nz.mem_1212_sv2v_reg ;
  assign \nz.mem [1211] = \nz.mem_1211_sv2v_reg ;
  assign \nz.mem [1210] = \nz.mem_1210_sv2v_reg ;
  assign \nz.mem [1209] = \nz.mem_1209_sv2v_reg ;
  assign \nz.mem [1208] = \nz.mem_1208_sv2v_reg ;
  assign \nz.mem [1207] = \nz.mem_1207_sv2v_reg ;
  assign \nz.mem [1206] = \nz.mem_1206_sv2v_reg ;
  assign \nz.mem [1205] = \nz.mem_1205_sv2v_reg ;
  assign \nz.mem [1204] = \nz.mem_1204_sv2v_reg ;
  assign \nz.mem [1203] = \nz.mem_1203_sv2v_reg ;
  assign \nz.mem [1202] = \nz.mem_1202_sv2v_reg ;
  assign \nz.mem [1201] = \nz.mem_1201_sv2v_reg ;
  assign \nz.mem [1200] = \nz.mem_1200_sv2v_reg ;
  assign \nz.mem [1199] = \nz.mem_1199_sv2v_reg ;
  assign \nz.mem [1198] = \nz.mem_1198_sv2v_reg ;
  assign \nz.mem [1197] = \nz.mem_1197_sv2v_reg ;
  assign \nz.mem [1196] = \nz.mem_1196_sv2v_reg ;
  assign \nz.mem [1195] = \nz.mem_1195_sv2v_reg ;
  assign \nz.mem [1194] = \nz.mem_1194_sv2v_reg ;
  assign \nz.mem [1193] = \nz.mem_1193_sv2v_reg ;
  assign \nz.mem [1192] = \nz.mem_1192_sv2v_reg ;
  assign \nz.mem [1191] = \nz.mem_1191_sv2v_reg ;
  assign \nz.mem [1190] = \nz.mem_1190_sv2v_reg ;
  assign \nz.mem [1189] = \nz.mem_1189_sv2v_reg ;
  assign \nz.mem [1188] = \nz.mem_1188_sv2v_reg ;
  assign \nz.mem [1187] = \nz.mem_1187_sv2v_reg ;
  assign \nz.mem [1186] = \nz.mem_1186_sv2v_reg ;
  assign \nz.mem [1185] = \nz.mem_1185_sv2v_reg ;
  assign \nz.mem [1184] = \nz.mem_1184_sv2v_reg ;
  assign \nz.mem [1183] = \nz.mem_1183_sv2v_reg ;
  assign \nz.mem [1182] = \nz.mem_1182_sv2v_reg ;
  assign \nz.mem [1181] = \nz.mem_1181_sv2v_reg ;
  assign \nz.mem [1180] = \nz.mem_1180_sv2v_reg ;
  assign \nz.mem [1179] = \nz.mem_1179_sv2v_reg ;
  assign \nz.mem [1178] = \nz.mem_1178_sv2v_reg ;
  assign \nz.mem [1177] = \nz.mem_1177_sv2v_reg ;
  assign \nz.mem [1176] = \nz.mem_1176_sv2v_reg ;
  assign \nz.mem [1175] = \nz.mem_1175_sv2v_reg ;
  assign \nz.mem [1174] = \nz.mem_1174_sv2v_reg ;
  assign \nz.mem [1173] = \nz.mem_1173_sv2v_reg ;
  assign \nz.mem [1172] = \nz.mem_1172_sv2v_reg ;
  assign \nz.mem [1171] = \nz.mem_1171_sv2v_reg ;
  assign \nz.mem [1170] = \nz.mem_1170_sv2v_reg ;
  assign \nz.mem [1169] = \nz.mem_1169_sv2v_reg ;
  assign \nz.mem [1168] = \nz.mem_1168_sv2v_reg ;
  assign \nz.mem [1167] = \nz.mem_1167_sv2v_reg ;
  assign \nz.mem [1166] = \nz.mem_1166_sv2v_reg ;
  assign \nz.mem [1165] = \nz.mem_1165_sv2v_reg ;
  assign \nz.mem [1164] = \nz.mem_1164_sv2v_reg ;
  assign \nz.mem [1163] = \nz.mem_1163_sv2v_reg ;
  assign \nz.mem [1162] = \nz.mem_1162_sv2v_reg ;
  assign \nz.mem [1161] = \nz.mem_1161_sv2v_reg ;
  assign \nz.mem [1160] = \nz.mem_1160_sv2v_reg ;
  assign \nz.mem [1159] = \nz.mem_1159_sv2v_reg ;
  assign \nz.mem [1158] = \nz.mem_1158_sv2v_reg ;
  assign \nz.mem [1157] = \nz.mem_1157_sv2v_reg ;
  assign \nz.mem [1156] = \nz.mem_1156_sv2v_reg ;
  assign \nz.mem [1155] = \nz.mem_1155_sv2v_reg ;
  assign \nz.mem [1154] = \nz.mem_1154_sv2v_reg ;
  assign \nz.mem [1153] = \nz.mem_1153_sv2v_reg ;
  assign \nz.mem [1152] = \nz.mem_1152_sv2v_reg ;
  assign \nz.mem [1151] = \nz.mem_1151_sv2v_reg ;
  assign \nz.mem [1150] = \nz.mem_1150_sv2v_reg ;
  assign \nz.mem [1149] = \nz.mem_1149_sv2v_reg ;
  assign \nz.mem [1148] = \nz.mem_1148_sv2v_reg ;
  assign \nz.mem [1147] = \nz.mem_1147_sv2v_reg ;
  assign \nz.mem [1146] = \nz.mem_1146_sv2v_reg ;
  assign \nz.mem [1145] = \nz.mem_1145_sv2v_reg ;
  assign \nz.mem [1144] = \nz.mem_1144_sv2v_reg ;
  assign \nz.mem [1143] = \nz.mem_1143_sv2v_reg ;
  assign \nz.mem [1142] = \nz.mem_1142_sv2v_reg ;
  assign \nz.mem [1141] = \nz.mem_1141_sv2v_reg ;
  assign \nz.mem [1140] = \nz.mem_1140_sv2v_reg ;
  assign \nz.mem [1139] = \nz.mem_1139_sv2v_reg ;
  assign \nz.mem [1138] = \nz.mem_1138_sv2v_reg ;
  assign \nz.mem [1137] = \nz.mem_1137_sv2v_reg ;
  assign \nz.mem [1136] = \nz.mem_1136_sv2v_reg ;
  assign \nz.mem [1135] = \nz.mem_1135_sv2v_reg ;
  assign \nz.mem [1134] = \nz.mem_1134_sv2v_reg ;
  assign \nz.mem [1133] = \nz.mem_1133_sv2v_reg ;
  assign \nz.mem [1132] = \nz.mem_1132_sv2v_reg ;
  assign \nz.mem [1131] = \nz.mem_1131_sv2v_reg ;
  assign \nz.mem [1130] = \nz.mem_1130_sv2v_reg ;
  assign \nz.mem [1129] = \nz.mem_1129_sv2v_reg ;
  assign \nz.mem [1128] = \nz.mem_1128_sv2v_reg ;
  assign \nz.mem [1127] = \nz.mem_1127_sv2v_reg ;
  assign \nz.mem [1126] = \nz.mem_1126_sv2v_reg ;
  assign \nz.mem [1125] = \nz.mem_1125_sv2v_reg ;
  assign \nz.mem [1124] = \nz.mem_1124_sv2v_reg ;
  assign \nz.mem [1123] = \nz.mem_1123_sv2v_reg ;
  assign \nz.mem [1122] = \nz.mem_1122_sv2v_reg ;
  assign \nz.mem [1121] = \nz.mem_1121_sv2v_reg ;
  assign \nz.mem [1120] = \nz.mem_1120_sv2v_reg ;
  assign \nz.mem [1119] = \nz.mem_1119_sv2v_reg ;
  assign \nz.mem [1118] = \nz.mem_1118_sv2v_reg ;
  assign \nz.mem [1117] = \nz.mem_1117_sv2v_reg ;
  assign \nz.mem [1116] = \nz.mem_1116_sv2v_reg ;
  assign \nz.mem [1115] = \nz.mem_1115_sv2v_reg ;
  assign \nz.mem [1114] = \nz.mem_1114_sv2v_reg ;
  assign \nz.mem [1113] = \nz.mem_1113_sv2v_reg ;
  assign \nz.mem [1112] = \nz.mem_1112_sv2v_reg ;
  assign \nz.mem [1111] = \nz.mem_1111_sv2v_reg ;
  assign \nz.mem [1110] = \nz.mem_1110_sv2v_reg ;
  assign \nz.mem [1109] = \nz.mem_1109_sv2v_reg ;
  assign \nz.mem [1108] = \nz.mem_1108_sv2v_reg ;
  assign \nz.mem [1107] = \nz.mem_1107_sv2v_reg ;
  assign \nz.mem [1106] = \nz.mem_1106_sv2v_reg ;
  assign \nz.mem [1105] = \nz.mem_1105_sv2v_reg ;
  assign \nz.mem [1104] = \nz.mem_1104_sv2v_reg ;
  assign \nz.mem [1103] = \nz.mem_1103_sv2v_reg ;
  assign \nz.mem [1102] = \nz.mem_1102_sv2v_reg ;
  assign \nz.mem [1101] = \nz.mem_1101_sv2v_reg ;
  assign \nz.mem [1100] = \nz.mem_1100_sv2v_reg ;
  assign \nz.mem [1099] = \nz.mem_1099_sv2v_reg ;
  assign \nz.mem [1098] = \nz.mem_1098_sv2v_reg ;
  assign \nz.mem [1097] = \nz.mem_1097_sv2v_reg ;
  assign \nz.mem [1096] = \nz.mem_1096_sv2v_reg ;
  assign \nz.mem [1095] = \nz.mem_1095_sv2v_reg ;
  assign \nz.mem [1094] = \nz.mem_1094_sv2v_reg ;
  assign \nz.mem [1093] = \nz.mem_1093_sv2v_reg ;
  assign \nz.mem [1092] = \nz.mem_1092_sv2v_reg ;
  assign \nz.mem [1091] = \nz.mem_1091_sv2v_reg ;
  assign \nz.mem [1090] = \nz.mem_1090_sv2v_reg ;
  assign \nz.mem [1089] = \nz.mem_1089_sv2v_reg ;
  assign \nz.mem [1088] = \nz.mem_1088_sv2v_reg ;
  assign \nz.mem [1087] = \nz.mem_1087_sv2v_reg ;
  assign \nz.mem [1086] = \nz.mem_1086_sv2v_reg ;
  assign \nz.mem [1085] = \nz.mem_1085_sv2v_reg ;
  assign \nz.mem [1084] = \nz.mem_1084_sv2v_reg ;
  assign \nz.mem [1083] = \nz.mem_1083_sv2v_reg ;
  assign \nz.mem [1082] = \nz.mem_1082_sv2v_reg ;
  assign \nz.mem [1081] = \nz.mem_1081_sv2v_reg ;
  assign \nz.mem [1080] = \nz.mem_1080_sv2v_reg ;
  assign \nz.mem [1079] = \nz.mem_1079_sv2v_reg ;
  assign \nz.mem [1078] = \nz.mem_1078_sv2v_reg ;
  assign \nz.mem [1077] = \nz.mem_1077_sv2v_reg ;
  assign \nz.mem [1076] = \nz.mem_1076_sv2v_reg ;
  assign \nz.mem [1075] = \nz.mem_1075_sv2v_reg ;
  assign \nz.mem [1074] = \nz.mem_1074_sv2v_reg ;
  assign \nz.mem [1073] = \nz.mem_1073_sv2v_reg ;
  assign \nz.mem [1072] = \nz.mem_1072_sv2v_reg ;
  assign \nz.mem [1071] = \nz.mem_1071_sv2v_reg ;
  assign \nz.mem [1070] = \nz.mem_1070_sv2v_reg ;
  assign \nz.mem [1069] = \nz.mem_1069_sv2v_reg ;
  assign \nz.mem [1068] = \nz.mem_1068_sv2v_reg ;
  assign \nz.mem [1067] = \nz.mem_1067_sv2v_reg ;
  assign \nz.mem [1066] = \nz.mem_1066_sv2v_reg ;
  assign \nz.mem [1065] = \nz.mem_1065_sv2v_reg ;
  assign \nz.mem [1064] = \nz.mem_1064_sv2v_reg ;
  assign \nz.mem [1063] = \nz.mem_1063_sv2v_reg ;
  assign \nz.mem [1062] = \nz.mem_1062_sv2v_reg ;
  assign \nz.mem [1061] = \nz.mem_1061_sv2v_reg ;
  assign \nz.mem [1060] = \nz.mem_1060_sv2v_reg ;
  assign \nz.mem [1059] = \nz.mem_1059_sv2v_reg ;
  assign \nz.mem [1058] = \nz.mem_1058_sv2v_reg ;
  assign \nz.mem [1057] = \nz.mem_1057_sv2v_reg ;
  assign \nz.mem [1056] = \nz.mem_1056_sv2v_reg ;
  assign \nz.mem [1055] = \nz.mem_1055_sv2v_reg ;
  assign \nz.mem [1054] = \nz.mem_1054_sv2v_reg ;
  assign \nz.mem [1053] = \nz.mem_1053_sv2v_reg ;
  assign \nz.mem [1052] = \nz.mem_1052_sv2v_reg ;
  assign \nz.mem [1051] = \nz.mem_1051_sv2v_reg ;
  assign \nz.mem [1050] = \nz.mem_1050_sv2v_reg ;
  assign \nz.mem [1049] = \nz.mem_1049_sv2v_reg ;
  assign \nz.mem [1048] = \nz.mem_1048_sv2v_reg ;
  assign \nz.mem [1047] = \nz.mem_1047_sv2v_reg ;
  assign \nz.mem [1046] = \nz.mem_1046_sv2v_reg ;
  assign \nz.mem [1045] = \nz.mem_1045_sv2v_reg ;
  assign \nz.mem [1044] = \nz.mem_1044_sv2v_reg ;
  assign \nz.mem [1043] = \nz.mem_1043_sv2v_reg ;
  assign \nz.mem [1042] = \nz.mem_1042_sv2v_reg ;
  assign \nz.mem [1041] = \nz.mem_1041_sv2v_reg ;
  assign \nz.mem [1040] = \nz.mem_1040_sv2v_reg ;
  assign \nz.mem [1039] = \nz.mem_1039_sv2v_reg ;
  assign \nz.mem [1038] = \nz.mem_1038_sv2v_reg ;
  assign \nz.mem [1037] = \nz.mem_1037_sv2v_reg ;
  assign \nz.mem [1036] = \nz.mem_1036_sv2v_reg ;
  assign \nz.mem [1035] = \nz.mem_1035_sv2v_reg ;
  assign \nz.mem [1034] = \nz.mem_1034_sv2v_reg ;
  assign \nz.mem [1033] = \nz.mem_1033_sv2v_reg ;
  assign \nz.mem [1032] = \nz.mem_1032_sv2v_reg ;
  assign \nz.mem [1031] = \nz.mem_1031_sv2v_reg ;
  assign \nz.mem [1030] = \nz.mem_1030_sv2v_reg ;
  assign \nz.mem [1029] = \nz.mem_1029_sv2v_reg ;
  assign \nz.mem [1028] = \nz.mem_1028_sv2v_reg ;
  assign \nz.mem [1027] = \nz.mem_1027_sv2v_reg ;
  assign \nz.mem [1026] = \nz.mem_1026_sv2v_reg ;
  assign \nz.mem [1025] = \nz.mem_1025_sv2v_reg ;
  assign \nz.mem [1024] = \nz.mem_1024_sv2v_reg ;
  assign \nz.mem [1023] = \nz.mem_1023_sv2v_reg ;
  assign \nz.mem [1022] = \nz.mem_1022_sv2v_reg ;
  assign \nz.mem [1021] = \nz.mem_1021_sv2v_reg ;
  assign \nz.mem [1020] = \nz.mem_1020_sv2v_reg ;
  assign \nz.mem [1019] = \nz.mem_1019_sv2v_reg ;
  assign \nz.mem [1018] = \nz.mem_1018_sv2v_reg ;
  assign \nz.mem [1017] = \nz.mem_1017_sv2v_reg ;
  assign \nz.mem [1016] = \nz.mem_1016_sv2v_reg ;
  assign \nz.mem [1015] = \nz.mem_1015_sv2v_reg ;
  assign \nz.mem [1014] = \nz.mem_1014_sv2v_reg ;
  assign \nz.mem [1013] = \nz.mem_1013_sv2v_reg ;
  assign \nz.mem [1012] = \nz.mem_1012_sv2v_reg ;
  assign \nz.mem [1011] = \nz.mem_1011_sv2v_reg ;
  assign \nz.mem [1010] = \nz.mem_1010_sv2v_reg ;
  assign \nz.mem [1009] = \nz.mem_1009_sv2v_reg ;
  assign \nz.mem [1008] = \nz.mem_1008_sv2v_reg ;
  assign \nz.mem [1007] = \nz.mem_1007_sv2v_reg ;
  assign \nz.mem [1006] = \nz.mem_1006_sv2v_reg ;
  assign \nz.mem [1005] = \nz.mem_1005_sv2v_reg ;
  assign \nz.mem [1004] = \nz.mem_1004_sv2v_reg ;
  assign \nz.mem [1003] = \nz.mem_1003_sv2v_reg ;
  assign \nz.mem [1002] = \nz.mem_1002_sv2v_reg ;
  assign \nz.mem [1001] = \nz.mem_1001_sv2v_reg ;
  assign \nz.mem [1000] = \nz.mem_1000_sv2v_reg ;
  assign \nz.mem [999] = \nz.mem_999_sv2v_reg ;
  assign \nz.mem [998] = \nz.mem_998_sv2v_reg ;
  assign \nz.mem [997] = \nz.mem_997_sv2v_reg ;
  assign \nz.mem [996] = \nz.mem_996_sv2v_reg ;
  assign \nz.mem [995] = \nz.mem_995_sv2v_reg ;
  assign \nz.mem [994] = \nz.mem_994_sv2v_reg ;
  assign \nz.mem [993] = \nz.mem_993_sv2v_reg ;
  assign \nz.mem [992] = \nz.mem_992_sv2v_reg ;
  assign \nz.mem [991] = \nz.mem_991_sv2v_reg ;
  assign \nz.mem [990] = \nz.mem_990_sv2v_reg ;
  assign \nz.mem [989] = \nz.mem_989_sv2v_reg ;
  assign \nz.mem [988] = \nz.mem_988_sv2v_reg ;
  assign \nz.mem [987] = \nz.mem_987_sv2v_reg ;
  assign \nz.mem [986] = \nz.mem_986_sv2v_reg ;
  assign \nz.mem [985] = \nz.mem_985_sv2v_reg ;
  assign \nz.mem [984] = \nz.mem_984_sv2v_reg ;
  assign \nz.mem [983] = \nz.mem_983_sv2v_reg ;
  assign \nz.mem [982] = \nz.mem_982_sv2v_reg ;
  assign \nz.mem [981] = \nz.mem_981_sv2v_reg ;
  assign \nz.mem [980] = \nz.mem_980_sv2v_reg ;
  assign \nz.mem [979] = \nz.mem_979_sv2v_reg ;
  assign \nz.mem [978] = \nz.mem_978_sv2v_reg ;
  assign \nz.mem [977] = \nz.mem_977_sv2v_reg ;
  assign \nz.mem [976] = \nz.mem_976_sv2v_reg ;
  assign \nz.mem [975] = \nz.mem_975_sv2v_reg ;
  assign \nz.mem [974] = \nz.mem_974_sv2v_reg ;
  assign \nz.mem [973] = \nz.mem_973_sv2v_reg ;
  assign \nz.mem [972] = \nz.mem_972_sv2v_reg ;
  assign \nz.mem [971] = \nz.mem_971_sv2v_reg ;
  assign \nz.mem [970] = \nz.mem_970_sv2v_reg ;
  assign \nz.mem [969] = \nz.mem_969_sv2v_reg ;
  assign \nz.mem [968] = \nz.mem_968_sv2v_reg ;
  assign \nz.mem [967] = \nz.mem_967_sv2v_reg ;
  assign \nz.mem [966] = \nz.mem_966_sv2v_reg ;
  assign \nz.mem [965] = \nz.mem_965_sv2v_reg ;
  assign \nz.mem [964] = \nz.mem_964_sv2v_reg ;
  assign \nz.mem [963] = \nz.mem_963_sv2v_reg ;
  assign \nz.mem [962] = \nz.mem_962_sv2v_reg ;
  assign \nz.mem [961] = \nz.mem_961_sv2v_reg ;
  assign \nz.mem [960] = \nz.mem_960_sv2v_reg ;
  assign \nz.mem [959] = \nz.mem_959_sv2v_reg ;
  assign \nz.mem [958] = \nz.mem_958_sv2v_reg ;
  assign \nz.mem [957] = \nz.mem_957_sv2v_reg ;
  assign \nz.mem [956] = \nz.mem_956_sv2v_reg ;
  assign \nz.mem [955] = \nz.mem_955_sv2v_reg ;
  assign \nz.mem [954] = \nz.mem_954_sv2v_reg ;
  assign \nz.mem [953] = \nz.mem_953_sv2v_reg ;
  assign \nz.mem [952] = \nz.mem_952_sv2v_reg ;
  assign \nz.mem [951] = \nz.mem_951_sv2v_reg ;
  assign \nz.mem [950] = \nz.mem_950_sv2v_reg ;
  assign \nz.mem [949] = \nz.mem_949_sv2v_reg ;
  assign \nz.mem [948] = \nz.mem_948_sv2v_reg ;
  assign \nz.mem [947] = \nz.mem_947_sv2v_reg ;
  assign \nz.mem [946] = \nz.mem_946_sv2v_reg ;
  assign \nz.mem [945] = \nz.mem_945_sv2v_reg ;
  assign \nz.mem [944] = \nz.mem_944_sv2v_reg ;
  assign \nz.mem [943] = \nz.mem_943_sv2v_reg ;
  assign \nz.mem [942] = \nz.mem_942_sv2v_reg ;
  assign \nz.mem [941] = \nz.mem_941_sv2v_reg ;
  assign \nz.mem [940] = \nz.mem_940_sv2v_reg ;
  assign \nz.mem [939] = \nz.mem_939_sv2v_reg ;
  assign \nz.mem [938] = \nz.mem_938_sv2v_reg ;
  assign \nz.mem [937] = \nz.mem_937_sv2v_reg ;
  assign \nz.mem [936] = \nz.mem_936_sv2v_reg ;
  assign \nz.mem [935] = \nz.mem_935_sv2v_reg ;
  assign \nz.mem [934] = \nz.mem_934_sv2v_reg ;
  assign \nz.mem [933] = \nz.mem_933_sv2v_reg ;
  assign \nz.mem [932] = \nz.mem_932_sv2v_reg ;
  assign \nz.mem [931] = \nz.mem_931_sv2v_reg ;
  assign \nz.mem [930] = \nz.mem_930_sv2v_reg ;
  assign \nz.mem [929] = \nz.mem_929_sv2v_reg ;
  assign \nz.mem [928] = \nz.mem_928_sv2v_reg ;
  assign \nz.mem [927] = \nz.mem_927_sv2v_reg ;
  assign \nz.mem [926] = \nz.mem_926_sv2v_reg ;
  assign \nz.mem [925] = \nz.mem_925_sv2v_reg ;
  assign \nz.mem [924] = \nz.mem_924_sv2v_reg ;
  assign \nz.mem [923] = \nz.mem_923_sv2v_reg ;
  assign \nz.mem [922] = \nz.mem_922_sv2v_reg ;
  assign \nz.mem [921] = \nz.mem_921_sv2v_reg ;
  assign \nz.mem [920] = \nz.mem_920_sv2v_reg ;
  assign \nz.mem [919] = \nz.mem_919_sv2v_reg ;
  assign \nz.mem [918] = \nz.mem_918_sv2v_reg ;
  assign \nz.mem [917] = \nz.mem_917_sv2v_reg ;
  assign \nz.mem [916] = \nz.mem_916_sv2v_reg ;
  assign \nz.mem [915] = \nz.mem_915_sv2v_reg ;
  assign \nz.mem [914] = \nz.mem_914_sv2v_reg ;
  assign \nz.mem [913] = \nz.mem_913_sv2v_reg ;
  assign \nz.mem [912] = \nz.mem_912_sv2v_reg ;
  assign \nz.mem [911] = \nz.mem_911_sv2v_reg ;
  assign \nz.mem [910] = \nz.mem_910_sv2v_reg ;
  assign \nz.mem [909] = \nz.mem_909_sv2v_reg ;
  assign \nz.mem [908] = \nz.mem_908_sv2v_reg ;
  assign \nz.mem [907] = \nz.mem_907_sv2v_reg ;
  assign \nz.mem [906] = \nz.mem_906_sv2v_reg ;
  assign \nz.mem [905] = \nz.mem_905_sv2v_reg ;
  assign \nz.mem [904] = \nz.mem_904_sv2v_reg ;
  assign \nz.mem [903] = \nz.mem_903_sv2v_reg ;
  assign \nz.mem [902] = \nz.mem_902_sv2v_reg ;
  assign \nz.mem [901] = \nz.mem_901_sv2v_reg ;
  assign \nz.mem [900] = \nz.mem_900_sv2v_reg ;
  assign \nz.mem [899] = \nz.mem_899_sv2v_reg ;
  assign \nz.mem [898] = \nz.mem_898_sv2v_reg ;
  assign \nz.mem [897] = \nz.mem_897_sv2v_reg ;
  assign \nz.mem [896] = \nz.mem_896_sv2v_reg ;
  assign \nz.mem [895] = \nz.mem_895_sv2v_reg ;
  assign \nz.mem [894] = \nz.mem_894_sv2v_reg ;
  assign \nz.mem [893] = \nz.mem_893_sv2v_reg ;
  assign \nz.mem [892] = \nz.mem_892_sv2v_reg ;
  assign \nz.mem [891] = \nz.mem_891_sv2v_reg ;
  assign \nz.mem [890] = \nz.mem_890_sv2v_reg ;
  assign \nz.mem [889] = \nz.mem_889_sv2v_reg ;
  assign \nz.mem [888] = \nz.mem_888_sv2v_reg ;
  assign \nz.mem [887] = \nz.mem_887_sv2v_reg ;
  assign \nz.mem [886] = \nz.mem_886_sv2v_reg ;
  assign \nz.mem [885] = \nz.mem_885_sv2v_reg ;
  assign \nz.mem [884] = \nz.mem_884_sv2v_reg ;
  assign \nz.mem [883] = \nz.mem_883_sv2v_reg ;
  assign \nz.mem [882] = \nz.mem_882_sv2v_reg ;
  assign \nz.mem [881] = \nz.mem_881_sv2v_reg ;
  assign \nz.mem [880] = \nz.mem_880_sv2v_reg ;
  assign \nz.mem [879] = \nz.mem_879_sv2v_reg ;
  assign \nz.mem [878] = \nz.mem_878_sv2v_reg ;
  assign \nz.mem [877] = \nz.mem_877_sv2v_reg ;
  assign \nz.mem [876] = \nz.mem_876_sv2v_reg ;
  assign \nz.mem [875] = \nz.mem_875_sv2v_reg ;
  assign \nz.mem [874] = \nz.mem_874_sv2v_reg ;
  assign \nz.mem [873] = \nz.mem_873_sv2v_reg ;
  assign \nz.mem [872] = \nz.mem_872_sv2v_reg ;
  assign \nz.mem [871] = \nz.mem_871_sv2v_reg ;
  assign \nz.mem [870] = \nz.mem_870_sv2v_reg ;
  assign \nz.mem [869] = \nz.mem_869_sv2v_reg ;
  assign \nz.mem [868] = \nz.mem_868_sv2v_reg ;
  assign \nz.mem [867] = \nz.mem_867_sv2v_reg ;
  assign \nz.mem [866] = \nz.mem_866_sv2v_reg ;
  assign \nz.mem [865] = \nz.mem_865_sv2v_reg ;
  assign \nz.mem [864] = \nz.mem_864_sv2v_reg ;
  assign \nz.mem [863] = \nz.mem_863_sv2v_reg ;
  assign \nz.mem [862] = \nz.mem_862_sv2v_reg ;
  assign \nz.mem [861] = \nz.mem_861_sv2v_reg ;
  assign \nz.mem [860] = \nz.mem_860_sv2v_reg ;
  assign \nz.mem [859] = \nz.mem_859_sv2v_reg ;
  assign \nz.mem [858] = \nz.mem_858_sv2v_reg ;
  assign \nz.mem [857] = \nz.mem_857_sv2v_reg ;
  assign \nz.mem [856] = \nz.mem_856_sv2v_reg ;
  assign \nz.mem [855] = \nz.mem_855_sv2v_reg ;
  assign \nz.mem [854] = \nz.mem_854_sv2v_reg ;
  assign \nz.mem [853] = \nz.mem_853_sv2v_reg ;
  assign \nz.mem [852] = \nz.mem_852_sv2v_reg ;
  assign \nz.mem [851] = \nz.mem_851_sv2v_reg ;
  assign \nz.mem [850] = \nz.mem_850_sv2v_reg ;
  assign \nz.mem [849] = \nz.mem_849_sv2v_reg ;
  assign \nz.mem [848] = \nz.mem_848_sv2v_reg ;
  assign \nz.mem [847] = \nz.mem_847_sv2v_reg ;
  assign \nz.mem [846] = \nz.mem_846_sv2v_reg ;
  assign \nz.mem [845] = \nz.mem_845_sv2v_reg ;
  assign \nz.mem [844] = \nz.mem_844_sv2v_reg ;
  assign \nz.mem [843] = \nz.mem_843_sv2v_reg ;
  assign \nz.mem [842] = \nz.mem_842_sv2v_reg ;
  assign \nz.mem [841] = \nz.mem_841_sv2v_reg ;
  assign \nz.mem [840] = \nz.mem_840_sv2v_reg ;
  assign \nz.mem [839] = \nz.mem_839_sv2v_reg ;
  assign \nz.mem [838] = \nz.mem_838_sv2v_reg ;
  assign \nz.mem [837] = \nz.mem_837_sv2v_reg ;
  assign \nz.mem [836] = \nz.mem_836_sv2v_reg ;
  assign \nz.mem [835] = \nz.mem_835_sv2v_reg ;
  assign \nz.mem [834] = \nz.mem_834_sv2v_reg ;
  assign \nz.mem [833] = \nz.mem_833_sv2v_reg ;
  assign \nz.mem [832] = \nz.mem_832_sv2v_reg ;
  assign \nz.mem [831] = \nz.mem_831_sv2v_reg ;
  assign \nz.mem [830] = \nz.mem_830_sv2v_reg ;
  assign \nz.mem [829] = \nz.mem_829_sv2v_reg ;
  assign \nz.mem [828] = \nz.mem_828_sv2v_reg ;
  assign \nz.mem [827] = \nz.mem_827_sv2v_reg ;
  assign \nz.mem [826] = \nz.mem_826_sv2v_reg ;
  assign \nz.mem [825] = \nz.mem_825_sv2v_reg ;
  assign \nz.mem [824] = \nz.mem_824_sv2v_reg ;
  assign \nz.mem [823] = \nz.mem_823_sv2v_reg ;
  assign \nz.mem [822] = \nz.mem_822_sv2v_reg ;
  assign \nz.mem [821] = \nz.mem_821_sv2v_reg ;
  assign \nz.mem [820] = \nz.mem_820_sv2v_reg ;
  assign \nz.mem [819] = \nz.mem_819_sv2v_reg ;
  assign \nz.mem [818] = \nz.mem_818_sv2v_reg ;
  assign \nz.mem [817] = \nz.mem_817_sv2v_reg ;
  assign \nz.mem [816] = \nz.mem_816_sv2v_reg ;
  assign \nz.mem [815] = \nz.mem_815_sv2v_reg ;
  assign \nz.mem [814] = \nz.mem_814_sv2v_reg ;
  assign \nz.mem [813] = \nz.mem_813_sv2v_reg ;
  assign \nz.mem [812] = \nz.mem_812_sv2v_reg ;
  assign \nz.mem [811] = \nz.mem_811_sv2v_reg ;
  assign \nz.mem [810] = \nz.mem_810_sv2v_reg ;
  assign \nz.mem [809] = \nz.mem_809_sv2v_reg ;
  assign \nz.mem [808] = \nz.mem_808_sv2v_reg ;
  assign \nz.mem [807] = \nz.mem_807_sv2v_reg ;
  assign \nz.mem [806] = \nz.mem_806_sv2v_reg ;
  assign \nz.mem [805] = \nz.mem_805_sv2v_reg ;
  assign \nz.mem [804] = \nz.mem_804_sv2v_reg ;
  assign \nz.mem [803] = \nz.mem_803_sv2v_reg ;
  assign \nz.mem [802] = \nz.mem_802_sv2v_reg ;
  assign \nz.mem [801] = \nz.mem_801_sv2v_reg ;
  assign \nz.mem [800] = \nz.mem_800_sv2v_reg ;
  assign \nz.mem [799] = \nz.mem_799_sv2v_reg ;
  assign \nz.mem [798] = \nz.mem_798_sv2v_reg ;
  assign \nz.mem [797] = \nz.mem_797_sv2v_reg ;
  assign \nz.mem [796] = \nz.mem_796_sv2v_reg ;
  assign \nz.mem [795] = \nz.mem_795_sv2v_reg ;
  assign \nz.mem [794] = \nz.mem_794_sv2v_reg ;
  assign \nz.mem [793] = \nz.mem_793_sv2v_reg ;
  assign \nz.mem [792] = \nz.mem_792_sv2v_reg ;
  assign \nz.mem [791] = \nz.mem_791_sv2v_reg ;
  assign \nz.mem [790] = \nz.mem_790_sv2v_reg ;
  assign \nz.mem [789] = \nz.mem_789_sv2v_reg ;
  assign \nz.mem [788] = \nz.mem_788_sv2v_reg ;
  assign \nz.mem [787] = \nz.mem_787_sv2v_reg ;
  assign \nz.mem [786] = \nz.mem_786_sv2v_reg ;
  assign \nz.mem [785] = \nz.mem_785_sv2v_reg ;
  assign \nz.mem [784] = \nz.mem_784_sv2v_reg ;
  assign \nz.mem [783] = \nz.mem_783_sv2v_reg ;
  assign \nz.mem [782] = \nz.mem_782_sv2v_reg ;
  assign \nz.mem [781] = \nz.mem_781_sv2v_reg ;
  assign \nz.mem [780] = \nz.mem_780_sv2v_reg ;
  assign \nz.mem [779] = \nz.mem_779_sv2v_reg ;
  assign \nz.mem [778] = \nz.mem_778_sv2v_reg ;
  assign \nz.mem [777] = \nz.mem_777_sv2v_reg ;
  assign \nz.mem [776] = \nz.mem_776_sv2v_reg ;
  assign \nz.mem [775] = \nz.mem_775_sv2v_reg ;
  assign \nz.mem [774] = \nz.mem_774_sv2v_reg ;
  assign \nz.mem [773] = \nz.mem_773_sv2v_reg ;
  assign \nz.mem [772] = \nz.mem_772_sv2v_reg ;
  assign \nz.mem [771] = \nz.mem_771_sv2v_reg ;
  assign \nz.mem [770] = \nz.mem_770_sv2v_reg ;
  assign \nz.mem [769] = \nz.mem_769_sv2v_reg ;
  assign \nz.mem [768] = \nz.mem_768_sv2v_reg ;
  assign \nz.mem [767] = \nz.mem_767_sv2v_reg ;
  assign \nz.mem [766] = \nz.mem_766_sv2v_reg ;
  assign \nz.mem [765] = \nz.mem_765_sv2v_reg ;
  assign \nz.mem [764] = \nz.mem_764_sv2v_reg ;
  assign \nz.mem [763] = \nz.mem_763_sv2v_reg ;
  assign \nz.mem [762] = \nz.mem_762_sv2v_reg ;
  assign \nz.mem [761] = \nz.mem_761_sv2v_reg ;
  assign \nz.mem [760] = \nz.mem_760_sv2v_reg ;
  assign \nz.mem [759] = \nz.mem_759_sv2v_reg ;
  assign \nz.mem [758] = \nz.mem_758_sv2v_reg ;
  assign \nz.mem [757] = \nz.mem_757_sv2v_reg ;
  assign \nz.mem [756] = \nz.mem_756_sv2v_reg ;
  assign \nz.mem [755] = \nz.mem_755_sv2v_reg ;
  assign \nz.mem [754] = \nz.mem_754_sv2v_reg ;
  assign \nz.mem [753] = \nz.mem_753_sv2v_reg ;
  assign \nz.mem [752] = \nz.mem_752_sv2v_reg ;
  assign \nz.mem [751] = \nz.mem_751_sv2v_reg ;
  assign \nz.mem [750] = \nz.mem_750_sv2v_reg ;
  assign \nz.mem [749] = \nz.mem_749_sv2v_reg ;
  assign \nz.mem [748] = \nz.mem_748_sv2v_reg ;
  assign \nz.mem [747] = \nz.mem_747_sv2v_reg ;
  assign \nz.mem [746] = \nz.mem_746_sv2v_reg ;
  assign \nz.mem [745] = \nz.mem_745_sv2v_reg ;
  assign \nz.mem [744] = \nz.mem_744_sv2v_reg ;
  assign \nz.mem [743] = \nz.mem_743_sv2v_reg ;
  assign \nz.mem [742] = \nz.mem_742_sv2v_reg ;
  assign \nz.mem [741] = \nz.mem_741_sv2v_reg ;
  assign \nz.mem [740] = \nz.mem_740_sv2v_reg ;
  assign \nz.mem [739] = \nz.mem_739_sv2v_reg ;
  assign \nz.mem [738] = \nz.mem_738_sv2v_reg ;
  assign \nz.mem [737] = \nz.mem_737_sv2v_reg ;
  assign \nz.mem [736] = \nz.mem_736_sv2v_reg ;
  assign \nz.mem [735] = \nz.mem_735_sv2v_reg ;
  assign \nz.mem [734] = \nz.mem_734_sv2v_reg ;
  assign \nz.mem [733] = \nz.mem_733_sv2v_reg ;
  assign \nz.mem [732] = \nz.mem_732_sv2v_reg ;
  assign \nz.mem [731] = \nz.mem_731_sv2v_reg ;
  assign \nz.mem [730] = \nz.mem_730_sv2v_reg ;
  assign \nz.mem [729] = \nz.mem_729_sv2v_reg ;
  assign \nz.mem [728] = \nz.mem_728_sv2v_reg ;
  assign \nz.mem [727] = \nz.mem_727_sv2v_reg ;
  assign \nz.mem [726] = \nz.mem_726_sv2v_reg ;
  assign \nz.mem [725] = \nz.mem_725_sv2v_reg ;
  assign \nz.mem [724] = \nz.mem_724_sv2v_reg ;
  assign \nz.mem [723] = \nz.mem_723_sv2v_reg ;
  assign \nz.mem [722] = \nz.mem_722_sv2v_reg ;
  assign \nz.mem [721] = \nz.mem_721_sv2v_reg ;
  assign \nz.mem [720] = \nz.mem_720_sv2v_reg ;
  assign \nz.mem [719] = \nz.mem_719_sv2v_reg ;
  assign \nz.mem [718] = \nz.mem_718_sv2v_reg ;
  assign \nz.mem [717] = \nz.mem_717_sv2v_reg ;
  assign \nz.mem [716] = \nz.mem_716_sv2v_reg ;
  assign \nz.mem [715] = \nz.mem_715_sv2v_reg ;
  assign \nz.mem [714] = \nz.mem_714_sv2v_reg ;
  assign \nz.mem [713] = \nz.mem_713_sv2v_reg ;
  assign \nz.mem [712] = \nz.mem_712_sv2v_reg ;
  assign \nz.mem [711] = \nz.mem_711_sv2v_reg ;
  assign \nz.mem [710] = \nz.mem_710_sv2v_reg ;
  assign \nz.mem [709] = \nz.mem_709_sv2v_reg ;
  assign \nz.mem [708] = \nz.mem_708_sv2v_reg ;
  assign \nz.mem [707] = \nz.mem_707_sv2v_reg ;
  assign \nz.mem [706] = \nz.mem_706_sv2v_reg ;
  assign \nz.mem [705] = \nz.mem_705_sv2v_reg ;
  assign \nz.mem [704] = \nz.mem_704_sv2v_reg ;
  assign \nz.mem [703] = \nz.mem_703_sv2v_reg ;
  assign \nz.mem [702] = \nz.mem_702_sv2v_reg ;
  assign \nz.mem [701] = \nz.mem_701_sv2v_reg ;
  assign \nz.mem [700] = \nz.mem_700_sv2v_reg ;
  assign \nz.mem [699] = \nz.mem_699_sv2v_reg ;
  assign \nz.mem [698] = \nz.mem_698_sv2v_reg ;
  assign \nz.mem [697] = \nz.mem_697_sv2v_reg ;
  assign \nz.mem [696] = \nz.mem_696_sv2v_reg ;
  assign \nz.mem [695] = \nz.mem_695_sv2v_reg ;
  assign \nz.mem [694] = \nz.mem_694_sv2v_reg ;
  assign \nz.mem [693] = \nz.mem_693_sv2v_reg ;
  assign \nz.mem [692] = \nz.mem_692_sv2v_reg ;
  assign \nz.mem [691] = \nz.mem_691_sv2v_reg ;
  assign \nz.mem [690] = \nz.mem_690_sv2v_reg ;
  assign \nz.mem [689] = \nz.mem_689_sv2v_reg ;
  assign \nz.mem [688] = \nz.mem_688_sv2v_reg ;
  assign \nz.mem [687] = \nz.mem_687_sv2v_reg ;
  assign \nz.mem [686] = \nz.mem_686_sv2v_reg ;
  assign \nz.mem [685] = \nz.mem_685_sv2v_reg ;
  assign \nz.mem [684] = \nz.mem_684_sv2v_reg ;
  assign \nz.mem [683] = \nz.mem_683_sv2v_reg ;
  assign \nz.mem [682] = \nz.mem_682_sv2v_reg ;
  assign \nz.mem [681] = \nz.mem_681_sv2v_reg ;
  assign \nz.mem [680] = \nz.mem_680_sv2v_reg ;
  assign \nz.mem [679] = \nz.mem_679_sv2v_reg ;
  assign \nz.mem [678] = \nz.mem_678_sv2v_reg ;
  assign \nz.mem [677] = \nz.mem_677_sv2v_reg ;
  assign \nz.mem [676] = \nz.mem_676_sv2v_reg ;
  assign \nz.mem [675] = \nz.mem_675_sv2v_reg ;
  assign \nz.mem [674] = \nz.mem_674_sv2v_reg ;
  assign \nz.mem [673] = \nz.mem_673_sv2v_reg ;
  assign \nz.mem [672] = \nz.mem_672_sv2v_reg ;
  assign \nz.mem [671] = \nz.mem_671_sv2v_reg ;
  assign \nz.mem [670] = \nz.mem_670_sv2v_reg ;
  assign \nz.mem [669] = \nz.mem_669_sv2v_reg ;
  assign \nz.mem [668] = \nz.mem_668_sv2v_reg ;
  assign \nz.mem [667] = \nz.mem_667_sv2v_reg ;
  assign \nz.mem [666] = \nz.mem_666_sv2v_reg ;
  assign \nz.mem [665] = \nz.mem_665_sv2v_reg ;
  assign \nz.mem [664] = \nz.mem_664_sv2v_reg ;
  assign \nz.mem [663] = \nz.mem_663_sv2v_reg ;
  assign \nz.mem [662] = \nz.mem_662_sv2v_reg ;
  assign \nz.mem [661] = \nz.mem_661_sv2v_reg ;
  assign \nz.mem [660] = \nz.mem_660_sv2v_reg ;
  assign \nz.mem [659] = \nz.mem_659_sv2v_reg ;
  assign \nz.mem [658] = \nz.mem_658_sv2v_reg ;
  assign \nz.mem [657] = \nz.mem_657_sv2v_reg ;
  assign \nz.mem [656] = \nz.mem_656_sv2v_reg ;
  assign \nz.mem [655] = \nz.mem_655_sv2v_reg ;
  assign \nz.mem [654] = \nz.mem_654_sv2v_reg ;
  assign \nz.mem [653] = \nz.mem_653_sv2v_reg ;
  assign \nz.mem [652] = \nz.mem_652_sv2v_reg ;
  assign \nz.mem [651] = \nz.mem_651_sv2v_reg ;
  assign \nz.mem [650] = \nz.mem_650_sv2v_reg ;
  assign \nz.mem [649] = \nz.mem_649_sv2v_reg ;
  assign \nz.mem [648] = \nz.mem_648_sv2v_reg ;
  assign \nz.mem [647] = \nz.mem_647_sv2v_reg ;
  assign \nz.mem [646] = \nz.mem_646_sv2v_reg ;
  assign \nz.mem [645] = \nz.mem_645_sv2v_reg ;
  assign \nz.mem [644] = \nz.mem_644_sv2v_reg ;
  assign \nz.mem [643] = \nz.mem_643_sv2v_reg ;
  assign \nz.mem [642] = \nz.mem_642_sv2v_reg ;
  assign \nz.mem [641] = \nz.mem_641_sv2v_reg ;
  assign \nz.mem [640] = \nz.mem_640_sv2v_reg ;
  assign \nz.mem [639] = \nz.mem_639_sv2v_reg ;
  assign \nz.mem [638] = \nz.mem_638_sv2v_reg ;
  assign \nz.mem [637] = \nz.mem_637_sv2v_reg ;
  assign \nz.mem [636] = \nz.mem_636_sv2v_reg ;
  assign \nz.mem [635] = \nz.mem_635_sv2v_reg ;
  assign \nz.mem [634] = \nz.mem_634_sv2v_reg ;
  assign \nz.mem [633] = \nz.mem_633_sv2v_reg ;
  assign \nz.mem [632] = \nz.mem_632_sv2v_reg ;
  assign \nz.mem [631] = \nz.mem_631_sv2v_reg ;
  assign \nz.mem [630] = \nz.mem_630_sv2v_reg ;
  assign \nz.mem [629] = \nz.mem_629_sv2v_reg ;
  assign \nz.mem [628] = \nz.mem_628_sv2v_reg ;
  assign \nz.mem [627] = \nz.mem_627_sv2v_reg ;
  assign \nz.mem [626] = \nz.mem_626_sv2v_reg ;
  assign \nz.mem [625] = \nz.mem_625_sv2v_reg ;
  assign \nz.mem [624] = \nz.mem_624_sv2v_reg ;
  assign \nz.mem [623] = \nz.mem_623_sv2v_reg ;
  assign \nz.mem [622] = \nz.mem_622_sv2v_reg ;
  assign \nz.mem [621] = \nz.mem_621_sv2v_reg ;
  assign \nz.mem [620] = \nz.mem_620_sv2v_reg ;
  assign \nz.mem [619] = \nz.mem_619_sv2v_reg ;
  assign \nz.mem [618] = \nz.mem_618_sv2v_reg ;
  assign \nz.mem [617] = \nz.mem_617_sv2v_reg ;
  assign \nz.mem [616] = \nz.mem_616_sv2v_reg ;
  assign \nz.mem [615] = \nz.mem_615_sv2v_reg ;
  assign \nz.mem [614] = \nz.mem_614_sv2v_reg ;
  assign \nz.mem [613] = \nz.mem_613_sv2v_reg ;
  assign \nz.mem [612] = \nz.mem_612_sv2v_reg ;
  assign \nz.mem [611] = \nz.mem_611_sv2v_reg ;
  assign \nz.mem [610] = \nz.mem_610_sv2v_reg ;
  assign \nz.mem [609] = \nz.mem_609_sv2v_reg ;
  assign \nz.mem [608] = \nz.mem_608_sv2v_reg ;
  assign \nz.mem [607] = \nz.mem_607_sv2v_reg ;
  assign \nz.mem [606] = \nz.mem_606_sv2v_reg ;
  assign \nz.mem [605] = \nz.mem_605_sv2v_reg ;
  assign \nz.mem [604] = \nz.mem_604_sv2v_reg ;
  assign \nz.mem [603] = \nz.mem_603_sv2v_reg ;
  assign \nz.mem [602] = \nz.mem_602_sv2v_reg ;
  assign \nz.mem [601] = \nz.mem_601_sv2v_reg ;
  assign \nz.mem [600] = \nz.mem_600_sv2v_reg ;
  assign \nz.mem [599] = \nz.mem_599_sv2v_reg ;
  assign \nz.mem [598] = \nz.mem_598_sv2v_reg ;
  assign \nz.mem [597] = \nz.mem_597_sv2v_reg ;
  assign \nz.mem [596] = \nz.mem_596_sv2v_reg ;
  assign \nz.mem [595] = \nz.mem_595_sv2v_reg ;
  assign \nz.mem [594] = \nz.mem_594_sv2v_reg ;
  assign \nz.mem [593] = \nz.mem_593_sv2v_reg ;
  assign \nz.mem [592] = \nz.mem_592_sv2v_reg ;
  assign \nz.mem [591] = \nz.mem_591_sv2v_reg ;
  assign \nz.mem [590] = \nz.mem_590_sv2v_reg ;
  assign \nz.mem [589] = \nz.mem_589_sv2v_reg ;
  assign \nz.mem [588] = \nz.mem_588_sv2v_reg ;
  assign \nz.mem [587] = \nz.mem_587_sv2v_reg ;
  assign \nz.mem [586] = \nz.mem_586_sv2v_reg ;
  assign \nz.mem [585] = \nz.mem_585_sv2v_reg ;
  assign \nz.mem [584] = \nz.mem_584_sv2v_reg ;
  assign \nz.mem [583] = \nz.mem_583_sv2v_reg ;
  assign \nz.mem [582] = \nz.mem_582_sv2v_reg ;
  assign \nz.mem [581] = \nz.mem_581_sv2v_reg ;
  assign \nz.mem [580] = \nz.mem_580_sv2v_reg ;
  assign \nz.mem [579] = \nz.mem_579_sv2v_reg ;
  assign \nz.mem [578] = \nz.mem_578_sv2v_reg ;
  assign \nz.mem [577] = \nz.mem_577_sv2v_reg ;
  assign \nz.mem [576] = \nz.mem_576_sv2v_reg ;
  assign \nz.mem [575] = \nz.mem_575_sv2v_reg ;
  assign \nz.mem [574] = \nz.mem_574_sv2v_reg ;
  assign \nz.mem [573] = \nz.mem_573_sv2v_reg ;
  assign \nz.mem [572] = \nz.mem_572_sv2v_reg ;
  assign \nz.mem [571] = \nz.mem_571_sv2v_reg ;
  assign \nz.mem [570] = \nz.mem_570_sv2v_reg ;
  assign \nz.mem [569] = \nz.mem_569_sv2v_reg ;
  assign \nz.mem [568] = \nz.mem_568_sv2v_reg ;
  assign \nz.mem [567] = \nz.mem_567_sv2v_reg ;
  assign \nz.mem [566] = \nz.mem_566_sv2v_reg ;
  assign \nz.mem [565] = \nz.mem_565_sv2v_reg ;
  assign \nz.mem [564] = \nz.mem_564_sv2v_reg ;
  assign \nz.mem [563] = \nz.mem_563_sv2v_reg ;
  assign \nz.mem [562] = \nz.mem_562_sv2v_reg ;
  assign \nz.mem [561] = \nz.mem_561_sv2v_reg ;
  assign \nz.mem [560] = \nz.mem_560_sv2v_reg ;
  assign \nz.mem [559] = \nz.mem_559_sv2v_reg ;
  assign \nz.mem [558] = \nz.mem_558_sv2v_reg ;
  assign \nz.mem [557] = \nz.mem_557_sv2v_reg ;
  assign \nz.mem [556] = \nz.mem_556_sv2v_reg ;
  assign \nz.mem [555] = \nz.mem_555_sv2v_reg ;
  assign \nz.mem [554] = \nz.mem_554_sv2v_reg ;
  assign \nz.mem [553] = \nz.mem_553_sv2v_reg ;
  assign \nz.mem [552] = \nz.mem_552_sv2v_reg ;
  assign \nz.mem [551] = \nz.mem_551_sv2v_reg ;
  assign \nz.mem [550] = \nz.mem_550_sv2v_reg ;
  assign \nz.mem [549] = \nz.mem_549_sv2v_reg ;
  assign \nz.mem [548] = \nz.mem_548_sv2v_reg ;
  assign \nz.mem [547] = \nz.mem_547_sv2v_reg ;
  assign \nz.mem [546] = \nz.mem_546_sv2v_reg ;
  assign \nz.mem [545] = \nz.mem_545_sv2v_reg ;
  assign \nz.mem [544] = \nz.mem_544_sv2v_reg ;
  assign \nz.mem [543] = \nz.mem_543_sv2v_reg ;
  assign \nz.mem [542] = \nz.mem_542_sv2v_reg ;
  assign \nz.mem [541] = \nz.mem_541_sv2v_reg ;
  assign \nz.mem [540] = \nz.mem_540_sv2v_reg ;
  assign \nz.mem [539] = \nz.mem_539_sv2v_reg ;
  assign \nz.mem [538] = \nz.mem_538_sv2v_reg ;
  assign \nz.mem [537] = \nz.mem_537_sv2v_reg ;
  assign \nz.mem [536] = \nz.mem_536_sv2v_reg ;
  assign \nz.mem [535] = \nz.mem_535_sv2v_reg ;
  assign \nz.mem [534] = \nz.mem_534_sv2v_reg ;
  assign \nz.mem [533] = \nz.mem_533_sv2v_reg ;
  assign \nz.mem [532] = \nz.mem_532_sv2v_reg ;
  assign \nz.mem [531] = \nz.mem_531_sv2v_reg ;
  assign \nz.mem [530] = \nz.mem_530_sv2v_reg ;
  assign \nz.mem [529] = \nz.mem_529_sv2v_reg ;
  assign \nz.mem [528] = \nz.mem_528_sv2v_reg ;
  assign \nz.mem [527] = \nz.mem_527_sv2v_reg ;
  assign \nz.mem [526] = \nz.mem_526_sv2v_reg ;
  assign \nz.mem [525] = \nz.mem_525_sv2v_reg ;
  assign \nz.mem [524] = \nz.mem_524_sv2v_reg ;
  assign \nz.mem [523] = \nz.mem_523_sv2v_reg ;
  assign \nz.mem [522] = \nz.mem_522_sv2v_reg ;
  assign \nz.mem [521] = \nz.mem_521_sv2v_reg ;
  assign \nz.mem [520] = \nz.mem_520_sv2v_reg ;
  assign \nz.mem [519] = \nz.mem_519_sv2v_reg ;
  assign \nz.mem [518] = \nz.mem_518_sv2v_reg ;
  assign \nz.mem [517] = \nz.mem_517_sv2v_reg ;
  assign \nz.mem [516] = \nz.mem_516_sv2v_reg ;
  assign \nz.mem [515] = \nz.mem_515_sv2v_reg ;
  assign \nz.mem [514] = \nz.mem_514_sv2v_reg ;
  assign \nz.mem [513] = \nz.mem_513_sv2v_reg ;
  assign \nz.mem [512] = \nz.mem_512_sv2v_reg ;
  assign \nz.mem [511] = \nz.mem_511_sv2v_reg ;
  assign \nz.mem [510] = \nz.mem_510_sv2v_reg ;
  assign \nz.mem [509] = \nz.mem_509_sv2v_reg ;
  assign \nz.mem [508] = \nz.mem_508_sv2v_reg ;
  assign \nz.mem [507] = \nz.mem_507_sv2v_reg ;
  assign \nz.mem [506] = \nz.mem_506_sv2v_reg ;
  assign \nz.mem [505] = \nz.mem_505_sv2v_reg ;
  assign \nz.mem [504] = \nz.mem_504_sv2v_reg ;
  assign \nz.mem [503] = \nz.mem_503_sv2v_reg ;
  assign \nz.mem [502] = \nz.mem_502_sv2v_reg ;
  assign \nz.mem [501] = \nz.mem_501_sv2v_reg ;
  assign \nz.mem [500] = \nz.mem_500_sv2v_reg ;
  assign \nz.mem [499] = \nz.mem_499_sv2v_reg ;
  assign \nz.mem [498] = \nz.mem_498_sv2v_reg ;
  assign \nz.mem [497] = \nz.mem_497_sv2v_reg ;
  assign \nz.mem [496] = \nz.mem_496_sv2v_reg ;
  assign \nz.mem [495] = \nz.mem_495_sv2v_reg ;
  assign \nz.mem [494] = \nz.mem_494_sv2v_reg ;
  assign \nz.mem [493] = \nz.mem_493_sv2v_reg ;
  assign \nz.mem [492] = \nz.mem_492_sv2v_reg ;
  assign \nz.mem [491] = \nz.mem_491_sv2v_reg ;
  assign \nz.mem [490] = \nz.mem_490_sv2v_reg ;
  assign \nz.mem [489] = \nz.mem_489_sv2v_reg ;
  assign \nz.mem [488] = \nz.mem_488_sv2v_reg ;
  assign \nz.mem [487] = \nz.mem_487_sv2v_reg ;
  assign \nz.mem [486] = \nz.mem_486_sv2v_reg ;
  assign \nz.mem [485] = \nz.mem_485_sv2v_reg ;
  assign \nz.mem [484] = \nz.mem_484_sv2v_reg ;
  assign \nz.mem [483] = \nz.mem_483_sv2v_reg ;
  assign \nz.mem [482] = \nz.mem_482_sv2v_reg ;
  assign \nz.mem [481] = \nz.mem_481_sv2v_reg ;
  assign \nz.mem [480] = \nz.mem_480_sv2v_reg ;
  assign \nz.mem [479] = \nz.mem_479_sv2v_reg ;
  assign \nz.mem [478] = \nz.mem_478_sv2v_reg ;
  assign \nz.mem [477] = \nz.mem_477_sv2v_reg ;
  assign \nz.mem [476] = \nz.mem_476_sv2v_reg ;
  assign \nz.mem [475] = \nz.mem_475_sv2v_reg ;
  assign \nz.mem [474] = \nz.mem_474_sv2v_reg ;
  assign \nz.mem [473] = \nz.mem_473_sv2v_reg ;
  assign \nz.mem [472] = \nz.mem_472_sv2v_reg ;
  assign \nz.mem [471] = \nz.mem_471_sv2v_reg ;
  assign \nz.mem [470] = \nz.mem_470_sv2v_reg ;
  assign \nz.mem [469] = \nz.mem_469_sv2v_reg ;
  assign \nz.mem [468] = \nz.mem_468_sv2v_reg ;
  assign \nz.mem [467] = \nz.mem_467_sv2v_reg ;
  assign \nz.mem [466] = \nz.mem_466_sv2v_reg ;
  assign \nz.mem [465] = \nz.mem_465_sv2v_reg ;
  assign \nz.mem [464] = \nz.mem_464_sv2v_reg ;
  assign \nz.mem [463] = \nz.mem_463_sv2v_reg ;
  assign \nz.mem [462] = \nz.mem_462_sv2v_reg ;
  assign \nz.mem [461] = \nz.mem_461_sv2v_reg ;
  assign \nz.mem [460] = \nz.mem_460_sv2v_reg ;
  assign \nz.mem [459] = \nz.mem_459_sv2v_reg ;
  assign \nz.mem [458] = \nz.mem_458_sv2v_reg ;
  assign \nz.mem [457] = \nz.mem_457_sv2v_reg ;
  assign \nz.mem [456] = \nz.mem_456_sv2v_reg ;
  assign \nz.mem [455] = \nz.mem_455_sv2v_reg ;
  assign \nz.mem [454] = \nz.mem_454_sv2v_reg ;
  assign \nz.mem [453] = \nz.mem_453_sv2v_reg ;
  assign \nz.mem [452] = \nz.mem_452_sv2v_reg ;
  assign \nz.mem [451] = \nz.mem_451_sv2v_reg ;
  assign \nz.mem [450] = \nz.mem_450_sv2v_reg ;
  assign \nz.mem [449] = \nz.mem_449_sv2v_reg ;
  assign \nz.mem [448] = \nz.mem_448_sv2v_reg ;
  assign \nz.mem [447] = \nz.mem_447_sv2v_reg ;
  assign \nz.mem [446] = \nz.mem_446_sv2v_reg ;
  assign \nz.mem [445] = \nz.mem_445_sv2v_reg ;
  assign \nz.mem [444] = \nz.mem_444_sv2v_reg ;
  assign \nz.mem [443] = \nz.mem_443_sv2v_reg ;
  assign \nz.mem [442] = \nz.mem_442_sv2v_reg ;
  assign \nz.mem [441] = \nz.mem_441_sv2v_reg ;
  assign \nz.mem [440] = \nz.mem_440_sv2v_reg ;
  assign \nz.mem [439] = \nz.mem_439_sv2v_reg ;
  assign \nz.mem [438] = \nz.mem_438_sv2v_reg ;
  assign \nz.mem [437] = \nz.mem_437_sv2v_reg ;
  assign \nz.mem [436] = \nz.mem_436_sv2v_reg ;
  assign \nz.mem [435] = \nz.mem_435_sv2v_reg ;
  assign \nz.mem [434] = \nz.mem_434_sv2v_reg ;
  assign \nz.mem [433] = \nz.mem_433_sv2v_reg ;
  assign \nz.mem [432] = \nz.mem_432_sv2v_reg ;
  assign \nz.mem [431] = \nz.mem_431_sv2v_reg ;
  assign \nz.mem [430] = \nz.mem_430_sv2v_reg ;
  assign \nz.mem [429] = \nz.mem_429_sv2v_reg ;
  assign \nz.mem [428] = \nz.mem_428_sv2v_reg ;
  assign \nz.mem [427] = \nz.mem_427_sv2v_reg ;
  assign \nz.mem [426] = \nz.mem_426_sv2v_reg ;
  assign \nz.mem [425] = \nz.mem_425_sv2v_reg ;
  assign \nz.mem [424] = \nz.mem_424_sv2v_reg ;
  assign \nz.mem [423] = \nz.mem_423_sv2v_reg ;
  assign \nz.mem [422] = \nz.mem_422_sv2v_reg ;
  assign \nz.mem [421] = \nz.mem_421_sv2v_reg ;
  assign \nz.mem [420] = \nz.mem_420_sv2v_reg ;
  assign \nz.mem [419] = \nz.mem_419_sv2v_reg ;
  assign \nz.mem [418] = \nz.mem_418_sv2v_reg ;
  assign \nz.mem [417] = \nz.mem_417_sv2v_reg ;
  assign \nz.mem [416] = \nz.mem_416_sv2v_reg ;
  assign \nz.mem [415] = \nz.mem_415_sv2v_reg ;
  assign \nz.mem [414] = \nz.mem_414_sv2v_reg ;
  assign \nz.mem [413] = \nz.mem_413_sv2v_reg ;
  assign \nz.mem [412] = \nz.mem_412_sv2v_reg ;
  assign \nz.mem [411] = \nz.mem_411_sv2v_reg ;
  assign \nz.mem [410] = \nz.mem_410_sv2v_reg ;
  assign \nz.mem [409] = \nz.mem_409_sv2v_reg ;
  assign \nz.mem [408] = \nz.mem_408_sv2v_reg ;
  assign \nz.mem [407] = \nz.mem_407_sv2v_reg ;
  assign \nz.mem [406] = \nz.mem_406_sv2v_reg ;
  assign \nz.mem [405] = \nz.mem_405_sv2v_reg ;
  assign \nz.mem [404] = \nz.mem_404_sv2v_reg ;
  assign \nz.mem [403] = \nz.mem_403_sv2v_reg ;
  assign \nz.mem [402] = \nz.mem_402_sv2v_reg ;
  assign \nz.mem [401] = \nz.mem_401_sv2v_reg ;
  assign \nz.mem [400] = \nz.mem_400_sv2v_reg ;
  assign \nz.mem [399] = \nz.mem_399_sv2v_reg ;
  assign \nz.mem [398] = \nz.mem_398_sv2v_reg ;
  assign \nz.mem [397] = \nz.mem_397_sv2v_reg ;
  assign \nz.mem [396] = \nz.mem_396_sv2v_reg ;
  assign \nz.mem [395] = \nz.mem_395_sv2v_reg ;
  assign \nz.mem [394] = \nz.mem_394_sv2v_reg ;
  assign \nz.mem [393] = \nz.mem_393_sv2v_reg ;
  assign \nz.mem [392] = \nz.mem_392_sv2v_reg ;
  assign \nz.mem [391] = \nz.mem_391_sv2v_reg ;
  assign \nz.mem [390] = \nz.mem_390_sv2v_reg ;
  assign \nz.mem [389] = \nz.mem_389_sv2v_reg ;
  assign \nz.mem [388] = \nz.mem_388_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[173] = (N17)? \nz.mem [173] : 
                         (N19)? \nz.mem [347] : 
                         (N21)? \nz.mem [521] : 
                         (N23)? \nz.mem [695] : 
                         (N18)? \nz.mem [869] : 
                         (N20)? \nz.mem [1043] : 
                         (N22)? \nz.mem [1217] : 
                         (N24)? \nz.mem [1391] : 1'b0;
  assign r_data_o[172] = (N17)? \nz.mem [172] : 
                         (N19)? \nz.mem [346] : 
                         (N21)? \nz.mem [520] : 
                         (N23)? \nz.mem [694] : 
                         (N18)? \nz.mem [868] : 
                         (N20)? \nz.mem [1042] : 
                         (N22)? \nz.mem [1216] : 
                         (N24)? \nz.mem [1390] : 1'b0;
  assign r_data_o[171] = (N17)? \nz.mem [171] : 
                         (N19)? \nz.mem [345] : 
                         (N21)? \nz.mem [519] : 
                         (N23)? \nz.mem [693] : 
                         (N18)? \nz.mem [867] : 
                         (N20)? \nz.mem [1041] : 
                         (N22)? \nz.mem [1215] : 
                         (N24)? \nz.mem [1389] : 1'b0;
  assign r_data_o[170] = (N17)? \nz.mem [170] : 
                         (N19)? \nz.mem [344] : 
                         (N21)? \nz.mem [518] : 
                         (N23)? \nz.mem [692] : 
                         (N18)? \nz.mem [866] : 
                         (N20)? \nz.mem [1040] : 
                         (N22)? \nz.mem [1214] : 
                         (N24)? \nz.mem [1388] : 1'b0;
  assign r_data_o[169] = (N17)? \nz.mem [169] : 
                         (N19)? \nz.mem [343] : 
                         (N21)? \nz.mem [517] : 
                         (N23)? \nz.mem [691] : 
                         (N18)? \nz.mem [865] : 
                         (N20)? \nz.mem [1039] : 
                         (N22)? \nz.mem [1213] : 
                         (N24)? \nz.mem [1387] : 1'b0;
  assign r_data_o[168] = (N17)? \nz.mem [168] : 
                         (N19)? \nz.mem [342] : 
                         (N21)? \nz.mem [516] : 
                         (N23)? \nz.mem [690] : 
                         (N18)? \nz.mem [864] : 
                         (N20)? \nz.mem [1038] : 
                         (N22)? \nz.mem [1212] : 
                         (N24)? \nz.mem [1386] : 1'b0;
  assign r_data_o[167] = (N17)? \nz.mem [167] : 
                         (N19)? \nz.mem [341] : 
                         (N21)? \nz.mem [515] : 
                         (N23)? \nz.mem [689] : 
                         (N18)? \nz.mem [863] : 
                         (N20)? \nz.mem [1037] : 
                         (N22)? \nz.mem [1211] : 
                         (N24)? \nz.mem [1385] : 1'b0;
  assign r_data_o[166] = (N17)? \nz.mem [166] : 
                         (N19)? \nz.mem [340] : 
                         (N21)? \nz.mem [514] : 
                         (N23)? \nz.mem [688] : 
                         (N18)? \nz.mem [862] : 
                         (N20)? \nz.mem [1036] : 
                         (N22)? \nz.mem [1210] : 
                         (N24)? \nz.mem [1384] : 1'b0;
  assign r_data_o[165] = (N17)? \nz.mem [165] : 
                         (N19)? \nz.mem [339] : 
                         (N21)? \nz.mem [513] : 
                         (N23)? \nz.mem [687] : 
                         (N18)? \nz.mem [861] : 
                         (N20)? \nz.mem [1035] : 
                         (N22)? \nz.mem [1209] : 
                         (N24)? \nz.mem [1383] : 1'b0;
  assign r_data_o[164] = (N17)? \nz.mem [164] : 
                         (N19)? \nz.mem [338] : 
                         (N21)? \nz.mem [512] : 
                         (N23)? \nz.mem [686] : 
                         (N18)? \nz.mem [860] : 
                         (N20)? \nz.mem [1034] : 
                         (N22)? \nz.mem [1208] : 
                         (N24)? \nz.mem [1382] : 1'b0;
  assign r_data_o[163] = (N17)? \nz.mem [163] : 
                         (N19)? \nz.mem [337] : 
                         (N21)? \nz.mem [511] : 
                         (N23)? \nz.mem [685] : 
                         (N18)? \nz.mem [859] : 
                         (N20)? \nz.mem [1033] : 
                         (N22)? \nz.mem [1207] : 
                         (N24)? \nz.mem [1381] : 1'b0;
  assign r_data_o[162] = (N17)? \nz.mem [162] : 
                         (N19)? \nz.mem [336] : 
                         (N21)? \nz.mem [510] : 
                         (N23)? \nz.mem [684] : 
                         (N18)? \nz.mem [858] : 
                         (N20)? \nz.mem [1032] : 
                         (N22)? \nz.mem [1206] : 
                         (N24)? \nz.mem [1380] : 1'b0;
  assign r_data_o[161] = (N17)? \nz.mem [161] : 
                         (N19)? \nz.mem [335] : 
                         (N21)? \nz.mem [509] : 
                         (N23)? \nz.mem [683] : 
                         (N18)? \nz.mem [857] : 
                         (N20)? \nz.mem [1031] : 
                         (N22)? \nz.mem [1205] : 
                         (N24)? \nz.mem [1379] : 1'b0;
  assign r_data_o[160] = (N17)? \nz.mem [160] : 
                         (N19)? \nz.mem [334] : 
                         (N21)? \nz.mem [508] : 
                         (N23)? \nz.mem [682] : 
                         (N18)? \nz.mem [856] : 
                         (N20)? \nz.mem [1030] : 
                         (N22)? \nz.mem [1204] : 
                         (N24)? \nz.mem [1378] : 1'b0;
  assign r_data_o[159] = (N17)? \nz.mem [159] : 
                         (N19)? \nz.mem [333] : 
                         (N21)? \nz.mem [507] : 
                         (N23)? \nz.mem [681] : 
                         (N18)? \nz.mem [855] : 
                         (N20)? \nz.mem [1029] : 
                         (N22)? \nz.mem [1203] : 
                         (N24)? \nz.mem [1377] : 1'b0;
  assign r_data_o[158] = (N17)? \nz.mem [158] : 
                         (N19)? \nz.mem [332] : 
                         (N21)? \nz.mem [506] : 
                         (N23)? \nz.mem [680] : 
                         (N18)? \nz.mem [854] : 
                         (N20)? \nz.mem [1028] : 
                         (N22)? \nz.mem [1202] : 
                         (N24)? \nz.mem [1376] : 1'b0;
  assign r_data_o[157] = (N17)? \nz.mem [157] : 
                         (N19)? \nz.mem [331] : 
                         (N21)? \nz.mem [505] : 
                         (N23)? \nz.mem [679] : 
                         (N18)? \nz.mem [853] : 
                         (N20)? \nz.mem [1027] : 
                         (N22)? \nz.mem [1201] : 
                         (N24)? \nz.mem [1375] : 1'b0;
  assign r_data_o[156] = (N17)? \nz.mem [156] : 
                         (N19)? \nz.mem [330] : 
                         (N21)? \nz.mem [504] : 
                         (N23)? \nz.mem [678] : 
                         (N18)? \nz.mem [852] : 
                         (N20)? \nz.mem [1026] : 
                         (N22)? \nz.mem [1200] : 
                         (N24)? \nz.mem [1374] : 1'b0;
  assign r_data_o[155] = (N17)? \nz.mem [155] : 
                         (N19)? \nz.mem [329] : 
                         (N21)? \nz.mem [503] : 
                         (N23)? \nz.mem [677] : 
                         (N18)? \nz.mem [851] : 
                         (N20)? \nz.mem [1025] : 
                         (N22)? \nz.mem [1199] : 
                         (N24)? \nz.mem [1373] : 1'b0;
  assign r_data_o[154] = (N17)? \nz.mem [154] : 
                         (N19)? \nz.mem [328] : 
                         (N21)? \nz.mem [502] : 
                         (N23)? \nz.mem [676] : 
                         (N18)? \nz.mem [850] : 
                         (N20)? \nz.mem [1024] : 
                         (N22)? \nz.mem [1198] : 
                         (N24)? \nz.mem [1372] : 1'b0;
  assign r_data_o[153] = (N17)? \nz.mem [153] : 
                         (N19)? \nz.mem [327] : 
                         (N21)? \nz.mem [501] : 
                         (N23)? \nz.mem [675] : 
                         (N18)? \nz.mem [849] : 
                         (N20)? \nz.mem [1023] : 
                         (N22)? \nz.mem [1197] : 
                         (N24)? \nz.mem [1371] : 1'b0;
  assign r_data_o[152] = (N17)? \nz.mem [152] : 
                         (N19)? \nz.mem [326] : 
                         (N21)? \nz.mem [500] : 
                         (N23)? \nz.mem [674] : 
                         (N18)? \nz.mem [848] : 
                         (N20)? \nz.mem [1022] : 
                         (N22)? \nz.mem [1196] : 
                         (N24)? \nz.mem [1370] : 1'b0;
  assign r_data_o[151] = (N17)? \nz.mem [151] : 
                         (N19)? \nz.mem [325] : 
                         (N21)? \nz.mem [499] : 
                         (N23)? \nz.mem [673] : 
                         (N18)? \nz.mem [847] : 
                         (N20)? \nz.mem [1021] : 
                         (N22)? \nz.mem [1195] : 
                         (N24)? \nz.mem [1369] : 1'b0;
  assign r_data_o[150] = (N17)? \nz.mem [150] : 
                         (N19)? \nz.mem [324] : 
                         (N21)? \nz.mem [498] : 
                         (N23)? \nz.mem [672] : 
                         (N18)? \nz.mem [846] : 
                         (N20)? \nz.mem [1020] : 
                         (N22)? \nz.mem [1194] : 
                         (N24)? \nz.mem [1368] : 1'b0;
  assign r_data_o[149] = (N17)? \nz.mem [149] : 
                         (N19)? \nz.mem [323] : 
                         (N21)? \nz.mem [497] : 
                         (N23)? \nz.mem [671] : 
                         (N18)? \nz.mem [845] : 
                         (N20)? \nz.mem [1019] : 
                         (N22)? \nz.mem [1193] : 
                         (N24)? \nz.mem [1367] : 1'b0;
  assign r_data_o[148] = (N17)? \nz.mem [148] : 
                         (N19)? \nz.mem [322] : 
                         (N21)? \nz.mem [496] : 
                         (N23)? \nz.mem [670] : 
                         (N18)? \nz.mem [844] : 
                         (N20)? \nz.mem [1018] : 
                         (N22)? \nz.mem [1192] : 
                         (N24)? \nz.mem [1366] : 1'b0;
  assign r_data_o[147] = (N17)? \nz.mem [147] : 
                         (N19)? \nz.mem [321] : 
                         (N21)? \nz.mem [495] : 
                         (N23)? \nz.mem [669] : 
                         (N18)? \nz.mem [843] : 
                         (N20)? \nz.mem [1017] : 
                         (N22)? \nz.mem [1191] : 
                         (N24)? \nz.mem [1365] : 1'b0;
  assign r_data_o[146] = (N17)? \nz.mem [146] : 
                         (N19)? \nz.mem [320] : 
                         (N21)? \nz.mem [494] : 
                         (N23)? \nz.mem [668] : 
                         (N18)? \nz.mem [842] : 
                         (N20)? \nz.mem [1016] : 
                         (N22)? \nz.mem [1190] : 
                         (N24)? \nz.mem [1364] : 1'b0;
  assign r_data_o[145] = (N17)? \nz.mem [145] : 
                         (N19)? \nz.mem [319] : 
                         (N21)? \nz.mem [493] : 
                         (N23)? \nz.mem [667] : 
                         (N18)? \nz.mem [841] : 
                         (N20)? \nz.mem [1015] : 
                         (N22)? \nz.mem [1189] : 
                         (N24)? \nz.mem [1363] : 1'b0;
  assign r_data_o[144] = (N17)? \nz.mem [144] : 
                         (N19)? \nz.mem [318] : 
                         (N21)? \nz.mem [492] : 
                         (N23)? \nz.mem [666] : 
                         (N18)? \nz.mem [840] : 
                         (N20)? \nz.mem [1014] : 
                         (N22)? \nz.mem [1188] : 
                         (N24)? \nz.mem [1362] : 1'b0;
  assign r_data_o[143] = (N17)? \nz.mem [143] : 
                         (N19)? \nz.mem [317] : 
                         (N21)? \nz.mem [491] : 
                         (N23)? \nz.mem [665] : 
                         (N18)? \nz.mem [839] : 
                         (N20)? \nz.mem [1013] : 
                         (N22)? \nz.mem [1187] : 
                         (N24)? \nz.mem [1361] : 1'b0;
  assign r_data_o[142] = (N17)? \nz.mem [142] : 
                         (N19)? \nz.mem [316] : 
                         (N21)? \nz.mem [490] : 
                         (N23)? \nz.mem [664] : 
                         (N18)? \nz.mem [838] : 
                         (N20)? \nz.mem [1012] : 
                         (N22)? \nz.mem [1186] : 
                         (N24)? \nz.mem [1360] : 1'b0;
  assign r_data_o[141] = (N17)? \nz.mem [141] : 
                         (N19)? \nz.mem [315] : 
                         (N21)? \nz.mem [489] : 
                         (N23)? \nz.mem [663] : 
                         (N18)? \nz.mem [837] : 
                         (N20)? \nz.mem [1011] : 
                         (N22)? \nz.mem [1185] : 
                         (N24)? \nz.mem [1359] : 1'b0;
  assign r_data_o[140] = (N17)? \nz.mem [140] : 
                         (N19)? \nz.mem [314] : 
                         (N21)? \nz.mem [488] : 
                         (N23)? \nz.mem [662] : 
                         (N18)? \nz.mem [836] : 
                         (N20)? \nz.mem [1010] : 
                         (N22)? \nz.mem [1184] : 
                         (N24)? \nz.mem [1358] : 1'b0;
  assign r_data_o[139] = (N17)? \nz.mem [139] : 
                         (N19)? \nz.mem [313] : 
                         (N21)? \nz.mem [487] : 
                         (N23)? \nz.mem [661] : 
                         (N18)? \nz.mem [835] : 
                         (N20)? \nz.mem [1009] : 
                         (N22)? \nz.mem [1183] : 
                         (N24)? \nz.mem [1357] : 1'b0;
  assign r_data_o[138] = (N17)? \nz.mem [138] : 
                         (N19)? \nz.mem [312] : 
                         (N21)? \nz.mem [486] : 
                         (N23)? \nz.mem [660] : 
                         (N18)? \nz.mem [834] : 
                         (N20)? \nz.mem [1008] : 
                         (N22)? \nz.mem [1182] : 
                         (N24)? \nz.mem [1356] : 1'b0;
  assign r_data_o[137] = (N17)? \nz.mem [137] : 
                         (N19)? \nz.mem [311] : 
                         (N21)? \nz.mem [485] : 
                         (N23)? \nz.mem [659] : 
                         (N18)? \nz.mem [833] : 
                         (N20)? \nz.mem [1007] : 
                         (N22)? \nz.mem [1181] : 
                         (N24)? \nz.mem [1355] : 1'b0;
  assign r_data_o[136] = (N17)? \nz.mem [136] : 
                         (N19)? \nz.mem [310] : 
                         (N21)? \nz.mem [484] : 
                         (N23)? \nz.mem [658] : 
                         (N18)? \nz.mem [832] : 
                         (N20)? \nz.mem [1006] : 
                         (N22)? \nz.mem [1180] : 
                         (N24)? \nz.mem [1354] : 1'b0;
  assign r_data_o[135] = (N17)? \nz.mem [135] : 
                         (N19)? \nz.mem [309] : 
                         (N21)? \nz.mem [483] : 
                         (N23)? \nz.mem [657] : 
                         (N18)? \nz.mem [831] : 
                         (N20)? \nz.mem [1005] : 
                         (N22)? \nz.mem [1179] : 
                         (N24)? \nz.mem [1353] : 1'b0;
  assign r_data_o[134] = (N17)? \nz.mem [134] : 
                         (N19)? \nz.mem [308] : 
                         (N21)? \nz.mem [482] : 
                         (N23)? \nz.mem [656] : 
                         (N18)? \nz.mem [830] : 
                         (N20)? \nz.mem [1004] : 
                         (N22)? \nz.mem [1178] : 
                         (N24)? \nz.mem [1352] : 1'b0;
  assign r_data_o[133] = (N17)? \nz.mem [133] : 
                         (N19)? \nz.mem [307] : 
                         (N21)? \nz.mem [481] : 
                         (N23)? \nz.mem [655] : 
                         (N18)? \nz.mem [829] : 
                         (N20)? \nz.mem [1003] : 
                         (N22)? \nz.mem [1177] : 
                         (N24)? \nz.mem [1351] : 1'b0;
  assign r_data_o[132] = (N17)? \nz.mem [132] : 
                         (N19)? \nz.mem [306] : 
                         (N21)? \nz.mem [480] : 
                         (N23)? \nz.mem [654] : 
                         (N18)? \nz.mem [828] : 
                         (N20)? \nz.mem [1002] : 
                         (N22)? \nz.mem [1176] : 
                         (N24)? \nz.mem [1350] : 1'b0;
  assign r_data_o[131] = (N17)? \nz.mem [131] : 
                         (N19)? \nz.mem [305] : 
                         (N21)? \nz.mem [479] : 
                         (N23)? \nz.mem [653] : 
                         (N18)? \nz.mem [827] : 
                         (N20)? \nz.mem [1001] : 
                         (N22)? \nz.mem [1175] : 
                         (N24)? \nz.mem [1349] : 1'b0;
  assign r_data_o[130] = (N17)? \nz.mem [130] : 
                         (N19)? \nz.mem [304] : 
                         (N21)? \nz.mem [478] : 
                         (N23)? \nz.mem [652] : 
                         (N18)? \nz.mem [826] : 
                         (N20)? \nz.mem [1000] : 
                         (N22)? \nz.mem [1174] : 
                         (N24)? \nz.mem [1348] : 1'b0;
  assign r_data_o[129] = (N17)? \nz.mem [129] : 
                         (N19)? \nz.mem [303] : 
                         (N21)? \nz.mem [477] : 
                         (N23)? \nz.mem [651] : 
                         (N18)? \nz.mem [825] : 
                         (N20)? \nz.mem [999] : 
                         (N22)? \nz.mem [1173] : 
                         (N24)? \nz.mem [1347] : 1'b0;
  assign r_data_o[128] = (N17)? \nz.mem [128] : 
                         (N19)? \nz.mem [302] : 
                         (N21)? \nz.mem [476] : 
                         (N23)? \nz.mem [650] : 
                         (N18)? \nz.mem [824] : 
                         (N20)? \nz.mem [998] : 
                         (N22)? \nz.mem [1172] : 
                         (N24)? \nz.mem [1346] : 1'b0;
  assign r_data_o[127] = (N17)? \nz.mem [127] : 
                         (N19)? \nz.mem [301] : 
                         (N21)? \nz.mem [475] : 
                         (N23)? \nz.mem [649] : 
                         (N18)? \nz.mem [823] : 
                         (N20)? \nz.mem [997] : 
                         (N22)? \nz.mem [1171] : 
                         (N24)? \nz.mem [1345] : 1'b0;
  assign r_data_o[126] = (N17)? \nz.mem [126] : 
                         (N19)? \nz.mem [300] : 
                         (N21)? \nz.mem [474] : 
                         (N23)? \nz.mem [648] : 
                         (N18)? \nz.mem [822] : 
                         (N20)? \nz.mem [996] : 
                         (N22)? \nz.mem [1170] : 
                         (N24)? \nz.mem [1344] : 1'b0;
  assign r_data_o[125] = (N17)? \nz.mem [125] : 
                         (N19)? \nz.mem [299] : 
                         (N21)? \nz.mem [473] : 
                         (N23)? \nz.mem [647] : 
                         (N18)? \nz.mem [821] : 
                         (N20)? \nz.mem [995] : 
                         (N22)? \nz.mem [1169] : 
                         (N24)? \nz.mem [1343] : 1'b0;
  assign r_data_o[124] = (N17)? \nz.mem [124] : 
                         (N19)? \nz.mem [298] : 
                         (N21)? \nz.mem [472] : 
                         (N23)? \nz.mem [646] : 
                         (N18)? \nz.mem [820] : 
                         (N20)? \nz.mem [994] : 
                         (N22)? \nz.mem [1168] : 
                         (N24)? \nz.mem [1342] : 1'b0;
  assign r_data_o[123] = (N17)? \nz.mem [123] : 
                         (N19)? \nz.mem [297] : 
                         (N21)? \nz.mem [471] : 
                         (N23)? \nz.mem [645] : 
                         (N18)? \nz.mem [819] : 
                         (N20)? \nz.mem [993] : 
                         (N22)? \nz.mem [1167] : 
                         (N24)? \nz.mem [1341] : 1'b0;
  assign r_data_o[122] = (N17)? \nz.mem [122] : 
                         (N19)? \nz.mem [296] : 
                         (N21)? \nz.mem [470] : 
                         (N23)? \nz.mem [644] : 
                         (N18)? \nz.mem [818] : 
                         (N20)? \nz.mem [992] : 
                         (N22)? \nz.mem [1166] : 
                         (N24)? \nz.mem [1340] : 1'b0;
  assign r_data_o[121] = (N17)? \nz.mem [121] : 
                         (N19)? \nz.mem [295] : 
                         (N21)? \nz.mem [469] : 
                         (N23)? \nz.mem [643] : 
                         (N18)? \nz.mem [817] : 
                         (N20)? \nz.mem [991] : 
                         (N22)? \nz.mem [1165] : 
                         (N24)? \nz.mem [1339] : 1'b0;
  assign r_data_o[120] = (N17)? \nz.mem [120] : 
                         (N19)? \nz.mem [294] : 
                         (N21)? \nz.mem [468] : 
                         (N23)? \nz.mem [642] : 
                         (N18)? \nz.mem [816] : 
                         (N20)? \nz.mem [990] : 
                         (N22)? \nz.mem [1164] : 
                         (N24)? \nz.mem [1338] : 1'b0;
  assign r_data_o[119] = (N17)? \nz.mem [119] : 
                         (N19)? \nz.mem [293] : 
                         (N21)? \nz.mem [467] : 
                         (N23)? \nz.mem [641] : 
                         (N18)? \nz.mem [815] : 
                         (N20)? \nz.mem [989] : 
                         (N22)? \nz.mem [1163] : 
                         (N24)? \nz.mem [1337] : 1'b0;
  assign r_data_o[118] = (N17)? \nz.mem [118] : 
                         (N19)? \nz.mem [292] : 
                         (N21)? \nz.mem [466] : 
                         (N23)? \nz.mem [640] : 
                         (N18)? \nz.mem [814] : 
                         (N20)? \nz.mem [988] : 
                         (N22)? \nz.mem [1162] : 
                         (N24)? \nz.mem [1336] : 1'b0;
  assign r_data_o[117] = (N17)? \nz.mem [117] : 
                         (N19)? \nz.mem [291] : 
                         (N21)? \nz.mem [465] : 
                         (N23)? \nz.mem [639] : 
                         (N18)? \nz.mem [813] : 
                         (N20)? \nz.mem [987] : 
                         (N22)? \nz.mem [1161] : 
                         (N24)? \nz.mem [1335] : 1'b0;
  assign r_data_o[116] = (N17)? \nz.mem [116] : 
                         (N19)? \nz.mem [290] : 
                         (N21)? \nz.mem [464] : 
                         (N23)? \nz.mem [638] : 
                         (N18)? \nz.mem [812] : 
                         (N20)? \nz.mem [986] : 
                         (N22)? \nz.mem [1160] : 
                         (N24)? \nz.mem [1334] : 1'b0;
  assign r_data_o[115] = (N17)? \nz.mem [115] : 
                         (N19)? \nz.mem [289] : 
                         (N21)? \nz.mem [463] : 
                         (N23)? \nz.mem [637] : 
                         (N18)? \nz.mem [811] : 
                         (N20)? \nz.mem [985] : 
                         (N22)? \nz.mem [1159] : 
                         (N24)? \nz.mem [1333] : 1'b0;
  assign r_data_o[114] = (N17)? \nz.mem [114] : 
                         (N19)? \nz.mem [288] : 
                         (N21)? \nz.mem [462] : 
                         (N23)? \nz.mem [636] : 
                         (N18)? \nz.mem [810] : 
                         (N20)? \nz.mem [984] : 
                         (N22)? \nz.mem [1158] : 
                         (N24)? \nz.mem [1332] : 1'b0;
  assign r_data_o[113] = (N17)? \nz.mem [113] : 
                         (N19)? \nz.mem [287] : 
                         (N21)? \nz.mem [461] : 
                         (N23)? \nz.mem [635] : 
                         (N18)? \nz.mem [809] : 
                         (N20)? \nz.mem [983] : 
                         (N22)? \nz.mem [1157] : 
                         (N24)? \nz.mem [1331] : 1'b0;
  assign r_data_o[112] = (N17)? \nz.mem [112] : 
                         (N19)? \nz.mem [286] : 
                         (N21)? \nz.mem [460] : 
                         (N23)? \nz.mem [634] : 
                         (N18)? \nz.mem [808] : 
                         (N20)? \nz.mem [982] : 
                         (N22)? \nz.mem [1156] : 
                         (N24)? \nz.mem [1330] : 1'b0;
  assign r_data_o[111] = (N17)? \nz.mem [111] : 
                         (N19)? \nz.mem [285] : 
                         (N21)? \nz.mem [459] : 
                         (N23)? \nz.mem [633] : 
                         (N18)? \nz.mem [807] : 
                         (N20)? \nz.mem [981] : 
                         (N22)? \nz.mem [1155] : 
                         (N24)? \nz.mem [1329] : 1'b0;
  assign r_data_o[110] = (N17)? \nz.mem [110] : 
                         (N19)? \nz.mem [284] : 
                         (N21)? \nz.mem [458] : 
                         (N23)? \nz.mem [632] : 
                         (N18)? \nz.mem [806] : 
                         (N20)? \nz.mem [980] : 
                         (N22)? \nz.mem [1154] : 
                         (N24)? \nz.mem [1328] : 1'b0;
  assign r_data_o[109] = (N17)? \nz.mem [109] : 
                         (N19)? \nz.mem [283] : 
                         (N21)? \nz.mem [457] : 
                         (N23)? \nz.mem [631] : 
                         (N18)? \nz.mem [805] : 
                         (N20)? \nz.mem [979] : 
                         (N22)? \nz.mem [1153] : 
                         (N24)? \nz.mem [1327] : 1'b0;
  assign r_data_o[108] = (N17)? \nz.mem [108] : 
                         (N19)? \nz.mem [282] : 
                         (N21)? \nz.mem [456] : 
                         (N23)? \nz.mem [630] : 
                         (N18)? \nz.mem [804] : 
                         (N20)? \nz.mem [978] : 
                         (N22)? \nz.mem [1152] : 
                         (N24)? \nz.mem [1326] : 1'b0;
  assign r_data_o[107] = (N17)? \nz.mem [107] : 
                         (N19)? \nz.mem [281] : 
                         (N21)? \nz.mem [455] : 
                         (N23)? \nz.mem [629] : 
                         (N18)? \nz.mem [803] : 
                         (N20)? \nz.mem [977] : 
                         (N22)? \nz.mem [1151] : 
                         (N24)? \nz.mem [1325] : 1'b0;
  assign r_data_o[106] = (N17)? \nz.mem [106] : 
                         (N19)? \nz.mem [280] : 
                         (N21)? \nz.mem [454] : 
                         (N23)? \nz.mem [628] : 
                         (N18)? \nz.mem [802] : 
                         (N20)? \nz.mem [976] : 
                         (N22)? \nz.mem [1150] : 
                         (N24)? \nz.mem [1324] : 1'b0;
  assign r_data_o[105] = (N17)? \nz.mem [105] : 
                         (N19)? \nz.mem [279] : 
                         (N21)? \nz.mem [453] : 
                         (N23)? \nz.mem [627] : 
                         (N18)? \nz.mem [801] : 
                         (N20)? \nz.mem [975] : 
                         (N22)? \nz.mem [1149] : 
                         (N24)? \nz.mem [1323] : 1'b0;
  assign r_data_o[104] = (N17)? \nz.mem [104] : 
                         (N19)? \nz.mem [278] : 
                         (N21)? \nz.mem [452] : 
                         (N23)? \nz.mem [626] : 
                         (N18)? \nz.mem [800] : 
                         (N20)? \nz.mem [974] : 
                         (N22)? \nz.mem [1148] : 
                         (N24)? \nz.mem [1322] : 1'b0;
  assign r_data_o[103] = (N17)? \nz.mem [103] : 
                         (N19)? \nz.mem [277] : 
                         (N21)? \nz.mem [451] : 
                         (N23)? \nz.mem [625] : 
                         (N18)? \nz.mem [799] : 
                         (N20)? \nz.mem [973] : 
                         (N22)? \nz.mem [1147] : 
                         (N24)? \nz.mem [1321] : 1'b0;
  assign r_data_o[102] = (N17)? \nz.mem [102] : 
                         (N19)? \nz.mem [276] : 
                         (N21)? \nz.mem [450] : 
                         (N23)? \nz.mem [624] : 
                         (N18)? \nz.mem [798] : 
                         (N20)? \nz.mem [972] : 
                         (N22)? \nz.mem [1146] : 
                         (N24)? \nz.mem [1320] : 1'b0;
  assign r_data_o[101] = (N17)? \nz.mem [101] : 
                         (N19)? \nz.mem [275] : 
                         (N21)? \nz.mem [449] : 
                         (N23)? \nz.mem [623] : 
                         (N18)? \nz.mem [797] : 
                         (N20)? \nz.mem [971] : 
                         (N22)? \nz.mem [1145] : 
                         (N24)? \nz.mem [1319] : 1'b0;
  assign r_data_o[100] = (N17)? \nz.mem [100] : 
                         (N19)? \nz.mem [274] : 
                         (N21)? \nz.mem [448] : 
                         (N23)? \nz.mem [622] : 
                         (N18)? \nz.mem [796] : 
                         (N20)? \nz.mem [970] : 
                         (N22)? \nz.mem [1144] : 
                         (N24)? \nz.mem [1318] : 1'b0;
  assign r_data_o[99] = (N17)? \nz.mem [99] : 
                        (N19)? \nz.mem [273] : 
                        (N21)? \nz.mem [447] : 
                        (N23)? \nz.mem [621] : 
                        (N18)? \nz.mem [795] : 
                        (N20)? \nz.mem [969] : 
                        (N22)? \nz.mem [1143] : 
                        (N24)? \nz.mem [1317] : 1'b0;
  assign r_data_o[98] = (N17)? \nz.mem [98] : 
                        (N19)? \nz.mem [272] : 
                        (N21)? \nz.mem [446] : 
                        (N23)? \nz.mem [620] : 
                        (N18)? \nz.mem [794] : 
                        (N20)? \nz.mem [968] : 
                        (N22)? \nz.mem [1142] : 
                        (N24)? \nz.mem [1316] : 1'b0;
  assign r_data_o[97] = (N17)? \nz.mem [97] : 
                        (N19)? \nz.mem [271] : 
                        (N21)? \nz.mem [445] : 
                        (N23)? \nz.mem [619] : 
                        (N18)? \nz.mem [793] : 
                        (N20)? \nz.mem [967] : 
                        (N22)? \nz.mem [1141] : 
                        (N24)? \nz.mem [1315] : 1'b0;
  assign r_data_o[96] = (N17)? \nz.mem [96] : 
                        (N19)? \nz.mem [270] : 
                        (N21)? \nz.mem [444] : 
                        (N23)? \nz.mem [618] : 
                        (N18)? \nz.mem [792] : 
                        (N20)? \nz.mem [966] : 
                        (N22)? \nz.mem [1140] : 
                        (N24)? \nz.mem [1314] : 1'b0;
  assign r_data_o[95] = (N17)? \nz.mem [95] : 
                        (N19)? \nz.mem [269] : 
                        (N21)? \nz.mem [443] : 
                        (N23)? \nz.mem [617] : 
                        (N18)? \nz.mem [791] : 
                        (N20)? \nz.mem [965] : 
                        (N22)? \nz.mem [1139] : 
                        (N24)? \nz.mem [1313] : 1'b0;
  assign r_data_o[94] = (N17)? \nz.mem [94] : 
                        (N19)? \nz.mem [268] : 
                        (N21)? \nz.mem [442] : 
                        (N23)? \nz.mem [616] : 
                        (N18)? \nz.mem [790] : 
                        (N20)? \nz.mem [964] : 
                        (N22)? \nz.mem [1138] : 
                        (N24)? \nz.mem [1312] : 1'b0;
  assign r_data_o[93] = (N17)? \nz.mem [93] : 
                        (N19)? \nz.mem [267] : 
                        (N21)? \nz.mem [441] : 
                        (N23)? \nz.mem [615] : 
                        (N18)? \nz.mem [789] : 
                        (N20)? \nz.mem [963] : 
                        (N22)? \nz.mem [1137] : 
                        (N24)? \nz.mem [1311] : 1'b0;
  assign r_data_o[92] = (N17)? \nz.mem [92] : 
                        (N19)? \nz.mem [266] : 
                        (N21)? \nz.mem [440] : 
                        (N23)? \nz.mem [614] : 
                        (N18)? \nz.mem [788] : 
                        (N20)? \nz.mem [962] : 
                        (N22)? \nz.mem [1136] : 
                        (N24)? \nz.mem [1310] : 1'b0;
  assign r_data_o[91] = (N17)? \nz.mem [91] : 
                        (N19)? \nz.mem [265] : 
                        (N21)? \nz.mem [439] : 
                        (N23)? \nz.mem [613] : 
                        (N18)? \nz.mem [787] : 
                        (N20)? \nz.mem [961] : 
                        (N22)? \nz.mem [1135] : 
                        (N24)? \nz.mem [1309] : 1'b0;
  assign r_data_o[90] = (N17)? \nz.mem [90] : 
                        (N19)? \nz.mem [264] : 
                        (N21)? \nz.mem [438] : 
                        (N23)? \nz.mem [612] : 
                        (N18)? \nz.mem [786] : 
                        (N20)? \nz.mem [960] : 
                        (N22)? \nz.mem [1134] : 
                        (N24)? \nz.mem [1308] : 1'b0;
  assign r_data_o[89] = (N17)? \nz.mem [89] : 
                        (N19)? \nz.mem [263] : 
                        (N21)? \nz.mem [437] : 
                        (N23)? \nz.mem [611] : 
                        (N18)? \nz.mem [785] : 
                        (N20)? \nz.mem [959] : 
                        (N22)? \nz.mem [1133] : 
                        (N24)? \nz.mem [1307] : 1'b0;
  assign r_data_o[88] = (N17)? \nz.mem [88] : 
                        (N19)? \nz.mem [262] : 
                        (N21)? \nz.mem [436] : 
                        (N23)? \nz.mem [610] : 
                        (N18)? \nz.mem [784] : 
                        (N20)? \nz.mem [958] : 
                        (N22)? \nz.mem [1132] : 
                        (N24)? \nz.mem [1306] : 1'b0;
  assign r_data_o[87] = (N17)? \nz.mem [87] : 
                        (N19)? \nz.mem [261] : 
                        (N21)? \nz.mem [435] : 
                        (N23)? \nz.mem [609] : 
                        (N18)? \nz.mem [783] : 
                        (N20)? \nz.mem [957] : 
                        (N22)? \nz.mem [1131] : 
                        (N24)? \nz.mem [1305] : 1'b0;
  assign r_data_o[86] = (N17)? \nz.mem [86] : 
                        (N19)? \nz.mem [260] : 
                        (N21)? \nz.mem [434] : 
                        (N23)? \nz.mem [608] : 
                        (N18)? \nz.mem [782] : 
                        (N20)? \nz.mem [956] : 
                        (N22)? \nz.mem [1130] : 
                        (N24)? \nz.mem [1304] : 1'b0;
  assign r_data_o[85] = (N17)? \nz.mem [85] : 
                        (N19)? \nz.mem [259] : 
                        (N21)? \nz.mem [433] : 
                        (N23)? \nz.mem [607] : 
                        (N18)? \nz.mem [781] : 
                        (N20)? \nz.mem [955] : 
                        (N22)? \nz.mem [1129] : 
                        (N24)? \nz.mem [1303] : 1'b0;
  assign r_data_o[84] = (N17)? \nz.mem [84] : 
                        (N19)? \nz.mem [258] : 
                        (N21)? \nz.mem [432] : 
                        (N23)? \nz.mem [606] : 
                        (N18)? \nz.mem [780] : 
                        (N20)? \nz.mem [954] : 
                        (N22)? \nz.mem [1128] : 
                        (N24)? \nz.mem [1302] : 1'b0;
  assign r_data_o[83] = (N17)? \nz.mem [83] : 
                        (N19)? \nz.mem [257] : 
                        (N21)? \nz.mem [431] : 
                        (N23)? \nz.mem [605] : 
                        (N18)? \nz.mem [779] : 
                        (N20)? \nz.mem [953] : 
                        (N22)? \nz.mem [1127] : 
                        (N24)? \nz.mem [1301] : 1'b0;
  assign r_data_o[82] = (N17)? \nz.mem [82] : 
                        (N19)? \nz.mem [256] : 
                        (N21)? \nz.mem [430] : 
                        (N23)? \nz.mem [604] : 
                        (N18)? \nz.mem [778] : 
                        (N20)? \nz.mem [952] : 
                        (N22)? \nz.mem [1126] : 
                        (N24)? \nz.mem [1300] : 1'b0;
  assign r_data_o[81] = (N17)? \nz.mem [81] : 
                        (N19)? \nz.mem [255] : 
                        (N21)? \nz.mem [429] : 
                        (N23)? \nz.mem [603] : 
                        (N18)? \nz.mem [777] : 
                        (N20)? \nz.mem [951] : 
                        (N22)? \nz.mem [1125] : 
                        (N24)? \nz.mem [1299] : 1'b0;
  assign r_data_o[80] = (N17)? \nz.mem [80] : 
                        (N19)? \nz.mem [254] : 
                        (N21)? \nz.mem [428] : 
                        (N23)? \nz.mem [602] : 
                        (N18)? \nz.mem [776] : 
                        (N20)? \nz.mem [950] : 
                        (N22)? \nz.mem [1124] : 
                        (N24)? \nz.mem [1298] : 1'b0;
  assign r_data_o[79] = (N17)? \nz.mem [79] : 
                        (N19)? \nz.mem [253] : 
                        (N21)? \nz.mem [427] : 
                        (N23)? \nz.mem [601] : 
                        (N18)? \nz.mem [775] : 
                        (N20)? \nz.mem [949] : 
                        (N22)? \nz.mem [1123] : 
                        (N24)? \nz.mem [1297] : 1'b0;
  assign r_data_o[78] = (N17)? \nz.mem [78] : 
                        (N19)? \nz.mem [252] : 
                        (N21)? \nz.mem [426] : 
                        (N23)? \nz.mem [600] : 
                        (N18)? \nz.mem [774] : 
                        (N20)? \nz.mem [948] : 
                        (N22)? \nz.mem [1122] : 
                        (N24)? \nz.mem [1296] : 1'b0;
  assign r_data_o[77] = (N17)? \nz.mem [77] : 
                        (N19)? \nz.mem [251] : 
                        (N21)? \nz.mem [425] : 
                        (N23)? \nz.mem [599] : 
                        (N18)? \nz.mem [773] : 
                        (N20)? \nz.mem [947] : 
                        (N22)? \nz.mem [1121] : 
                        (N24)? \nz.mem [1295] : 1'b0;
  assign r_data_o[76] = (N17)? \nz.mem [76] : 
                        (N19)? \nz.mem [250] : 
                        (N21)? \nz.mem [424] : 
                        (N23)? \nz.mem [598] : 
                        (N18)? \nz.mem [772] : 
                        (N20)? \nz.mem [946] : 
                        (N22)? \nz.mem [1120] : 
                        (N24)? \nz.mem [1294] : 1'b0;
  assign r_data_o[75] = (N17)? \nz.mem [75] : 
                        (N19)? \nz.mem [249] : 
                        (N21)? \nz.mem [423] : 
                        (N23)? \nz.mem [597] : 
                        (N18)? \nz.mem [771] : 
                        (N20)? \nz.mem [945] : 
                        (N22)? \nz.mem [1119] : 
                        (N24)? \nz.mem [1293] : 1'b0;
  assign r_data_o[74] = (N17)? \nz.mem [74] : 
                        (N19)? \nz.mem [248] : 
                        (N21)? \nz.mem [422] : 
                        (N23)? \nz.mem [596] : 
                        (N18)? \nz.mem [770] : 
                        (N20)? \nz.mem [944] : 
                        (N22)? \nz.mem [1118] : 
                        (N24)? \nz.mem [1292] : 1'b0;
  assign r_data_o[73] = (N17)? \nz.mem [73] : 
                        (N19)? \nz.mem [247] : 
                        (N21)? \nz.mem [421] : 
                        (N23)? \nz.mem [595] : 
                        (N18)? \nz.mem [769] : 
                        (N20)? \nz.mem [943] : 
                        (N22)? \nz.mem [1117] : 
                        (N24)? \nz.mem [1291] : 1'b0;
  assign r_data_o[72] = (N17)? \nz.mem [72] : 
                        (N19)? \nz.mem [246] : 
                        (N21)? \nz.mem [420] : 
                        (N23)? \nz.mem [594] : 
                        (N18)? \nz.mem [768] : 
                        (N20)? \nz.mem [942] : 
                        (N22)? \nz.mem [1116] : 
                        (N24)? \nz.mem [1290] : 1'b0;
  assign r_data_o[71] = (N17)? \nz.mem [71] : 
                        (N19)? \nz.mem [245] : 
                        (N21)? \nz.mem [419] : 
                        (N23)? \nz.mem [593] : 
                        (N18)? \nz.mem [767] : 
                        (N20)? \nz.mem [941] : 
                        (N22)? \nz.mem [1115] : 
                        (N24)? \nz.mem [1289] : 1'b0;
  assign r_data_o[70] = (N17)? \nz.mem [70] : 
                        (N19)? \nz.mem [244] : 
                        (N21)? \nz.mem [418] : 
                        (N23)? \nz.mem [592] : 
                        (N18)? \nz.mem [766] : 
                        (N20)? \nz.mem [940] : 
                        (N22)? \nz.mem [1114] : 
                        (N24)? \nz.mem [1288] : 1'b0;
  assign r_data_o[69] = (N17)? \nz.mem [69] : 
                        (N19)? \nz.mem [243] : 
                        (N21)? \nz.mem [417] : 
                        (N23)? \nz.mem [591] : 
                        (N18)? \nz.mem [765] : 
                        (N20)? \nz.mem [939] : 
                        (N22)? \nz.mem [1113] : 
                        (N24)? \nz.mem [1287] : 1'b0;
  assign r_data_o[68] = (N17)? \nz.mem [68] : 
                        (N19)? \nz.mem [242] : 
                        (N21)? \nz.mem [416] : 
                        (N23)? \nz.mem [590] : 
                        (N18)? \nz.mem [764] : 
                        (N20)? \nz.mem [938] : 
                        (N22)? \nz.mem [1112] : 
                        (N24)? \nz.mem [1286] : 1'b0;
  assign r_data_o[67] = (N17)? \nz.mem [67] : 
                        (N19)? \nz.mem [241] : 
                        (N21)? \nz.mem [415] : 
                        (N23)? \nz.mem [589] : 
                        (N18)? \nz.mem [763] : 
                        (N20)? \nz.mem [937] : 
                        (N22)? \nz.mem [1111] : 
                        (N24)? \nz.mem [1285] : 1'b0;
  assign r_data_o[66] = (N17)? \nz.mem [66] : 
                        (N19)? \nz.mem [240] : 
                        (N21)? \nz.mem [414] : 
                        (N23)? \nz.mem [588] : 
                        (N18)? \nz.mem [762] : 
                        (N20)? \nz.mem [936] : 
                        (N22)? \nz.mem [1110] : 
                        (N24)? \nz.mem [1284] : 1'b0;
  assign r_data_o[65] = (N17)? \nz.mem [65] : 
                        (N19)? \nz.mem [239] : 
                        (N21)? \nz.mem [413] : 
                        (N23)? \nz.mem [587] : 
                        (N18)? \nz.mem [761] : 
                        (N20)? \nz.mem [935] : 
                        (N22)? \nz.mem [1109] : 
                        (N24)? \nz.mem [1283] : 1'b0;
  assign r_data_o[64] = (N17)? \nz.mem [64] : 
                        (N19)? \nz.mem [238] : 
                        (N21)? \nz.mem [412] : 
                        (N23)? \nz.mem [586] : 
                        (N18)? \nz.mem [760] : 
                        (N20)? \nz.mem [934] : 
                        (N22)? \nz.mem [1108] : 
                        (N24)? \nz.mem [1282] : 1'b0;
  assign r_data_o[63] = (N17)? \nz.mem [63] : 
                        (N19)? \nz.mem [237] : 
                        (N21)? \nz.mem [411] : 
                        (N23)? \nz.mem [585] : 
                        (N18)? \nz.mem [759] : 
                        (N20)? \nz.mem [933] : 
                        (N22)? \nz.mem [1107] : 
                        (N24)? \nz.mem [1281] : 1'b0;
  assign r_data_o[62] = (N17)? \nz.mem [62] : 
                        (N19)? \nz.mem [236] : 
                        (N21)? \nz.mem [410] : 
                        (N23)? \nz.mem [584] : 
                        (N18)? \nz.mem [758] : 
                        (N20)? \nz.mem [932] : 
                        (N22)? \nz.mem [1106] : 
                        (N24)? \nz.mem [1280] : 1'b0;
  assign r_data_o[61] = (N17)? \nz.mem [61] : 
                        (N19)? \nz.mem [235] : 
                        (N21)? \nz.mem [409] : 
                        (N23)? \nz.mem [583] : 
                        (N18)? \nz.mem [757] : 
                        (N20)? \nz.mem [931] : 
                        (N22)? \nz.mem [1105] : 
                        (N24)? \nz.mem [1279] : 1'b0;
  assign r_data_o[60] = (N17)? \nz.mem [60] : 
                        (N19)? \nz.mem [234] : 
                        (N21)? \nz.mem [408] : 
                        (N23)? \nz.mem [582] : 
                        (N18)? \nz.mem [756] : 
                        (N20)? \nz.mem [930] : 
                        (N22)? \nz.mem [1104] : 
                        (N24)? \nz.mem [1278] : 1'b0;
  assign r_data_o[59] = (N17)? \nz.mem [59] : 
                        (N19)? \nz.mem [233] : 
                        (N21)? \nz.mem [407] : 
                        (N23)? \nz.mem [581] : 
                        (N18)? \nz.mem [755] : 
                        (N20)? \nz.mem [929] : 
                        (N22)? \nz.mem [1103] : 
                        (N24)? \nz.mem [1277] : 1'b0;
  assign r_data_o[58] = (N17)? \nz.mem [58] : 
                        (N19)? \nz.mem [232] : 
                        (N21)? \nz.mem [406] : 
                        (N23)? \nz.mem [580] : 
                        (N18)? \nz.mem [754] : 
                        (N20)? \nz.mem [928] : 
                        (N22)? \nz.mem [1102] : 
                        (N24)? \nz.mem [1276] : 1'b0;
  assign r_data_o[57] = (N17)? \nz.mem [57] : 
                        (N19)? \nz.mem [231] : 
                        (N21)? \nz.mem [405] : 
                        (N23)? \nz.mem [579] : 
                        (N18)? \nz.mem [753] : 
                        (N20)? \nz.mem [927] : 
                        (N22)? \nz.mem [1101] : 
                        (N24)? \nz.mem [1275] : 1'b0;
  assign r_data_o[56] = (N17)? \nz.mem [56] : 
                        (N19)? \nz.mem [230] : 
                        (N21)? \nz.mem [404] : 
                        (N23)? \nz.mem [578] : 
                        (N18)? \nz.mem [752] : 
                        (N20)? \nz.mem [926] : 
                        (N22)? \nz.mem [1100] : 
                        (N24)? \nz.mem [1274] : 1'b0;
  assign r_data_o[55] = (N17)? \nz.mem [55] : 
                        (N19)? \nz.mem [229] : 
                        (N21)? \nz.mem [403] : 
                        (N23)? \nz.mem [577] : 
                        (N18)? \nz.mem [751] : 
                        (N20)? \nz.mem [925] : 
                        (N22)? \nz.mem [1099] : 
                        (N24)? \nz.mem [1273] : 1'b0;
  assign r_data_o[54] = (N17)? \nz.mem [54] : 
                        (N19)? \nz.mem [228] : 
                        (N21)? \nz.mem [402] : 
                        (N23)? \nz.mem [576] : 
                        (N18)? \nz.mem [750] : 
                        (N20)? \nz.mem [924] : 
                        (N22)? \nz.mem [1098] : 
                        (N24)? \nz.mem [1272] : 1'b0;
  assign r_data_o[53] = (N17)? \nz.mem [53] : 
                        (N19)? \nz.mem [227] : 
                        (N21)? \nz.mem [401] : 
                        (N23)? \nz.mem [575] : 
                        (N18)? \nz.mem [749] : 
                        (N20)? \nz.mem [923] : 
                        (N22)? \nz.mem [1097] : 
                        (N24)? \nz.mem [1271] : 1'b0;
  assign r_data_o[52] = (N17)? \nz.mem [52] : 
                        (N19)? \nz.mem [226] : 
                        (N21)? \nz.mem [400] : 
                        (N23)? \nz.mem [574] : 
                        (N18)? \nz.mem [748] : 
                        (N20)? \nz.mem [922] : 
                        (N22)? \nz.mem [1096] : 
                        (N24)? \nz.mem [1270] : 1'b0;
  assign r_data_o[51] = (N17)? \nz.mem [51] : 
                        (N19)? \nz.mem [225] : 
                        (N21)? \nz.mem [399] : 
                        (N23)? \nz.mem [573] : 
                        (N18)? \nz.mem [747] : 
                        (N20)? \nz.mem [921] : 
                        (N22)? \nz.mem [1095] : 
                        (N24)? \nz.mem [1269] : 1'b0;
  assign r_data_o[50] = (N17)? \nz.mem [50] : 
                        (N19)? \nz.mem [224] : 
                        (N21)? \nz.mem [398] : 
                        (N23)? \nz.mem [572] : 
                        (N18)? \nz.mem [746] : 
                        (N20)? \nz.mem [920] : 
                        (N22)? \nz.mem [1094] : 
                        (N24)? \nz.mem [1268] : 1'b0;
  assign r_data_o[49] = (N17)? \nz.mem [49] : 
                        (N19)? \nz.mem [223] : 
                        (N21)? \nz.mem [397] : 
                        (N23)? \nz.mem [571] : 
                        (N18)? \nz.mem [745] : 
                        (N20)? \nz.mem [919] : 
                        (N22)? \nz.mem [1093] : 
                        (N24)? \nz.mem [1267] : 1'b0;
  assign r_data_o[48] = (N17)? \nz.mem [48] : 
                        (N19)? \nz.mem [222] : 
                        (N21)? \nz.mem [396] : 
                        (N23)? \nz.mem [570] : 
                        (N18)? \nz.mem [744] : 
                        (N20)? \nz.mem [918] : 
                        (N22)? \nz.mem [1092] : 
                        (N24)? \nz.mem [1266] : 1'b0;
  assign r_data_o[47] = (N17)? \nz.mem [47] : 
                        (N19)? \nz.mem [221] : 
                        (N21)? \nz.mem [395] : 
                        (N23)? \nz.mem [569] : 
                        (N18)? \nz.mem [743] : 
                        (N20)? \nz.mem [917] : 
                        (N22)? \nz.mem [1091] : 
                        (N24)? \nz.mem [1265] : 1'b0;
  assign r_data_o[46] = (N17)? \nz.mem [46] : 
                        (N19)? \nz.mem [220] : 
                        (N21)? \nz.mem [394] : 
                        (N23)? \nz.mem [568] : 
                        (N18)? \nz.mem [742] : 
                        (N20)? \nz.mem [916] : 
                        (N22)? \nz.mem [1090] : 
                        (N24)? \nz.mem [1264] : 1'b0;
  assign r_data_o[45] = (N17)? \nz.mem [45] : 
                        (N19)? \nz.mem [219] : 
                        (N21)? \nz.mem [393] : 
                        (N23)? \nz.mem [567] : 
                        (N18)? \nz.mem [741] : 
                        (N20)? \nz.mem [915] : 
                        (N22)? \nz.mem [1089] : 
                        (N24)? \nz.mem [1263] : 1'b0;
  assign r_data_o[44] = (N17)? \nz.mem [44] : 
                        (N19)? \nz.mem [218] : 
                        (N21)? \nz.mem [392] : 
                        (N23)? \nz.mem [566] : 
                        (N18)? \nz.mem [740] : 
                        (N20)? \nz.mem [914] : 
                        (N22)? \nz.mem [1088] : 
                        (N24)? \nz.mem [1262] : 1'b0;
  assign r_data_o[43] = (N17)? \nz.mem [43] : 
                        (N19)? \nz.mem [217] : 
                        (N21)? \nz.mem [391] : 
                        (N23)? \nz.mem [565] : 
                        (N18)? \nz.mem [739] : 
                        (N20)? \nz.mem [913] : 
                        (N22)? \nz.mem [1087] : 
                        (N24)? \nz.mem [1261] : 1'b0;
  assign r_data_o[42] = (N17)? \nz.mem [42] : 
                        (N19)? \nz.mem [216] : 
                        (N21)? \nz.mem [390] : 
                        (N23)? \nz.mem [564] : 
                        (N18)? \nz.mem [738] : 
                        (N20)? \nz.mem [912] : 
                        (N22)? \nz.mem [1086] : 
                        (N24)? \nz.mem [1260] : 1'b0;
  assign r_data_o[41] = (N17)? \nz.mem [41] : 
                        (N19)? \nz.mem [215] : 
                        (N21)? \nz.mem [389] : 
                        (N23)? \nz.mem [563] : 
                        (N18)? \nz.mem [737] : 
                        (N20)? \nz.mem [911] : 
                        (N22)? \nz.mem [1085] : 
                        (N24)? \nz.mem [1259] : 1'b0;
  assign r_data_o[40] = (N17)? \nz.mem [40] : 
                        (N19)? \nz.mem [214] : 
                        (N21)? \nz.mem [388] : 
                        (N23)? \nz.mem [562] : 
                        (N18)? \nz.mem [736] : 
                        (N20)? \nz.mem [910] : 
                        (N22)? \nz.mem [1084] : 
                        (N24)? \nz.mem [1258] : 1'b0;
  assign r_data_o[39] = (N17)? \nz.mem [39] : 
                        (N19)? \nz.mem [213] : 
                        (N21)? \nz.mem [387] : 
                        (N23)? \nz.mem [561] : 
                        (N18)? \nz.mem [735] : 
                        (N20)? \nz.mem [909] : 
                        (N22)? \nz.mem [1083] : 
                        (N24)? \nz.mem [1257] : 1'b0;
  assign r_data_o[38] = (N17)? \nz.mem [38] : 
                        (N19)? \nz.mem [212] : 
                        (N21)? \nz.mem [386] : 
                        (N23)? \nz.mem [560] : 
                        (N18)? \nz.mem [734] : 
                        (N20)? \nz.mem [908] : 
                        (N22)? \nz.mem [1082] : 
                        (N24)? \nz.mem [1256] : 1'b0;
  assign r_data_o[37] = (N17)? \nz.mem [37] : 
                        (N19)? \nz.mem [211] : 
                        (N21)? \nz.mem [385] : 
                        (N23)? \nz.mem [559] : 
                        (N18)? \nz.mem [733] : 
                        (N20)? \nz.mem [907] : 
                        (N22)? \nz.mem [1081] : 
                        (N24)? \nz.mem [1255] : 1'b0;
  assign r_data_o[36] = (N17)? \nz.mem [36] : 
                        (N19)? \nz.mem [210] : 
                        (N21)? \nz.mem [384] : 
                        (N23)? \nz.mem [558] : 
                        (N18)? \nz.mem [732] : 
                        (N20)? \nz.mem [906] : 
                        (N22)? \nz.mem [1080] : 
                        (N24)? \nz.mem [1254] : 1'b0;
  assign r_data_o[35] = (N17)? \nz.mem [35] : 
                        (N19)? \nz.mem [209] : 
                        (N21)? \nz.mem [383] : 
                        (N23)? \nz.mem [557] : 
                        (N18)? \nz.mem [731] : 
                        (N20)? \nz.mem [905] : 
                        (N22)? \nz.mem [1079] : 
                        (N24)? \nz.mem [1253] : 1'b0;
  assign r_data_o[34] = (N17)? \nz.mem [34] : 
                        (N19)? \nz.mem [208] : 
                        (N21)? \nz.mem [382] : 
                        (N23)? \nz.mem [556] : 
                        (N18)? \nz.mem [730] : 
                        (N20)? \nz.mem [904] : 
                        (N22)? \nz.mem [1078] : 
                        (N24)? \nz.mem [1252] : 1'b0;
  assign r_data_o[33] = (N17)? \nz.mem [33] : 
                        (N19)? \nz.mem [207] : 
                        (N21)? \nz.mem [381] : 
                        (N23)? \nz.mem [555] : 
                        (N18)? \nz.mem [729] : 
                        (N20)? \nz.mem [903] : 
                        (N22)? \nz.mem [1077] : 
                        (N24)? \nz.mem [1251] : 1'b0;
  assign r_data_o[32] = (N17)? \nz.mem [32] : 
                        (N19)? \nz.mem [206] : 
                        (N21)? \nz.mem [380] : 
                        (N23)? \nz.mem [554] : 
                        (N18)? \nz.mem [728] : 
                        (N20)? \nz.mem [902] : 
                        (N22)? \nz.mem [1076] : 
                        (N24)? \nz.mem [1250] : 1'b0;
  assign r_data_o[31] = (N17)? \nz.mem [31] : 
                        (N19)? \nz.mem [205] : 
                        (N21)? \nz.mem [379] : 
                        (N23)? \nz.mem [553] : 
                        (N18)? \nz.mem [727] : 
                        (N20)? \nz.mem [901] : 
                        (N22)? \nz.mem [1075] : 
                        (N24)? \nz.mem [1249] : 1'b0;
  assign r_data_o[30] = (N17)? \nz.mem [30] : 
                        (N19)? \nz.mem [204] : 
                        (N21)? \nz.mem [378] : 
                        (N23)? \nz.mem [552] : 
                        (N18)? \nz.mem [726] : 
                        (N20)? \nz.mem [900] : 
                        (N22)? \nz.mem [1074] : 
                        (N24)? \nz.mem [1248] : 1'b0;
  assign r_data_o[29] = (N17)? \nz.mem [29] : 
                        (N19)? \nz.mem [203] : 
                        (N21)? \nz.mem [377] : 
                        (N23)? \nz.mem [551] : 
                        (N18)? \nz.mem [725] : 
                        (N20)? \nz.mem [899] : 
                        (N22)? \nz.mem [1073] : 
                        (N24)? \nz.mem [1247] : 1'b0;
  assign r_data_o[28] = (N17)? \nz.mem [28] : 
                        (N19)? \nz.mem [202] : 
                        (N21)? \nz.mem [376] : 
                        (N23)? \nz.mem [550] : 
                        (N18)? \nz.mem [724] : 
                        (N20)? \nz.mem [898] : 
                        (N22)? \nz.mem [1072] : 
                        (N24)? \nz.mem [1246] : 1'b0;
  assign r_data_o[27] = (N17)? \nz.mem [27] : 
                        (N19)? \nz.mem [201] : 
                        (N21)? \nz.mem [375] : 
                        (N23)? \nz.mem [549] : 
                        (N18)? \nz.mem [723] : 
                        (N20)? \nz.mem [897] : 
                        (N22)? \nz.mem [1071] : 
                        (N24)? \nz.mem [1245] : 1'b0;
  assign r_data_o[26] = (N17)? \nz.mem [26] : 
                        (N19)? \nz.mem [200] : 
                        (N21)? \nz.mem [374] : 
                        (N23)? \nz.mem [548] : 
                        (N18)? \nz.mem [722] : 
                        (N20)? \nz.mem [896] : 
                        (N22)? \nz.mem [1070] : 
                        (N24)? \nz.mem [1244] : 1'b0;
  assign r_data_o[25] = (N17)? \nz.mem [25] : 
                        (N19)? \nz.mem [199] : 
                        (N21)? \nz.mem [373] : 
                        (N23)? \nz.mem [547] : 
                        (N18)? \nz.mem [721] : 
                        (N20)? \nz.mem [895] : 
                        (N22)? \nz.mem [1069] : 
                        (N24)? \nz.mem [1243] : 1'b0;
  assign r_data_o[24] = (N17)? \nz.mem [24] : 
                        (N19)? \nz.mem [198] : 
                        (N21)? \nz.mem [372] : 
                        (N23)? \nz.mem [546] : 
                        (N18)? \nz.mem [720] : 
                        (N20)? \nz.mem [894] : 
                        (N22)? \nz.mem [1068] : 
                        (N24)? \nz.mem [1242] : 1'b0;
  assign r_data_o[23] = (N17)? \nz.mem [23] : 
                        (N19)? \nz.mem [197] : 
                        (N21)? \nz.mem [371] : 
                        (N23)? \nz.mem [545] : 
                        (N18)? \nz.mem [719] : 
                        (N20)? \nz.mem [893] : 
                        (N22)? \nz.mem [1067] : 
                        (N24)? \nz.mem [1241] : 1'b0;
  assign r_data_o[22] = (N17)? \nz.mem [22] : 
                        (N19)? \nz.mem [196] : 
                        (N21)? \nz.mem [370] : 
                        (N23)? \nz.mem [544] : 
                        (N18)? \nz.mem [718] : 
                        (N20)? \nz.mem [892] : 
                        (N22)? \nz.mem [1066] : 
                        (N24)? \nz.mem [1240] : 1'b0;
  assign r_data_o[21] = (N17)? \nz.mem [21] : 
                        (N19)? \nz.mem [195] : 
                        (N21)? \nz.mem [369] : 
                        (N23)? \nz.mem [543] : 
                        (N18)? \nz.mem [717] : 
                        (N20)? \nz.mem [891] : 
                        (N22)? \nz.mem [1065] : 
                        (N24)? \nz.mem [1239] : 1'b0;
  assign r_data_o[20] = (N17)? \nz.mem [20] : 
                        (N19)? \nz.mem [194] : 
                        (N21)? \nz.mem [368] : 
                        (N23)? \nz.mem [542] : 
                        (N18)? \nz.mem [716] : 
                        (N20)? \nz.mem [890] : 
                        (N22)? \nz.mem [1064] : 
                        (N24)? \nz.mem [1238] : 1'b0;
  assign r_data_o[19] = (N17)? \nz.mem [19] : 
                        (N19)? \nz.mem [193] : 
                        (N21)? \nz.mem [367] : 
                        (N23)? \nz.mem [541] : 
                        (N18)? \nz.mem [715] : 
                        (N20)? \nz.mem [889] : 
                        (N22)? \nz.mem [1063] : 
                        (N24)? \nz.mem [1237] : 1'b0;
  assign r_data_o[18] = (N17)? \nz.mem [18] : 
                        (N19)? \nz.mem [192] : 
                        (N21)? \nz.mem [366] : 
                        (N23)? \nz.mem [540] : 
                        (N18)? \nz.mem [714] : 
                        (N20)? \nz.mem [888] : 
                        (N22)? \nz.mem [1062] : 
                        (N24)? \nz.mem [1236] : 1'b0;
  assign r_data_o[17] = (N17)? \nz.mem [17] : 
                        (N19)? \nz.mem [191] : 
                        (N21)? \nz.mem [365] : 
                        (N23)? \nz.mem [539] : 
                        (N18)? \nz.mem [713] : 
                        (N20)? \nz.mem [887] : 
                        (N22)? \nz.mem [1061] : 
                        (N24)? \nz.mem [1235] : 1'b0;
  assign r_data_o[16] = (N17)? \nz.mem [16] : 
                        (N19)? \nz.mem [190] : 
                        (N21)? \nz.mem [364] : 
                        (N23)? \nz.mem [538] : 
                        (N18)? \nz.mem [712] : 
                        (N20)? \nz.mem [886] : 
                        (N22)? \nz.mem [1060] : 
                        (N24)? \nz.mem [1234] : 1'b0;
  assign r_data_o[15] = (N17)? \nz.mem [15] : 
                        (N19)? \nz.mem [189] : 
                        (N21)? \nz.mem [363] : 
                        (N23)? \nz.mem [537] : 
                        (N18)? \nz.mem [711] : 
                        (N20)? \nz.mem [885] : 
                        (N22)? \nz.mem [1059] : 
                        (N24)? \nz.mem [1233] : 1'b0;
  assign r_data_o[14] = (N17)? \nz.mem [14] : 
                        (N19)? \nz.mem [188] : 
                        (N21)? \nz.mem [362] : 
                        (N23)? \nz.mem [536] : 
                        (N18)? \nz.mem [710] : 
                        (N20)? \nz.mem [884] : 
                        (N22)? \nz.mem [1058] : 
                        (N24)? \nz.mem [1232] : 1'b0;
  assign r_data_o[13] = (N17)? \nz.mem [13] : 
                        (N19)? \nz.mem [187] : 
                        (N21)? \nz.mem [361] : 
                        (N23)? \nz.mem [535] : 
                        (N18)? \nz.mem [709] : 
                        (N20)? \nz.mem [883] : 
                        (N22)? \nz.mem [1057] : 
                        (N24)? \nz.mem [1231] : 1'b0;
  assign r_data_o[12] = (N17)? \nz.mem [12] : 
                        (N19)? \nz.mem [186] : 
                        (N21)? \nz.mem [360] : 
                        (N23)? \nz.mem [534] : 
                        (N18)? \nz.mem [708] : 
                        (N20)? \nz.mem [882] : 
                        (N22)? \nz.mem [1056] : 
                        (N24)? \nz.mem [1230] : 1'b0;
  assign r_data_o[11] = (N17)? \nz.mem [11] : 
                        (N19)? \nz.mem [185] : 
                        (N21)? \nz.mem [359] : 
                        (N23)? \nz.mem [533] : 
                        (N18)? \nz.mem [707] : 
                        (N20)? \nz.mem [881] : 
                        (N22)? \nz.mem [1055] : 
                        (N24)? \nz.mem [1229] : 1'b0;
  assign r_data_o[10] = (N17)? \nz.mem [10] : 
                        (N19)? \nz.mem [184] : 
                        (N21)? \nz.mem [358] : 
                        (N23)? \nz.mem [532] : 
                        (N18)? \nz.mem [706] : 
                        (N20)? \nz.mem [880] : 
                        (N22)? \nz.mem [1054] : 
                        (N24)? \nz.mem [1228] : 1'b0;
  assign r_data_o[9] = (N17)? \nz.mem [9] : 
                       (N19)? \nz.mem [183] : 
                       (N21)? \nz.mem [357] : 
                       (N23)? \nz.mem [531] : 
                       (N18)? \nz.mem [705] : 
                       (N20)? \nz.mem [879] : 
                       (N22)? \nz.mem [1053] : 
                       (N24)? \nz.mem [1227] : 1'b0;
  assign r_data_o[8] = (N17)? \nz.mem [8] : 
                       (N19)? \nz.mem [182] : 
                       (N21)? \nz.mem [356] : 
                       (N23)? \nz.mem [530] : 
                       (N18)? \nz.mem [704] : 
                       (N20)? \nz.mem [878] : 
                       (N22)? \nz.mem [1052] : 
                       (N24)? \nz.mem [1226] : 1'b0;
  assign r_data_o[7] = (N17)? \nz.mem [7] : 
                       (N19)? \nz.mem [181] : 
                       (N21)? \nz.mem [355] : 
                       (N23)? \nz.mem [529] : 
                       (N18)? \nz.mem [703] : 
                       (N20)? \nz.mem [877] : 
                       (N22)? \nz.mem [1051] : 
                       (N24)? \nz.mem [1225] : 1'b0;
  assign r_data_o[6] = (N17)? \nz.mem [6] : 
                       (N19)? \nz.mem [180] : 
                       (N21)? \nz.mem [354] : 
                       (N23)? \nz.mem [528] : 
                       (N18)? \nz.mem [702] : 
                       (N20)? \nz.mem [876] : 
                       (N22)? \nz.mem [1050] : 
                       (N24)? \nz.mem [1224] : 1'b0;
  assign r_data_o[5] = (N17)? \nz.mem [5] : 
                       (N19)? \nz.mem [179] : 
                       (N21)? \nz.mem [353] : 
                       (N23)? \nz.mem [527] : 
                       (N18)? \nz.mem [701] : 
                       (N20)? \nz.mem [875] : 
                       (N22)? \nz.mem [1049] : 
                       (N24)? \nz.mem [1223] : 1'b0;
  assign r_data_o[4] = (N17)? \nz.mem [4] : 
                       (N19)? \nz.mem [178] : 
                       (N21)? \nz.mem [352] : 
                       (N23)? \nz.mem [526] : 
                       (N18)? \nz.mem [700] : 
                       (N20)? \nz.mem [874] : 
                       (N22)? \nz.mem [1048] : 
                       (N24)? \nz.mem [1222] : 1'b0;
  assign r_data_o[3] = (N17)? \nz.mem [3] : 
                       (N19)? \nz.mem [177] : 
                       (N21)? \nz.mem [351] : 
                       (N23)? \nz.mem [525] : 
                       (N18)? \nz.mem [699] : 
                       (N20)? \nz.mem [873] : 
                       (N22)? \nz.mem [1047] : 
                       (N24)? \nz.mem [1221] : 1'b0;
  assign r_data_o[2] = (N17)? \nz.mem [2] : 
                       (N19)? \nz.mem [176] : 
                       (N21)? \nz.mem [350] : 
                       (N23)? \nz.mem [524] : 
                       (N18)? \nz.mem [698] : 
                       (N20)? \nz.mem [872] : 
                       (N22)? \nz.mem [1046] : 
                       (N24)? \nz.mem [1220] : 1'b0;
  assign r_data_o[1] = (N17)? \nz.mem [1] : 
                       (N19)? \nz.mem [175] : 
                       (N21)? \nz.mem [349] : 
                       (N23)? \nz.mem [523] : 
                       (N18)? \nz.mem [697] : 
                       (N20)? \nz.mem [871] : 
                       (N22)? \nz.mem [1045] : 
                       (N24)? \nz.mem [1219] : 1'b0;
  assign r_data_o[0] = (N17)? \nz.mem [0] : 
                       (N19)? \nz.mem [174] : 
                       (N21)? \nz.mem [348] : 
                       (N23)? \nz.mem [522] : 
                       (N18)? \nz.mem [696] : 
                       (N20)? \nz.mem [870] : 
                       (N22)? \nz.mem [1044] : 
                       (N24)? \nz.mem [1218] : 1'b0;
  assign N50 = w_addr_i[0] & w_addr_i[1];
  assign N33 = N50 & w_addr_i[2];
  assign N51 = N0 & w_addr_i[1];
  assign N0 = ~w_addr_i[0];
  assign N32 = N51 & w_addr_i[2];
  assign N52 = w_addr_i[0] & N1;
  assign N1 = ~w_addr_i[1];
  assign N31 = N52 & w_addr_i[2];
  assign N53 = N2 & N3;
  assign N2 = ~w_addr_i[0];
  assign N3 = ~w_addr_i[1];
  assign N30 = N53 & w_addr_i[2];
  assign N29 = N50 & N4;
  assign N4 = ~w_addr_i[2];
  assign N28 = N51 & N5;
  assign N5 = ~w_addr_i[2];
  assign N27 = N52 & N6;
  assign N6 = ~w_addr_i[2];
  assign N26 = N53 & N7;
  assign N7 = ~w_addr_i[2];
  assign { N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34 } = (N8)? { N33, N33, N32, N32, N31, N31, N30, N30, N29, N29, N28, N28, N27, N27, N26, N26 } : 
                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N25;
  assign N10 = ~r_addr_i[0];
  assign N11 = ~r_addr_i[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r_addr_i[1];
  assign N14 = r_addr_i[0] & N11;
  assign N15 = r_addr_i[0] & r_addr_i[1];
  assign N16 = ~r_addr_i[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r_addr_i[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r_addr_i[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r_addr_i[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r_addr_i[2];
  assign N25 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N48) begin
      \nz.mem_1391_sv2v_reg  <= w_data_i[173];
      \nz.mem_1390_sv2v_reg  <= w_data_i[172];
      \nz.mem_1389_sv2v_reg  <= w_data_i[171];
      \nz.mem_1388_sv2v_reg  <= w_data_i[170];
      \nz.mem_1387_sv2v_reg  <= w_data_i[169];
      \nz.mem_1386_sv2v_reg  <= w_data_i[168];
      \nz.mem_1385_sv2v_reg  <= w_data_i[167];
      \nz.mem_1384_sv2v_reg  <= w_data_i[166];
      \nz.mem_1383_sv2v_reg  <= w_data_i[165];
      \nz.mem_1382_sv2v_reg  <= w_data_i[164];
      \nz.mem_1381_sv2v_reg  <= w_data_i[163];
      \nz.mem_1380_sv2v_reg  <= w_data_i[162];
      \nz.mem_1379_sv2v_reg  <= w_data_i[161];
      \nz.mem_1378_sv2v_reg  <= w_data_i[160];
      \nz.mem_1377_sv2v_reg  <= w_data_i[159];
      \nz.mem_1376_sv2v_reg  <= w_data_i[158];
      \nz.mem_1375_sv2v_reg  <= w_data_i[157];
      \nz.mem_1374_sv2v_reg  <= w_data_i[156];
      \nz.mem_1373_sv2v_reg  <= w_data_i[155];
      \nz.mem_1372_sv2v_reg  <= w_data_i[154];
      \nz.mem_1371_sv2v_reg  <= w_data_i[153];
      \nz.mem_1370_sv2v_reg  <= w_data_i[152];
      \nz.mem_1369_sv2v_reg  <= w_data_i[151];
      \nz.mem_1368_sv2v_reg  <= w_data_i[150];
      \nz.mem_1367_sv2v_reg  <= w_data_i[149];
      \nz.mem_1366_sv2v_reg  <= w_data_i[148];
      \nz.mem_1365_sv2v_reg  <= w_data_i[147];
      \nz.mem_1364_sv2v_reg  <= w_data_i[146];
      \nz.mem_1363_sv2v_reg  <= w_data_i[145];
      \nz.mem_1362_sv2v_reg  <= w_data_i[144];
      \nz.mem_1361_sv2v_reg  <= w_data_i[143];
      \nz.mem_1360_sv2v_reg  <= w_data_i[142];
      \nz.mem_1359_sv2v_reg  <= w_data_i[141];
      \nz.mem_1358_sv2v_reg  <= w_data_i[140];
      \nz.mem_1357_sv2v_reg  <= w_data_i[139];
      \nz.mem_1356_sv2v_reg  <= w_data_i[138];
      \nz.mem_1355_sv2v_reg  <= w_data_i[137];
      \nz.mem_1354_sv2v_reg  <= w_data_i[136];
      \nz.mem_1353_sv2v_reg  <= w_data_i[135];
      \nz.mem_1352_sv2v_reg  <= w_data_i[134];
      \nz.mem_1351_sv2v_reg  <= w_data_i[133];
      \nz.mem_1350_sv2v_reg  <= w_data_i[132];
      \nz.mem_1349_sv2v_reg  <= w_data_i[131];
      \nz.mem_1348_sv2v_reg  <= w_data_i[130];
      \nz.mem_1347_sv2v_reg  <= w_data_i[129];
      \nz.mem_1346_sv2v_reg  <= w_data_i[128];
      \nz.mem_1345_sv2v_reg  <= w_data_i[127];
      \nz.mem_1344_sv2v_reg  <= w_data_i[126];
      \nz.mem_1343_sv2v_reg  <= w_data_i[125];
      \nz.mem_1342_sv2v_reg  <= w_data_i[124];
      \nz.mem_1341_sv2v_reg  <= w_data_i[123];
      \nz.mem_1340_sv2v_reg  <= w_data_i[122];
      \nz.mem_1339_sv2v_reg  <= w_data_i[121];
      \nz.mem_1338_sv2v_reg  <= w_data_i[120];
      \nz.mem_1337_sv2v_reg  <= w_data_i[119];
      \nz.mem_1336_sv2v_reg  <= w_data_i[118];
      \nz.mem_1335_sv2v_reg  <= w_data_i[117];
      \nz.mem_1334_sv2v_reg  <= w_data_i[116];
      \nz.mem_1333_sv2v_reg  <= w_data_i[115];
      \nz.mem_1332_sv2v_reg  <= w_data_i[114];
      \nz.mem_1331_sv2v_reg  <= w_data_i[113];
      \nz.mem_1330_sv2v_reg  <= w_data_i[112];
      \nz.mem_1329_sv2v_reg  <= w_data_i[111];
      \nz.mem_1328_sv2v_reg  <= w_data_i[110];
      \nz.mem_1327_sv2v_reg  <= w_data_i[109];
      \nz.mem_1326_sv2v_reg  <= w_data_i[108];
      \nz.mem_1325_sv2v_reg  <= w_data_i[107];
      \nz.mem_1324_sv2v_reg  <= w_data_i[106];
      \nz.mem_1323_sv2v_reg  <= w_data_i[105];
      \nz.mem_1322_sv2v_reg  <= w_data_i[104];
      \nz.mem_1321_sv2v_reg  <= w_data_i[103];
      \nz.mem_1320_sv2v_reg  <= w_data_i[102];
      \nz.mem_1319_sv2v_reg  <= w_data_i[101];
      \nz.mem_1318_sv2v_reg  <= w_data_i[100];
      \nz.mem_1317_sv2v_reg  <= w_data_i[99];
      \nz.mem_1316_sv2v_reg  <= w_data_i[98];
      \nz.mem_1315_sv2v_reg  <= w_data_i[97];
      \nz.mem_1314_sv2v_reg  <= w_data_i[96];
      \nz.mem_1313_sv2v_reg  <= w_data_i[95];
      \nz.mem_1312_sv2v_reg  <= w_data_i[94];
      \nz.mem_1311_sv2v_reg  <= w_data_i[93];
      \nz.mem_1310_sv2v_reg  <= w_data_i[92];
      \nz.mem_1309_sv2v_reg  <= w_data_i[91];
      \nz.mem_1308_sv2v_reg  <= w_data_i[90];
      \nz.mem_1307_sv2v_reg  <= w_data_i[89];
      \nz.mem_1306_sv2v_reg  <= w_data_i[88];
      \nz.mem_1305_sv2v_reg  <= w_data_i[87];
      \nz.mem_1304_sv2v_reg  <= w_data_i[86];
      \nz.mem_1303_sv2v_reg  <= w_data_i[85];
      \nz.mem_1302_sv2v_reg  <= w_data_i[84];
      \nz.mem_1301_sv2v_reg  <= w_data_i[83];
      \nz.mem_1300_sv2v_reg  <= w_data_i[82];
      \nz.mem_1299_sv2v_reg  <= w_data_i[81];
      \nz.mem_1298_sv2v_reg  <= w_data_i[80];
      \nz.mem_1297_sv2v_reg  <= w_data_i[79];
      \nz.mem_1296_sv2v_reg  <= w_data_i[78];
      \nz.mem_1295_sv2v_reg  <= w_data_i[77];
      \nz.mem_1294_sv2v_reg  <= w_data_i[76];
      \nz.mem_1293_sv2v_reg  <= w_data_i[75];
      \nz.mem_1218_sv2v_reg  <= w_data_i[0];
    end 
    if(N49) begin
      \nz.mem_1292_sv2v_reg  <= w_data_i[74];
      \nz.mem_1291_sv2v_reg  <= w_data_i[73];
      \nz.mem_1290_sv2v_reg  <= w_data_i[72];
      \nz.mem_1289_sv2v_reg  <= w_data_i[71];
      \nz.mem_1288_sv2v_reg  <= w_data_i[70];
      \nz.mem_1287_sv2v_reg  <= w_data_i[69];
      \nz.mem_1286_sv2v_reg  <= w_data_i[68];
      \nz.mem_1285_sv2v_reg  <= w_data_i[67];
      \nz.mem_1284_sv2v_reg  <= w_data_i[66];
      \nz.mem_1283_sv2v_reg  <= w_data_i[65];
      \nz.mem_1282_sv2v_reg  <= w_data_i[64];
      \nz.mem_1281_sv2v_reg  <= w_data_i[63];
      \nz.mem_1280_sv2v_reg  <= w_data_i[62];
      \nz.mem_1279_sv2v_reg  <= w_data_i[61];
      \nz.mem_1278_sv2v_reg  <= w_data_i[60];
      \nz.mem_1277_sv2v_reg  <= w_data_i[59];
      \nz.mem_1276_sv2v_reg  <= w_data_i[58];
      \nz.mem_1275_sv2v_reg  <= w_data_i[57];
      \nz.mem_1274_sv2v_reg  <= w_data_i[56];
      \nz.mem_1273_sv2v_reg  <= w_data_i[55];
      \nz.mem_1272_sv2v_reg  <= w_data_i[54];
      \nz.mem_1271_sv2v_reg  <= w_data_i[53];
      \nz.mem_1270_sv2v_reg  <= w_data_i[52];
      \nz.mem_1269_sv2v_reg  <= w_data_i[51];
      \nz.mem_1268_sv2v_reg  <= w_data_i[50];
      \nz.mem_1267_sv2v_reg  <= w_data_i[49];
      \nz.mem_1266_sv2v_reg  <= w_data_i[48];
      \nz.mem_1265_sv2v_reg  <= w_data_i[47];
      \nz.mem_1264_sv2v_reg  <= w_data_i[46];
      \nz.mem_1263_sv2v_reg  <= w_data_i[45];
      \nz.mem_1262_sv2v_reg  <= w_data_i[44];
      \nz.mem_1261_sv2v_reg  <= w_data_i[43];
      \nz.mem_1260_sv2v_reg  <= w_data_i[42];
      \nz.mem_1259_sv2v_reg  <= w_data_i[41];
      \nz.mem_1258_sv2v_reg  <= w_data_i[40];
      \nz.mem_1257_sv2v_reg  <= w_data_i[39];
      \nz.mem_1256_sv2v_reg  <= w_data_i[38];
      \nz.mem_1255_sv2v_reg  <= w_data_i[37];
      \nz.mem_1254_sv2v_reg  <= w_data_i[36];
      \nz.mem_1253_sv2v_reg  <= w_data_i[35];
      \nz.mem_1252_sv2v_reg  <= w_data_i[34];
      \nz.mem_1251_sv2v_reg  <= w_data_i[33];
      \nz.mem_1250_sv2v_reg  <= w_data_i[32];
      \nz.mem_1249_sv2v_reg  <= w_data_i[31];
      \nz.mem_1248_sv2v_reg  <= w_data_i[30];
      \nz.mem_1247_sv2v_reg  <= w_data_i[29];
      \nz.mem_1246_sv2v_reg  <= w_data_i[28];
      \nz.mem_1245_sv2v_reg  <= w_data_i[27];
      \nz.mem_1244_sv2v_reg  <= w_data_i[26];
      \nz.mem_1243_sv2v_reg  <= w_data_i[25];
      \nz.mem_1242_sv2v_reg  <= w_data_i[24];
      \nz.mem_1241_sv2v_reg  <= w_data_i[23];
      \nz.mem_1240_sv2v_reg  <= w_data_i[22];
      \nz.mem_1239_sv2v_reg  <= w_data_i[21];
      \nz.mem_1238_sv2v_reg  <= w_data_i[20];
      \nz.mem_1237_sv2v_reg  <= w_data_i[19];
      \nz.mem_1236_sv2v_reg  <= w_data_i[18];
      \nz.mem_1235_sv2v_reg  <= w_data_i[17];
      \nz.mem_1234_sv2v_reg  <= w_data_i[16];
      \nz.mem_1233_sv2v_reg  <= w_data_i[15];
      \nz.mem_1232_sv2v_reg  <= w_data_i[14];
      \nz.mem_1231_sv2v_reg  <= w_data_i[13];
      \nz.mem_1230_sv2v_reg  <= w_data_i[12];
      \nz.mem_1229_sv2v_reg  <= w_data_i[11];
      \nz.mem_1228_sv2v_reg  <= w_data_i[10];
      \nz.mem_1227_sv2v_reg  <= w_data_i[9];
      \nz.mem_1226_sv2v_reg  <= w_data_i[8];
      \nz.mem_1225_sv2v_reg  <= w_data_i[7];
      \nz.mem_1224_sv2v_reg  <= w_data_i[6];
      \nz.mem_1223_sv2v_reg  <= w_data_i[5];
      \nz.mem_1222_sv2v_reg  <= w_data_i[4];
      \nz.mem_1221_sv2v_reg  <= w_data_i[3];
      \nz.mem_1220_sv2v_reg  <= w_data_i[2];
      \nz.mem_1219_sv2v_reg  <= w_data_i[1];
    end 
    if(N46) begin
      \nz.mem_1217_sv2v_reg  <= w_data_i[173];
      \nz.mem_1216_sv2v_reg  <= w_data_i[172];
      \nz.mem_1215_sv2v_reg  <= w_data_i[171];
      \nz.mem_1214_sv2v_reg  <= w_data_i[170];
      \nz.mem_1213_sv2v_reg  <= w_data_i[169];
      \nz.mem_1212_sv2v_reg  <= w_data_i[168];
      \nz.mem_1211_sv2v_reg  <= w_data_i[167];
      \nz.mem_1210_sv2v_reg  <= w_data_i[166];
      \nz.mem_1209_sv2v_reg  <= w_data_i[165];
      \nz.mem_1208_sv2v_reg  <= w_data_i[164];
      \nz.mem_1207_sv2v_reg  <= w_data_i[163];
      \nz.mem_1206_sv2v_reg  <= w_data_i[162];
      \nz.mem_1205_sv2v_reg  <= w_data_i[161];
      \nz.mem_1204_sv2v_reg  <= w_data_i[160];
      \nz.mem_1203_sv2v_reg  <= w_data_i[159];
      \nz.mem_1202_sv2v_reg  <= w_data_i[158];
      \nz.mem_1201_sv2v_reg  <= w_data_i[157];
      \nz.mem_1200_sv2v_reg  <= w_data_i[156];
      \nz.mem_1199_sv2v_reg  <= w_data_i[155];
      \nz.mem_1198_sv2v_reg  <= w_data_i[154];
      \nz.mem_1197_sv2v_reg  <= w_data_i[153];
      \nz.mem_1196_sv2v_reg  <= w_data_i[152];
      \nz.mem_1195_sv2v_reg  <= w_data_i[151];
      \nz.mem_1194_sv2v_reg  <= w_data_i[150];
      \nz.mem_1193_sv2v_reg  <= w_data_i[149];
      \nz.mem_1192_sv2v_reg  <= w_data_i[148];
      \nz.mem_1191_sv2v_reg  <= w_data_i[147];
      \nz.mem_1190_sv2v_reg  <= w_data_i[146];
      \nz.mem_1189_sv2v_reg  <= w_data_i[145];
      \nz.mem_1188_sv2v_reg  <= w_data_i[144];
      \nz.mem_1187_sv2v_reg  <= w_data_i[143];
      \nz.mem_1186_sv2v_reg  <= w_data_i[142];
      \nz.mem_1185_sv2v_reg  <= w_data_i[141];
      \nz.mem_1184_sv2v_reg  <= w_data_i[140];
      \nz.mem_1183_sv2v_reg  <= w_data_i[139];
      \nz.mem_1182_sv2v_reg  <= w_data_i[138];
      \nz.mem_1181_sv2v_reg  <= w_data_i[137];
      \nz.mem_1180_sv2v_reg  <= w_data_i[136];
      \nz.mem_1179_sv2v_reg  <= w_data_i[135];
      \nz.mem_1178_sv2v_reg  <= w_data_i[134];
      \nz.mem_1177_sv2v_reg  <= w_data_i[133];
      \nz.mem_1176_sv2v_reg  <= w_data_i[132];
      \nz.mem_1175_sv2v_reg  <= w_data_i[131];
      \nz.mem_1174_sv2v_reg  <= w_data_i[130];
      \nz.mem_1173_sv2v_reg  <= w_data_i[129];
      \nz.mem_1172_sv2v_reg  <= w_data_i[128];
      \nz.mem_1171_sv2v_reg  <= w_data_i[127];
      \nz.mem_1170_sv2v_reg  <= w_data_i[126];
      \nz.mem_1169_sv2v_reg  <= w_data_i[125];
      \nz.mem_1168_sv2v_reg  <= w_data_i[124];
      \nz.mem_1167_sv2v_reg  <= w_data_i[123];
      \nz.mem_1166_sv2v_reg  <= w_data_i[122];
      \nz.mem_1165_sv2v_reg  <= w_data_i[121];
      \nz.mem_1164_sv2v_reg  <= w_data_i[120];
      \nz.mem_1163_sv2v_reg  <= w_data_i[119];
      \nz.mem_1162_sv2v_reg  <= w_data_i[118];
      \nz.mem_1161_sv2v_reg  <= w_data_i[117];
      \nz.mem_1160_sv2v_reg  <= w_data_i[116];
      \nz.mem_1159_sv2v_reg  <= w_data_i[115];
      \nz.mem_1158_sv2v_reg  <= w_data_i[114];
      \nz.mem_1157_sv2v_reg  <= w_data_i[113];
      \nz.mem_1156_sv2v_reg  <= w_data_i[112];
      \nz.mem_1155_sv2v_reg  <= w_data_i[111];
      \nz.mem_1154_sv2v_reg  <= w_data_i[110];
      \nz.mem_1153_sv2v_reg  <= w_data_i[109];
      \nz.mem_1152_sv2v_reg  <= w_data_i[108];
      \nz.mem_1151_sv2v_reg  <= w_data_i[107];
      \nz.mem_1150_sv2v_reg  <= w_data_i[106];
      \nz.mem_1149_sv2v_reg  <= w_data_i[105];
      \nz.mem_1148_sv2v_reg  <= w_data_i[104];
      \nz.mem_1147_sv2v_reg  <= w_data_i[103];
      \nz.mem_1146_sv2v_reg  <= w_data_i[102];
      \nz.mem_1145_sv2v_reg  <= w_data_i[101];
      \nz.mem_1144_sv2v_reg  <= w_data_i[100];
      \nz.mem_1143_sv2v_reg  <= w_data_i[99];
      \nz.mem_1142_sv2v_reg  <= w_data_i[98];
      \nz.mem_1141_sv2v_reg  <= w_data_i[97];
      \nz.mem_1140_sv2v_reg  <= w_data_i[96];
      \nz.mem_1139_sv2v_reg  <= w_data_i[95];
      \nz.mem_1138_sv2v_reg  <= w_data_i[94];
      \nz.mem_1137_sv2v_reg  <= w_data_i[93];
      \nz.mem_1136_sv2v_reg  <= w_data_i[92];
      \nz.mem_1135_sv2v_reg  <= w_data_i[91];
      \nz.mem_1134_sv2v_reg  <= w_data_i[90];
      \nz.mem_1133_sv2v_reg  <= w_data_i[89];
      \nz.mem_1132_sv2v_reg  <= w_data_i[88];
      \nz.mem_1131_sv2v_reg  <= w_data_i[87];
      \nz.mem_1130_sv2v_reg  <= w_data_i[86];
      \nz.mem_1129_sv2v_reg  <= w_data_i[85];
      \nz.mem_1128_sv2v_reg  <= w_data_i[84];
      \nz.mem_1127_sv2v_reg  <= w_data_i[83];
      \nz.mem_1126_sv2v_reg  <= w_data_i[82];
      \nz.mem_1125_sv2v_reg  <= w_data_i[81];
      \nz.mem_1124_sv2v_reg  <= w_data_i[80];
      \nz.mem_1123_sv2v_reg  <= w_data_i[79];
      \nz.mem_1122_sv2v_reg  <= w_data_i[78];
      \nz.mem_1121_sv2v_reg  <= w_data_i[77];
      \nz.mem_1120_sv2v_reg  <= w_data_i[76];
      \nz.mem_1119_sv2v_reg  <= w_data_i[75];
      \nz.mem_1044_sv2v_reg  <= w_data_i[0];
    end 
    if(N47) begin
      \nz.mem_1118_sv2v_reg  <= w_data_i[74];
      \nz.mem_1117_sv2v_reg  <= w_data_i[73];
      \nz.mem_1116_sv2v_reg  <= w_data_i[72];
      \nz.mem_1115_sv2v_reg  <= w_data_i[71];
      \nz.mem_1114_sv2v_reg  <= w_data_i[70];
      \nz.mem_1113_sv2v_reg  <= w_data_i[69];
      \nz.mem_1112_sv2v_reg  <= w_data_i[68];
      \nz.mem_1111_sv2v_reg  <= w_data_i[67];
      \nz.mem_1110_sv2v_reg  <= w_data_i[66];
      \nz.mem_1109_sv2v_reg  <= w_data_i[65];
      \nz.mem_1108_sv2v_reg  <= w_data_i[64];
      \nz.mem_1107_sv2v_reg  <= w_data_i[63];
      \nz.mem_1106_sv2v_reg  <= w_data_i[62];
      \nz.mem_1105_sv2v_reg  <= w_data_i[61];
      \nz.mem_1104_sv2v_reg  <= w_data_i[60];
      \nz.mem_1103_sv2v_reg  <= w_data_i[59];
      \nz.mem_1102_sv2v_reg  <= w_data_i[58];
      \nz.mem_1101_sv2v_reg  <= w_data_i[57];
      \nz.mem_1100_sv2v_reg  <= w_data_i[56];
      \nz.mem_1099_sv2v_reg  <= w_data_i[55];
      \nz.mem_1098_sv2v_reg  <= w_data_i[54];
      \nz.mem_1097_sv2v_reg  <= w_data_i[53];
      \nz.mem_1096_sv2v_reg  <= w_data_i[52];
      \nz.mem_1095_sv2v_reg  <= w_data_i[51];
      \nz.mem_1094_sv2v_reg  <= w_data_i[50];
      \nz.mem_1093_sv2v_reg  <= w_data_i[49];
      \nz.mem_1092_sv2v_reg  <= w_data_i[48];
      \nz.mem_1091_sv2v_reg  <= w_data_i[47];
      \nz.mem_1090_sv2v_reg  <= w_data_i[46];
      \nz.mem_1089_sv2v_reg  <= w_data_i[45];
      \nz.mem_1088_sv2v_reg  <= w_data_i[44];
      \nz.mem_1087_sv2v_reg  <= w_data_i[43];
      \nz.mem_1086_sv2v_reg  <= w_data_i[42];
      \nz.mem_1085_sv2v_reg  <= w_data_i[41];
      \nz.mem_1084_sv2v_reg  <= w_data_i[40];
      \nz.mem_1083_sv2v_reg  <= w_data_i[39];
      \nz.mem_1082_sv2v_reg  <= w_data_i[38];
      \nz.mem_1081_sv2v_reg  <= w_data_i[37];
      \nz.mem_1080_sv2v_reg  <= w_data_i[36];
      \nz.mem_1079_sv2v_reg  <= w_data_i[35];
      \nz.mem_1078_sv2v_reg  <= w_data_i[34];
      \nz.mem_1077_sv2v_reg  <= w_data_i[33];
      \nz.mem_1076_sv2v_reg  <= w_data_i[32];
      \nz.mem_1075_sv2v_reg  <= w_data_i[31];
      \nz.mem_1074_sv2v_reg  <= w_data_i[30];
      \nz.mem_1073_sv2v_reg  <= w_data_i[29];
      \nz.mem_1072_sv2v_reg  <= w_data_i[28];
      \nz.mem_1071_sv2v_reg  <= w_data_i[27];
      \nz.mem_1070_sv2v_reg  <= w_data_i[26];
      \nz.mem_1069_sv2v_reg  <= w_data_i[25];
      \nz.mem_1068_sv2v_reg  <= w_data_i[24];
      \nz.mem_1067_sv2v_reg  <= w_data_i[23];
      \nz.mem_1066_sv2v_reg  <= w_data_i[22];
      \nz.mem_1065_sv2v_reg  <= w_data_i[21];
      \nz.mem_1064_sv2v_reg  <= w_data_i[20];
      \nz.mem_1063_sv2v_reg  <= w_data_i[19];
      \nz.mem_1062_sv2v_reg  <= w_data_i[18];
      \nz.mem_1061_sv2v_reg  <= w_data_i[17];
      \nz.mem_1060_sv2v_reg  <= w_data_i[16];
      \nz.mem_1059_sv2v_reg  <= w_data_i[15];
      \nz.mem_1058_sv2v_reg  <= w_data_i[14];
      \nz.mem_1057_sv2v_reg  <= w_data_i[13];
      \nz.mem_1056_sv2v_reg  <= w_data_i[12];
      \nz.mem_1055_sv2v_reg  <= w_data_i[11];
      \nz.mem_1054_sv2v_reg  <= w_data_i[10];
      \nz.mem_1053_sv2v_reg  <= w_data_i[9];
      \nz.mem_1052_sv2v_reg  <= w_data_i[8];
      \nz.mem_1051_sv2v_reg  <= w_data_i[7];
      \nz.mem_1050_sv2v_reg  <= w_data_i[6];
      \nz.mem_1049_sv2v_reg  <= w_data_i[5];
      \nz.mem_1048_sv2v_reg  <= w_data_i[4];
      \nz.mem_1047_sv2v_reg  <= w_data_i[3];
      \nz.mem_1046_sv2v_reg  <= w_data_i[2];
      \nz.mem_1045_sv2v_reg  <= w_data_i[1];
    end 
    if(N44) begin
      \nz.mem_1043_sv2v_reg  <= w_data_i[173];
      \nz.mem_1042_sv2v_reg  <= w_data_i[172];
      \nz.mem_1041_sv2v_reg  <= w_data_i[171];
      \nz.mem_1040_sv2v_reg  <= w_data_i[170];
      \nz.mem_1039_sv2v_reg  <= w_data_i[169];
      \nz.mem_1038_sv2v_reg  <= w_data_i[168];
      \nz.mem_1037_sv2v_reg  <= w_data_i[167];
      \nz.mem_1036_sv2v_reg  <= w_data_i[166];
      \nz.mem_1035_sv2v_reg  <= w_data_i[165];
      \nz.mem_1034_sv2v_reg  <= w_data_i[164];
      \nz.mem_1033_sv2v_reg  <= w_data_i[163];
      \nz.mem_1032_sv2v_reg  <= w_data_i[162];
      \nz.mem_1031_sv2v_reg  <= w_data_i[161];
      \nz.mem_1030_sv2v_reg  <= w_data_i[160];
      \nz.mem_1029_sv2v_reg  <= w_data_i[159];
      \nz.mem_1028_sv2v_reg  <= w_data_i[158];
      \nz.mem_1027_sv2v_reg  <= w_data_i[157];
      \nz.mem_1026_sv2v_reg  <= w_data_i[156];
      \nz.mem_1025_sv2v_reg  <= w_data_i[155];
      \nz.mem_1024_sv2v_reg  <= w_data_i[154];
      \nz.mem_1023_sv2v_reg  <= w_data_i[153];
      \nz.mem_1022_sv2v_reg  <= w_data_i[152];
      \nz.mem_1021_sv2v_reg  <= w_data_i[151];
      \nz.mem_1020_sv2v_reg  <= w_data_i[150];
      \nz.mem_1019_sv2v_reg  <= w_data_i[149];
      \nz.mem_1018_sv2v_reg  <= w_data_i[148];
      \nz.mem_1017_sv2v_reg  <= w_data_i[147];
      \nz.mem_1016_sv2v_reg  <= w_data_i[146];
      \nz.mem_1015_sv2v_reg  <= w_data_i[145];
      \nz.mem_1014_sv2v_reg  <= w_data_i[144];
      \nz.mem_1013_sv2v_reg  <= w_data_i[143];
      \nz.mem_1012_sv2v_reg  <= w_data_i[142];
      \nz.mem_1011_sv2v_reg  <= w_data_i[141];
      \nz.mem_1010_sv2v_reg  <= w_data_i[140];
      \nz.mem_1009_sv2v_reg  <= w_data_i[139];
      \nz.mem_1008_sv2v_reg  <= w_data_i[138];
      \nz.mem_1007_sv2v_reg  <= w_data_i[137];
      \nz.mem_1006_sv2v_reg  <= w_data_i[136];
      \nz.mem_1005_sv2v_reg  <= w_data_i[135];
      \nz.mem_1004_sv2v_reg  <= w_data_i[134];
      \nz.mem_1003_sv2v_reg  <= w_data_i[133];
      \nz.mem_1002_sv2v_reg  <= w_data_i[132];
      \nz.mem_1001_sv2v_reg  <= w_data_i[131];
      \nz.mem_1000_sv2v_reg  <= w_data_i[130];
      \nz.mem_999_sv2v_reg  <= w_data_i[129];
      \nz.mem_998_sv2v_reg  <= w_data_i[128];
      \nz.mem_997_sv2v_reg  <= w_data_i[127];
      \nz.mem_996_sv2v_reg  <= w_data_i[126];
      \nz.mem_995_sv2v_reg  <= w_data_i[125];
      \nz.mem_994_sv2v_reg  <= w_data_i[124];
      \nz.mem_993_sv2v_reg  <= w_data_i[123];
      \nz.mem_992_sv2v_reg  <= w_data_i[122];
      \nz.mem_991_sv2v_reg  <= w_data_i[121];
      \nz.mem_990_sv2v_reg  <= w_data_i[120];
      \nz.mem_989_sv2v_reg  <= w_data_i[119];
      \nz.mem_988_sv2v_reg  <= w_data_i[118];
      \nz.mem_987_sv2v_reg  <= w_data_i[117];
      \nz.mem_986_sv2v_reg  <= w_data_i[116];
      \nz.mem_985_sv2v_reg  <= w_data_i[115];
      \nz.mem_984_sv2v_reg  <= w_data_i[114];
      \nz.mem_983_sv2v_reg  <= w_data_i[113];
      \nz.mem_982_sv2v_reg  <= w_data_i[112];
      \nz.mem_981_sv2v_reg  <= w_data_i[111];
      \nz.mem_980_sv2v_reg  <= w_data_i[110];
      \nz.mem_979_sv2v_reg  <= w_data_i[109];
      \nz.mem_978_sv2v_reg  <= w_data_i[108];
      \nz.mem_977_sv2v_reg  <= w_data_i[107];
      \nz.mem_976_sv2v_reg  <= w_data_i[106];
      \nz.mem_975_sv2v_reg  <= w_data_i[105];
      \nz.mem_974_sv2v_reg  <= w_data_i[104];
      \nz.mem_973_sv2v_reg  <= w_data_i[103];
      \nz.mem_972_sv2v_reg  <= w_data_i[102];
      \nz.mem_971_sv2v_reg  <= w_data_i[101];
      \nz.mem_970_sv2v_reg  <= w_data_i[100];
      \nz.mem_969_sv2v_reg  <= w_data_i[99];
      \nz.mem_968_sv2v_reg  <= w_data_i[98];
      \nz.mem_967_sv2v_reg  <= w_data_i[97];
      \nz.mem_966_sv2v_reg  <= w_data_i[96];
      \nz.mem_965_sv2v_reg  <= w_data_i[95];
      \nz.mem_964_sv2v_reg  <= w_data_i[94];
      \nz.mem_963_sv2v_reg  <= w_data_i[93];
      \nz.mem_962_sv2v_reg  <= w_data_i[92];
      \nz.mem_961_sv2v_reg  <= w_data_i[91];
      \nz.mem_960_sv2v_reg  <= w_data_i[90];
      \nz.mem_959_sv2v_reg  <= w_data_i[89];
      \nz.mem_958_sv2v_reg  <= w_data_i[88];
      \nz.mem_957_sv2v_reg  <= w_data_i[87];
      \nz.mem_956_sv2v_reg  <= w_data_i[86];
      \nz.mem_955_sv2v_reg  <= w_data_i[85];
      \nz.mem_954_sv2v_reg  <= w_data_i[84];
      \nz.mem_953_sv2v_reg  <= w_data_i[83];
      \nz.mem_952_sv2v_reg  <= w_data_i[82];
      \nz.mem_951_sv2v_reg  <= w_data_i[81];
      \nz.mem_950_sv2v_reg  <= w_data_i[80];
      \nz.mem_949_sv2v_reg  <= w_data_i[79];
      \nz.mem_948_sv2v_reg  <= w_data_i[78];
      \nz.mem_947_sv2v_reg  <= w_data_i[77];
      \nz.mem_946_sv2v_reg  <= w_data_i[76];
      \nz.mem_945_sv2v_reg  <= w_data_i[75];
      \nz.mem_870_sv2v_reg  <= w_data_i[0];
    end 
    if(N45) begin
      \nz.mem_944_sv2v_reg  <= w_data_i[74];
      \nz.mem_943_sv2v_reg  <= w_data_i[73];
      \nz.mem_942_sv2v_reg  <= w_data_i[72];
      \nz.mem_941_sv2v_reg  <= w_data_i[71];
      \nz.mem_940_sv2v_reg  <= w_data_i[70];
      \nz.mem_939_sv2v_reg  <= w_data_i[69];
      \nz.mem_938_sv2v_reg  <= w_data_i[68];
      \nz.mem_937_sv2v_reg  <= w_data_i[67];
      \nz.mem_936_sv2v_reg  <= w_data_i[66];
      \nz.mem_935_sv2v_reg  <= w_data_i[65];
      \nz.mem_934_sv2v_reg  <= w_data_i[64];
      \nz.mem_933_sv2v_reg  <= w_data_i[63];
      \nz.mem_932_sv2v_reg  <= w_data_i[62];
      \nz.mem_931_sv2v_reg  <= w_data_i[61];
      \nz.mem_930_sv2v_reg  <= w_data_i[60];
      \nz.mem_929_sv2v_reg  <= w_data_i[59];
      \nz.mem_928_sv2v_reg  <= w_data_i[58];
      \nz.mem_927_sv2v_reg  <= w_data_i[57];
      \nz.mem_926_sv2v_reg  <= w_data_i[56];
      \nz.mem_925_sv2v_reg  <= w_data_i[55];
      \nz.mem_924_sv2v_reg  <= w_data_i[54];
      \nz.mem_923_sv2v_reg  <= w_data_i[53];
      \nz.mem_922_sv2v_reg  <= w_data_i[52];
      \nz.mem_921_sv2v_reg  <= w_data_i[51];
      \nz.mem_920_sv2v_reg  <= w_data_i[50];
      \nz.mem_919_sv2v_reg  <= w_data_i[49];
      \nz.mem_918_sv2v_reg  <= w_data_i[48];
      \nz.mem_917_sv2v_reg  <= w_data_i[47];
      \nz.mem_916_sv2v_reg  <= w_data_i[46];
      \nz.mem_915_sv2v_reg  <= w_data_i[45];
      \nz.mem_914_sv2v_reg  <= w_data_i[44];
      \nz.mem_913_sv2v_reg  <= w_data_i[43];
      \nz.mem_912_sv2v_reg  <= w_data_i[42];
      \nz.mem_911_sv2v_reg  <= w_data_i[41];
      \nz.mem_910_sv2v_reg  <= w_data_i[40];
      \nz.mem_909_sv2v_reg  <= w_data_i[39];
      \nz.mem_908_sv2v_reg  <= w_data_i[38];
      \nz.mem_907_sv2v_reg  <= w_data_i[37];
      \nz.mem_906_sv2v_reg  <= w_data_i[36];
      \nz.mem_905_sv2v_reg  <= w_data_i[35];
      \nz.mem_904_sv2v_reg  <= w_data_i[34];
      \nz.mem_903_sv2v_reg  <= w_data_i[33];
      \nz.mem_902_sv2v_reg  <= w_data_i[32];
      \nz.mem_901_sv2v_reg  <= w_data_i[31];
      \nz.mem_900_sv2v_reg  <= w_data_i[30];
      \nz.mem_899_sv2v_reg  <= w_data_i[29];
      \nz.mem_898_sv2v_reg  <= w_data_i[28];
      \nz.mem_897_sv2v_reg  <= w_data_i[27];
      \nz.mem_896_sv2v_reg  <= w_data_i[26];
      \nz.mem_895_sv2v_reg  <= w_data_i[25];
      \nz.mem_894_sv2v_reg  <= w_data_i[24];
      \nz.mem_893_sv2v_reg  <= w_data_i[23];
      \nz.mem_892_sv2v_reg  <= w_data_i[22];
      \nz.mem_891_sv2v_reg  <= w_data_i[21];
      \nz.mem_890_sv2v_reg  <= w_data_i[20];
      \nz.mem_889_sv2v_reg  <= w_data_i[19];
      \nz.mem_888_sv2v_reg  <= w_data_i[18];
      \nz.mem_887_sv2v_reg  <= w_data_i[17];
      \nz.mem_886_sv2v_reg  <= w_data_i[16];
      \nz.mem_885_sv2v_reg  <= w_data_i[15];
      \nz.mem_884_sv2v_reg  <= w_data_i[14];
      \nz.mem_883_sv2v_reg  <= w_data_i[13];
      \nz.mem_882_sv2v_reg  <= w_data_i[12];
      \nz.mem_881_sv2v_reg  <= w_data_i[11];
      \nz.mem_880_sv2v_reg  <= w_data_i[10];
      \nz.mem_879_sv2v_reg  <= w_data_i[9];
      \nz.mem_878_sv2v_reg  <= w_data_i[8];
      \nz.mem_877_sv2v_reg  <= w_data_i[7];
      \nz.mem_876_sv2v_reg  <= w_data_i[6];
      \nz.mem_875_sv2v_reg  <= w_data_i[5];
      \nz.mem_874_sv2v_reg  <= w_data_i[4];
      \nz.mem_873_sv2v_reg  <= w_data_i[3];
      \nz.mem_872_sv2v_reg  <= w_data_i[2];
      \nz.mem_871_sv2v_reg  <= w_data_i[1];
    end 
    if(N42) begin
      \nz.mem_869_sv2v_reg  <= w_data_i[173];
      \nz.mem_868_sv2v_reg  <= w_data_i[172];
      \nz.mem_867_sv2v_reg  <= w_data_i[171];
      \nz.mem_866_sv2v_reg  <= w_data_i[170];
      \nz.mem_865_sv2v_reg  <= w_data_i[169];
      \nz.mem_864_sv2v_reg  <= w_data_i[168];
      \nz.mem_863_sv2v_reg  <= w_data_i[167];
      \nz.mem_862_sv2v_reg  <= w_data_i[166];
      \nz.mem_861_sv2v_reg  <= w_data_i[165];
      \nz.mem_860_sv2v_reg  <= w_data_i[164];
      \nz.mem_859_sv2v_reg  <= w_data_i[163];
      \nz.mem_858_sv2v_reg  <= w_data_i[162];
      \nz.mem_857_sv2v_reg  <= w_data_i[161];
      \nz.mem_856_sv2v_reg  <= w_data_i[160];
      \nz.mem_855_sv2v_reg  <= w_data_i[159];
      \nz.mem_854_sv2v_reg  <= w_data_i[158];
      \nz.mem_853_sv2v_reg  <= w_data_i[157];
      \nz.mem_852_sv2v_reg  <= w_data_i[156];
      \nz.mem_851_sv2v_reg  <= w_data_i[155];
      \nz.mem_850_sv2v_reg  <= w_data_i[154];
      \nz.mem_849_sv2v_reg  <= w_data_i[153];
      \nz.mem_848_sv2v_reg  <= w_data_i[152];
      \nz.mem_847_sv2v_reg  <= w_data_i[151];
      \nz.mem_846_sv2v_reg  <= w_data_i[150];
      \nz.mem_845_sv2v_reg  <= w_data_i[149];
      \nz.mem_844_sv2v_reg  <= w_data_i[148];
      \nz.mem_843_sv2v_reg  <= w_data_i[147];
      \nz.mem_842_sv2v_reg  <= w_data_i[146];
      \nz.mem_841_sv2v_reg  <= w_data_i[145];
      \nz.mem_840_sv2v_reg  <= w_data_i[144];
      \nz.mem_839_sv2v_reg  <= w_data_i[143];
      \nz.mem_838_sv2v_reg  <= w_data_i[142];
      \nz.mem_837_sv2v_reg  <= w_data_i[141];
      \nz.mem_836_sv2v_reg  <= w_data_i[140];
      \nz.mem_835_sv2v_reg  <= w_data_i[139];
      \nz.mem_834_sv2v_reg  <= w_data_i[138];
      \nz.mem_833_sv2v_reg  <= w_data_i[137];
      \nz.mem_832_sv2v_reg  <= w_data_i[136];
      \nz.mem_831_sv2v_reg  <= w_data_i[135];
      \nz.mem_830_sv2v_reg  <= w_data_i[134];
      \nz.mem_829_sv2v_reg  <= w_data_i[133];
      \nz.mem_828_sv2v_reg  <= w_data_i[132];
      \nz.mem_827_sv2v_reg  <= w_data_i[131];
      \nz.mem_826_sv2v_reg  <= w_data_i[130];
      \nz.mem_825_sv2v_reg  <= w_data_i[129];
      \nz.mem_824_sv2v_reg  <= w_data_i[128];
      \nz.mem_823_sv2v_reg  <= w_data_i[127];
      \nz.mem_822_sv2v_reg  <= w_data_i[126];
      \nz.mem_821_sv2v_reg  <= w_data_i[125];
      \nz.mem_820_sv2v_reg  <= w_data_i[124];
      \nz.mem_819_sv2v_reg  <= w_data_i[123];
      \nz.mem_818_sv2v_reg  <= w_data_i[122];
      \nz.mem_817_sv2v_reg  <= w_data_i[121];
      \nz.mem_816_sv2v_reg  <= w_data_i[120];
      \nz.mem_815_sv2v_reg  <= w_data_i[119];
      \nz.mem_814_sv2v_reg  <= w_data_i[118];
      \nz.mem_813_sv2v_reg  <= w_data_i[117];
      \nz.mem_812_sv2v_reg  <= w_data_i[116];
      \nz.mem_811_sv2v_reg  <= w_data_i[115];
      \nz.mem_810_sv2v_reg  <= w_data_i[114];
      \nz.mem_809_sv2v_reg  <= w_data_i[113];
      \nz.mem_808_sv2v_reg  <= w_data_i[112];
      \nz.mem_807_sv2v_reg  <= w_data_i[111];
      \nz.mem_806_sv2v_reg  <= w_data_i[110];
      \nz.mem_805_sv2v_reg  <= w_data_i[109];
      \nz.mem_804_sv2v_reg  <= w_data_i[108];
      \nz.mem_803_sv2v_reg  <= w_data_i[107];
      \nz.mem_802_sv2v_reg  <= w_data_i[106];
      \nz.mem_801_sv2v_reg  <= w_data_i[105];
      \nz.mem_800_sv2v_reg  <= w_data_i[104];
      \nz.mem_799_sv2v_reg  <= w_data_i[103];
      \nz.mem_798_sv2v_reg  <= w_data_i[102];
      \nz.mem_797_sv2v_reg  <= w_data_i[101];
      \nz.mem_796_sv2v_reg  <= w_data_i[100];
      \nz.mem_795_sv2v_reg  <= w_data_i[99];
      \nz.mem_794_sv2v_reg  <= w_data_i[98];
      \nz.mem_793_sv2v_reg  <= w_data_i[97];
      \nz.mem_792_sv2v_reg  <= w_data_i[96];
      \nz.mem_791_sv2v_reg  <= w_data_i[95];
      \nz.mem_790_sv2v_reg  <= w_data_i[94];
      \nz.mem_789_sv2v_reg  <= w_data_i[93];
      \nz.mem_788_sv2v_reg  <= w_data_i[92];
      \nz.mem_787_sv2v_reg  <= w_data_i[91];
      \nz.mem_786_sv2v_reg  <= w_data_i[90];
      \nz.mem_785_sv2v_reg  <= w_data_i[89];
      \nz.mem_784_sv2v_reg  <= w_data_i[88];
      \nz.mem_783_sv2v_reg  <= w_data_i[87];
      \nz.mem_782_sv2v_reg  <= w_data_i[86];
      \nz.mem_781_sv2v_reg  <= w_data_i[85];
      \nz.mem_780_sv2v_reg  <= w_data_i[84];
      \nz.mem_779_sv2v_reg  <= w_data_i[83];
      \nz.mem_778_sv2v_reg  <= w_data_i[82];
      \nz.mem_777_sv2v_reg  <= w_data_i[81];
      \nz.mem_776_sv2v_reg  <= w_data_i[80];
      \nz.mem_775_sv2v_reg  <= w_data_i[79];
      \nz.mem_774_sv2v_reg  <= w_data_i[78];
      \nz.mem_773_sv2v_reg  <= w_data_i[77];
      \nz.mem_772_sv2v_reg  <= w_data_i[76];
      \nz.mem_771_sv2v_reg  <= w_data_i[75];
      \nz.mem_696_sv2v_reg  <= w_data_i[0];
    end 
    if(N43) begin
      \nz.mem_770_sv2v_reg  <= w_data_i[74];
      \nz.mem_769_sv2v_reg  <= w_data_i[73];
      \nz.mem_768_sv2v_reg  <= w_data_i[72];
      \nz.mem_767_sv2v_reg  <= w_data_i[71];
      \nz.mem_766_sv2v_reg  <= w_data_i[70];
      \nz.mem_765_sv2v_reg  <= w_data_i[69];
      \nz.mem_764_sv2v_reg  <= w_data_i[68];
      \nz.mem_763_sv2v_reg  <= w_data_i[67];
      \nz.mem_762_sv2v_reg  <= w_data_i[66];
      \nz.mem_761_sv2v_reg  <= w_data_i[65];
      \nz.mem_760_sv2v_reg  <= w_data_i[64];
      \nz.mem_759_sv2v_reg  <= w_data_i[63];
      \nz.mem_758_sv2v_reg  <= w_data_i[62];
      \nz.mem_757_sv2v_reg  <= w_data_i[61];
      \nz.mem_756_sv2v_reg  <= w_data_i[60];
      \nz.mem_755_sv2v_reg  <= w_data_i[59];
      \nz.mem_754_sv2v_reg  <= w_data_i[58];
      \nz.mem_753_sv2v_reg  <= w_data_i[57];
      \nz.mem_752_sv2v_reg  <= w_data_i[56];
      \nz.mem_751_sv2v_reg  <= w_data_i[55];
      \nz.mem_750_sv2v_reg  <= w_data_i[54];
      \nz.mem_749_sv2v_reg  <= w_data_i[53];
      \nz.mem_748_sv2v_reg  <= w_data_i[52];
      \nz.mem_747_sv2v_reg  <= w_data_i[51];
      \nz.mem_746_sv2v_reg  <= w_data_i[50];
      \nz.mem_745_sv2v_reg  <= w_data_i[49];
      \nz.mem_744_sv2v_reg  <= w_data_i[48];
      \nz.mem_743_sv2v_reg  <= w_data_i[47];
      \nz.mem_742_sv2v_reg  <= w_data_i[46];
      \nz.mem_741_sv2v_reg  <= w_data_i[45];
      \nz.mem_740_sv2v_reg  <= w_data_i[44];
      \nz.mem_739_sv2v_reg  <= w_data_i[43];
      \nz.mem_738_sv2v_reg  <= w_data_i[42];
      \nz.mem_737_sv2v_reg  <= w_data_i[41];
      \nz.mem_736_sv2v_reg  <= w_data_i[40];
      \nz.mem_735_sv2v_reg  <= w_data_i[39];
      \nz.mem_734_sv2v_reg  <= w_data_i[38];
      \nz.mem_733_sv2v_reg  <= w_data_i[37];
      \nz.mem_732_sv2v_reg  <= w_data_i[36];
      \nz.mem_731_sv2v_reg  <= w_data_i[35];
      \nz.mem_730_sv2v_reg  <= w_data_i[34];
      \nz.mem_729_sv2v_reg  <= w_data_i[33];
      \nz.mem_728_sv2v_reg  <= w_data_i[32];
      \nz.mem_727_sv2v_reg  <= w_data_i[31];
      \nz.mem_726_sv2v_reg  <= w_data_i[30];
      \nz.mem_725_sv2v_reg  <= w_data_i[29];
      \nz.mem_724_sv2v_reg  <= w_data_i[28];
      \nz.mem_723_sv2v_reg  <= w_data_i[27];
      \nz.mem_722_sv2v_reg  <= w_data_i[26];
      \nz.mem_721_sv2v_reg  <= w_data_i[25];
      \nz.mem_720_sv2v_reg  <= w_data_i[24];
      \nz.mem_719_sv2v_reg  <= w_data_i[23];
      \nz.mem_718_sv2v_reg  <= w_data_i[22];
      \nz.mem_717_sv2v_reg  <= w_data_i[21];
      \nz.mem_716_sv2v_reg  <= w_data_i[20];
      \nz.mem_715_sv2v_reg  <= w_data_i[19];
      \nz.mem_714_sv2v_reg  <= w_data_i[18];
      \nz.mem_713_sv2v_reg  <= w_data_i[17];
      \nz.mem_712_sv2v_reg  <= w_data_i[16];
      \nz.mem_711_sv2v_reg  <= w_data_i[15];
      \nz.mem_710_sv2v_reg  <= w_data_i[14];
      \nz.mem_709_sv2v_reg  <= w_data_i[13];
      \nz.mem_708_sv2v_reg  <= w_data_i[12];
      \nz.mem_707_sv2v_reg  <= w_data_i[11];
      \nz.mem_706_sv2v_reg  <= w_data_i[10];
      \nz.mem_705_sv2v_reg  <= w_data_i[9];
      \nz.mem_704_sv2v_reg  <= w_data_i[8];
      \nz.mem_703_sv2v_reg  <= w_data_i[7];
      \nz.mem_702_sv2v_reg  <= w_data_i[6];
      \nz.mem_701_sv2v_reg  <= w_data_i[5];
      \nz.mem_700_sv2v_reg  <= w_data_i[4];
      \nz.mem_699_sv2v_reg  <= w_data_i[3];
      \nz.mem_698_sv2v_reg  <= w_data_i[2];
      \nz.mem_697_sv2v_reg  <= w_data_i[1];
    end 
    if(N40) begin
      \nz.mem_695_sv2v_reg  <= w_data_i[173];
      \nz.mem_694_sv2v_reg  <= w_data_i[172];
      \nz.mem_693_sv2v_reg  <= w_data_i[171];
      \nz.mem_692_sv2v_reg  <= w_data_i[170];
      \nz.mem_691_sv2v_reg  <= w_data_i[169];
      \nz.mem_690_sv2v_reg  <= w_data_i[168];
      \nz.mem_689_sv2v_reg  <= w_data_i[167];
      \nz.mem_688_sv2v_reg  <= w_data_i[166];
      \nz.mem_687_sv2v_reg  <= w_data_i[165];
      \nz.mem_686_sv2v_reg  <= w_data_i[164];
      \nz.mem_685_sv2v_reg  <= w_data_i[163];
      \nz.mem_684_sv2v_reg  <= w_data_i[162];
      \nz.mem_683_sv2v_reg  <= w_data_i[161];
      \nz.mem_682_sv2v_reg  <= w_data_i[160];
      \nz.mem_681_sv2v_reg  <= w_data_i[159];
      \nz.mem_680_sv2v_reg  <= w_data_i[158];
      \nz.mem_679_sv2v_reg  <= w_data_i[157];
      \nz.mem_678_sv2v_reg  <= w_data_i[156];
      \nz.mem_677_sv2v_reg  <= w_data_i[155];
      \nz.mem_676_sv2v_reg  <= w_data_i[154];
      \nz.mem_675_sv2v_reg  <= w_data_i[153];
      \nz.mem_674_sv2v_reg  <= w_data_i[152];
      \nz.mem_673_sv2v_reg  <= w_data_i[151];
      \nz.mem_672_sv2v_reg  <= w_data_i[150];
      \nz.mem_671_sv2v_reg  <= w_data_i[149];
      \nz.mem_670_sv2v_reg  <= w_data_i[148];
      \nz.mem_669_sv2v_reg  <= w_data_i[147];
      \nz.mem_668_sv2v_reg  <= w_data_i[146];
      \nz.mem_667_sv2v_reg  <= w_data_i[145];
      \nz.mem_666_sv2v_reg  <= w_data_i[144];
      \nz.mem_665_sv2v_reg  <= w_data_i[143];
      \nz.mem_664_sv2v_reg  <= w_data_i[142];
      \nz.mem_663_sv2v_reg  <= w_data_i[141];
      \nz.mem_662_sv2v_reg  <= w_data_i[140];
      \nz.mem_661_sv2v_reg  <= w_data_i[139];
      \nz.mem_660_sv2v_reg  <= w_data_i[138];
      \nz.mem_659_sv2v_reg  <= w_data_i[137];
      \nz.mem_658_sv2v_reg  <= w_data_i[136];
      \nz.mem_657_sv2v_reg  <= w_data_i[135];
      \nz.mem_656_sv2v_reg  <= w_data_i[134];
      \nz.mem_655_sv2v_reg  <= w_data_i[133];
      \nz.mem_654_sv2v_reg  <= w_data_i[132];
      \nz.mem_653_sv2v_reg  <= w_data_i[131];
      \nz.mem_652_sv2v_reg  <= w_data_i[130];
      \nz.mem_651_sv2v_reg  <= w_data_i[129];
      \nz.mem_650_sv2v_reg  <= w_data_i[128];
      \nz.mem_649_sv2v_reg  <= w_data_i[127];
      \nz.mem_648_sv2v_reg  <= w_data_i[126];
      \nz.mem_647_sv2v_reg  <= w_data_i[125];
      \nz.mem_646_sv2v_reg  <= w_data_i[124];
      \nz.mem_645_sv2v_reg  <= w_data_i[123];
      \nz.mem_644_sv2v_reg  <= w_data_i[122];
      \nz.mem_643_sv2v_reg  <= w_data_i[121];
      \nz.mem_642_sv2v_reg  <= w_data_i[120];
      \nz.mem_641_sv2v_reg  <= w_data_i[119];
      \nz.mem_640_sv2v_reg  <= w_data_i[118];
      \nz.mem_639_sv2v_reg  <= w_data_i[117];
      \nz.mem_638_sv2v_reg  <= w_data_i[116];
      \nz.mem_637_sv2v_reg  <= w_data_i[115];
      \nz.mem_636_sv2v_reg  <= w_data_i[114];
      \nz.mem_635_sv2v_reg  <= w_data_i[113];
      \nz.mem_634_sv2v_reg  <= w_data_i[112];
      \nz.mem_633_sv2v_reg  <= w_data_i[111];
      \nz.mem_632_sv2v_reg  <= w_data_i[110];
      \nz.mem_631_sv2v_reg  <= w_data_i[109];
      \nz.mem_630_sv2v_reg  <= w_data_i[108];
      \nz.mem_629_sv2v_reg  <= w_data_i[107];
      \nz.mem_628_sv2v_reg  <= w_data_i[106];
      \nz.mem_627_sv2v_reg  <= w_data_i[105];
      \nz.mem_626_sv2v_reg  <= w_data_i[104];
      \nz.mem_625_sv2v_reg  <= w_data_i[103];
      \nz.mem_624_sv2v_reg  <= w_data_i[102];
      \nz.mem_623_sv2v_reg  <= w_data_i[101];
      \nz.mem_622_sv2v_reg  <= w_data_i[100];
      \nz.mem_621_sv2v_reg  <= w_data_i[99];
      \nz.mem_620_sv2v_reg  <= w_data_i[98];
      \nz.mem_619_sv2v_reg  <= w_data_i[97];
      \nz.mem_618_sv2v_reg  <= w_data_i[96];
      \nz.mem_617_sv2v_reg  <= w_data_i[95];
      \nz.mem_616_sv2v_reg  <= w_data_i[94];
      \nz.mem_615_sv2v_reg  <= w_data_i[93];
      \nz.mem_614_sv2v_reg  <= w_data_i[92];
      \nz.mem_613_sv2v_reg  <= w_data_i[91];
      \nz.mem_612_sv2v_reg  <= w_data_i[90];
      \nz.mem_611_sv2v_reg  <= w_data_i[89];
      \nz.mem_610_sv2v_reg  <= w_data_i[88];
      \nz.mem_609_sv2v_reg  <= w_data_i[87];
      \nz.mem_608_sv2v_reg  <= w_data_i[86];
      \nz.mem_607_sv2v_reg  <= w_data_i[85];
      \nz.mem_606_sv2v_reg  <= w_data_i[84];
      \nz.mem_605_sv2v_reg  <= w_data_i[83];
      \nz.mem_604_sv2v_reg  <= w_data_i[82];
      \nz.mem_603_sv2v_reg  <= w_data_i[81];
      \nz.mem_602_sv2v_reg  <= w_data_i[80];
      \nz.mem_601_sv2v_reg  <= w_data_i[79];
      \nz.mem_600_sv2v_reg  <= w_data_i[78];
      \nz.mem_599_sv2v_reg  <= w_data_i[77];
      \nz.mem_598_sv2v_reg  <= w_data_i[76];
      \nz.mem_597_sv2v_reg  <= w_data_i[75];
      \nz.mem_522_sv2v_reg  <= w_data_i[0];
    end 
    if(N41) begin
      \nz.mem_596_sv2v_reg  <= w_data_i[74];
      \nz.mem_595_sv2v_reg  <= w_data_i[73];
      \nz.mem_594_sv2v_reg  <= w_data_i[72];
      \nz.mem_593_sv2v_reg  <= w_data_i[71];
      \nz.mem_592_sv2v_reg  <= w_data_i[70];
      \nz.mem_591_sv2v_reg  <= w_data_i[69];
      \nz.mem_590_sv2v_reg  <= w_data_i[68];
      \nz.mem_589_sv2v_reg  <= w_data_i[67];
      \nz.mem_588_sv2v_reg  <= w_data_i[66];
      \nz.mem_587_sv2v_reg  <= w_data_i[65];
      \nz.mem_586_sv2v_reg  <= w_data_i[64];
      \nz.mem_585_sv2v_reg  <= w_data_i[63];
      \nz.mem_584_sv2v_reg  <= w_data_i[62];
      \nz.mem_583_sv2v_reg  <= w_data_i[61];
      \nz.mem_582_sv2v_reg  <= w_data_i[60];
      \nz.mem_581_sv2v_reg  <= w_data_i[59];
      \nz.mem_580_sv2v_reg  <= w_data_i[58];
      \nz.mem_579_sv2v_reg  <= w_data_i[57];
      \nz.mem_578_sv2v_reg  <= w_data_i[56];
      \nz.mem_577_sv2v_reg  <= w_data_i[55];
      \nz.mem_576_sv2v_reg  <= w_data_i[54];
      \nz.mem_575_sv2v_reg  <= w_data_i[53];
      \nz.mem_574_sv2v_reg  <= w_data_i[52];
      \nz.mem_573_sv2v_reg  <= w_data_i[51];
      \nz.mem_572_sv2v_reg  <= w_data_i[50];
      \nz.mem_571_sv2v_reg  <= w_data_i[49];
      \nz.mem_570_sv2v_reg  <= w_data_i[48];
      \nz.mem_569_sv2v_reg  <= w_data_i[47];
      \nz.mem_568_sv2v_reg  <= w_data_i[46];
      \nz.mem_567_sv2v_reg  <= w_data_i[45];
      \nz.mem_566_sv2v_reg  <= w_data_i[44];
      \nz.mem_565_sv2v_reg  <= w_data_i[43];
      \nz.mem_564_sv2v_reg  <= w_data_i[42];
      \nz.mem_563_sv2v_reg  <= w_data_i[41];
      \nz.mem_562_sv2v_reg  <= w_data_i[40];
      \nz.mem_561_sv2v_reg  <= w_data_i[39];
      \nz.mem_560_sv2v_reg  <= w_data_i[38];
      \nz.mem_559_sv2v_reg  <= w_data_i[37];
      \nz.mem_558_sv2v_reg  <= w_data_i[36];
      \nz.mem_557_sv2v_reg  <= w_data_i[35];
      \nz.mem_556_sv2v_reg  <= w_data_i[34];
      \nz.mem_555_sv2v_reg  <= w_data_i[33];
      \nz.mem_554_sv2v_reg  <= w_data_i[32];
      \nz.mem_553_sv2v_reg  <= w_data_i[31];
      \nz.mem_552_sv2v_reg  <= w_data_i[30];
      \nz.mem_551_sv2v_reg  <= w_data_i[29];
      \nz.mem_550_sv2v_reg  <= w_data_i[28];
      \nz.mem_549_sv2v_reg  <= w_data_i[27];
      \nz.mem_548_sv2v_reg  <= w_data_i[26];
      \nz.mem_547_sv2v_reg  <= w_data_i[25];
      \nz.mem_546_sv2v_reg  <= w_data_i[24];
      \nz.mem_545_sv2v_reg  <= w_data_i[23];
      \nz.mem_544_sv2v_reg  <= w_data_i[22];
      \nz.mem_543_sv2v_reg  <= w_data_i[21];
      \nz.mem_542_sv2v_reg  <= w_data_i[20];
      \nz.mem_541_sv2v_reg  <= w_data_i[19];
      \nz.mem_540_sv2v_reg  <= w_data_i[18];
      \nz.mem_539_sv2v_reg  <= w_data_i[17];
      \nz.mem_538_sv2v_reg  <= w_data_i[16];
      \nz.mem_537_sv2v_reg  <= w_data_i[15];
      \nz.mem_536_sv2v_reg  <= w_data_i[14];
      \nz.mem_535_sv2v_reg  <= w_data_i[13];
      \nz.mem_534_sv2v_reg  <= w_data_i[12];
      \nz.mem_533_sv2v_reg  <= w_data_i[11];
      \nz.mem_532_sv2v_reg  <= w_data_i[10];
      \nz.mem_531_sv2v_reg  <= w_data_i[9];
      \nz.mem_530_sv2v_reg  <= w_data_i[8];
      \nz.mem_529_sv2v_reg  <= w_data_i[7];
      \nz.mem_528_sv2v_reg  <= w_data_i[6];
      \nz.mem_527_sv2v_reg  <= w_data_i[5];
      \nz.mem_526_sv2v_reg  <= w_data_i[4];
      \nz.mem_525_sv2v_reg  <= w_data_i[3];
      \nz.mem_524_sv2v_reg  <= w_data_i[2];
      \nz.mem_523_sv2v_reg  <= w_data_i[1];
    end 
    if(N38) begin
      \nz.mem_521_sv2v_reg  <= w_data_i[173];
      \nz.mem_520_sv2v_reg  <= w_data_i[172];
      \nz.mem_519_sv2v_reg  <= w_data_i[171];
      \nz.mem_518_sv2v_reg  <= w_data_i[170];
      \nz.mem_517_sv2v_reg  <= w_data_i[169];
      \nz.mem_516_sv2v_reg  <= w_data_i[168];
      \nz.mem_515_sv2v_reg  <= w_data_i[167];
      \nz.mem_514_sv2v_reg  <= w_data_i[166];
      \nz.mem_513_sv2v_reg  <= w_data_i[165];
      \nz.mem_512_sv2v_reg  <= w_data_i[164];
      \nz.mem_511_sv2v_reg  <= w_data_i[163];
      \nz.mem_510_sv2v_reg  <= w_data_i[162];
      \nz.mem_509_sv2v_reg  <= w_data_i[161];
      \nz.mem_508_sv2v_reg  <= w_data_i[160];
      \nz.mem_507_sv2v_reg  <= w_data_i[159];
      \nz.mem_506_sv2v_reg  <= w_data_i[158];
      \nz.mem_505_sv2v_reg  <= w_data_i[157];
      \nz.mem_504_sv2v_reg  <= w_data_i[156];
      \nz.mem_503_sv2v_reg  <= w_data_i[155];
      \nz.mem_502_sv2v_reg  <= w_data_i[154];
      \nz.mem_501_sv2v_reg  <= w_data_i[153];
      \nz.mem_500_sv2v_reg  <= w_data_i[152];
      \nz.mem_499_sv2v_reg  <= w_data_i[151];
      \nz.mem_498_sv2v_reg  <= w_data_i[150];
      \nz.mem_497_sv2v_reg  <= w_data_i[149];
      \nz.mem_496_sv2v_reg  <= w_data_i[148];
      \nz.mem_495_sv2v_reg  <= w_data_i[147];
      \nz.mem_494_sv2v_reg  <= w_data_i[146];
      \nz.mem_493_sv2v_reg  <= w_data_i[145];
      \nz.mem_492_sv2v_reg  <= w_data_i[144];
      \nz.mem_491_sv2v_reg  <= w_data_i[143];
      \nz.mem_490_sv2v_reg  <= w_data_i[142];
      \nz.mem_489_sv2v_reg  <= w_data_i[141];
      \nz.mem_488_sv2v_reg  <= w_data_i[140];
      \nz.mem_487_sv2v_reg  <= w_data_i[139];
      \nz.mem_486_sv2v_reg  <= w_data_i[138];
      \nz.mem_485_sv2v_reg  <= w_data_i[137];
      \nz.mem_484_sv2v_reg  <= w_data_i[136];
      \nz.mem_483_sv2v_reg  <= w_data_i[135];
      \nz.mem_482_sv2v_reg  <= w_data_i[134];
      \nz.mem_481_sv2v_reg  <= w_data_i[133];
      \nz.mem_480_sv2v_reg  <= w_data_i[132];
      \nz.mem_479_sv2v_reg  <= w_data_i[131];
      \nz.mem_478_sv2v_reg  <= w_data_i[130];
      \nz.mem_477_sv2v_reg  <= w_data_i[129];
      \nz.mem_476_sv2v_reg  <= w_data_i[128];
      \nz.mem_475_sv2v_reg  <= w_data_i[127];
      \nz.mem_474_sv2v_reg  <= w_data_i[126];
      \nz.mem_473_sv2v_reg  <= w_data_i[125];
      \nz.mem_472_sv2v_reg  <= w_data_i[124];
      \nz.mem_471_sv2v_reg  <= w_data_i[123];
      \nz.mem_470_sv2v_reg  <= w_data_i[122];
      \nz.mem_469_sv2v_reg  <= w_data_i[121];
      \nz.mem_468_sv2v_reg  <= w_data_i[120];
      \nz.mem_467_sv2v_reg  <= w_data_i[119];
      \nz.mem_466_sv2v_reg  <= w_data_i[118];
      \nz.mem_465_sv2v_reg  <= w_data_i[117];
      \nz.mem_464_sv2v_reg  <= w_data_i[116];
      \nz.mem_463_sv2v_reg  <= w_data_i[115];
      \nz.mem_462_sv2v_reg  <= w_data_i[114];
      \nz.mem_461_sv2v_reg  <= w_data_i[113];
      \nz.mem_460_sv2v_reg  <= w_data_i[112];
      \nz.mem_459_sv2v_reg  <= w_data_i[111];
      \nz.mem_458_sv2v_reg  <= w_data_i[110];
      \nz.mem_457_sv2v_reg  <= w_data_i[109];
      \nz.mem_456_sv2v_reg  <= w_data_i[108];
      \nz.mem_455_sv2v_reg  <= w_data_i[107];
      \nz.mem_454_sv2v_reg  <= w_data_i[106];
      \nz.mem_453_sv2v_reg  <= w_data_i[105];
      \nz.mem_452_sv2v_reg  <= w_data_i[104];
      \nz.mem_451_sv2v_reg  <= w_data_i[103];
      \nz.mem_450_sv2v_reg  <= w_data_i[102];
      \nz.mem_449_sv2v_reg  <= w_data_i[101];
      \nz.mem_448_sv2v_reg  <= w_data_i[100];
      \nz.mem_447_sv2v_reg  <= w_data_i[99];
      \nz.mem_446_sv2v_reg  <= w_data_i[98];
      \nz.mem_445_sv2v_reg  <= w_data_i[97];
      \nz.mem_444_sv2v_reg  <= w_data_i[96];
      \nz.mem_443_sv2v_reg  <= w_data_i[95];
      \nz.mem_442_sv2v_reg  <= w_data_i[94];
      \nz.mem_441_sv2v_reg  <= w_data_i[93];
      \nz.mem_440_sv2v_reg  <= w_data_i[92];
      \nz.mem_439_sv2v_reg  <= w_data_i[91];
      \nz.mem_438_sv2v_reg  <= w_data_i[90];
      \nz.mem_437_sv2v_reg  <= w_data_i[89];
      \nz.mem_436_sv2v_reg  <= w_data_i[88];
      \nz.mem_435_sv2v_reg  <= w_data_i[87];
      \nz.mem_434_sv2v_reg  <= w_data_i[86];
      \nz.mem_433_sv2v_reg  <= w_data_i[85];
      \nz.mem_432_sv2v_reg  <= w_data_i[84];
      \nz.mem_431_sv2v_reg  <= w_data_i[83];
      \nz.mem_430_sv2v_reg  <= w_data_i[82];
      \nz.mem_429_sv2v_reg  <= w_data_i[81];
      \nz.mem_428_sv2v_reg  <= w_data_i[80];
      \nz.mem_427_sv2v_reg  <= w_data_i[79];
      \nz.mem_426_sv2v_reg  <= w_data_i[78];
      \nz.mem_425_sv2v_reg  <= w_data_i[77];
      \nz.mem_424_sv2v_reg  <= w_data_i[76];
      \nz.mem_423_sv2v_reg  <= w_data_i[75];
      \nz.mem_348_sv2v_reg  <= w_data_i[0];
    end 
    if(N39) begin
      \nz.mem_422_sv2v_reg  <= w_data_i[74];
      \nz.mem_421_sv2v_reg  <= w_data_i[73];
      \nz.mem_420_sv2v_reg  <= w_data_i[72];
      \nz.mem_419_sv2v_reg  <= w_data_i[71];
      \nz.mem_418_sv2v_reg  <= w_data_i[70];
      \nz.mem_417_sv2v_reg  <= w_data_i[69];
      \nz.mem_416_sv2v_reg  <= w_data_i[68];
      \nz.mem_415_sv2v_reg  <= w_data_i[67];
      \nz.mem_414_sv2v_reg  <= w_data_i[66];
      \nz.mem_413_sv2v_reg  <= w_data_i[65];
      \nz.mem_412_sv2v_reg  <= w_data_i[64];
      \nz.mem_411_sv2v_reg  <= w_data_i[63];
      \nz.mem_410_sv2v_reg  <= w_data_i[62];
      \nz.mem_409_sv2v_reg  <= w_data_i[61];
      \nz.mem_408_sv2v_reg  <= w_data_i[60];
      \nz.mem_407_sv2v_reg  <= w_data_i[59];
      \nz.mem_406_sv2v_reg  <= w_data_i[58];
      \nz.mem_405_sv2v_reg  <= w_data_i[57];
      \nz.mem_404_sv2v_reg  <= w_data_i[56];
      \nz.mem_403_sv2v_reg  <= w_data_i[55];
      \nz.mem_402_sv2v_reg  <= w_data_i[54];
      \nz.mem_401_sv2v_reg  <= w_data_i[53];
      \nz.mem_400_sv2v_reg  <= w_data_i[52];
      \nz.mem_399_sv2v_reg  <= w_data_i[51];
      \nz.mem_398_sv2v_reg  <= w_data_i[50];
      \nz.mem_397_sv2v_reg  <= w_data_i[49];
      \nz.mem_396_sv2v_reg  <= w_data_i[48];
      \nz.mem_395_sv2v_reg  <= w_data_i[47];
      \nz.mem_394_sv2v_reg  <= w_data_i[46];
      \nz.mem_393_sv2v_reg  <= w_data_i[45];
      \nz.mem_392_sv2v_reg  <= w_data_i[44];
      \nz.mem_391_sv2v_reg  <= w_data_i[43];
      \nz.mem_390_sv2v_reg  <= w_data_i[42];
      \nz.mem_389_sv2v_reg  <= w_data_i[41];
      \nz.mem_388_sv2v_reg  <= w_data_i[40];
      \nz.mem_387_sv2v_reg  <= w_data_i[39];
      \nz.mem_386_sv2v_reg  <= w_data_i[38];
      \nz.mem_385_sv2v_reg  <= w_data_i[37];
      \nz.mem_384_sv2v_reg  <= w_data_i[36];
      \nz.mem_383_sv2v_reg  <= w_data_i[35];
      \nz.mem_382_sv2v_reg  <= w_data_i[34];
      \nz.mem_381_sv2v_reg  <= w_data_i[33];
      \nz.mem_380_sv2v_reg  <= w_data_i[32];
      \nz.mem_379_sv2v_reg  <= w_data_i[31];
      \nz.mem_378_sv2v_reg  <= w_data_i[30];
      \nz.mem_377_sv2v_reg  <= w_data_i[29];
      \nz.mem_376_sv2v_reg  <= w_data_i[28];
      \nz.mem_375_sv2v_reg  <= w_data_i[27];
      \nz.mem_374_sv2v_reg  <= w_data_i[26];
      \nz.mem_373_sv2v_reg  <= w_data_i[25];
      \nz.mem_372_sv2v_reg  <= w_data_i[24];
      \nz.mem_371_sv2v_reg  <= w_data_i[23];
      \nz.mem_370_sv2v_reg  <= w_data_i[22];
      \nz.mem_369_sv2v_reg  <= w_data_i[21];
      \nz.mem_368_sv2v_reg  <= w_data_i[20];
      \nz.mem_367_sv2v_reg  <= w_data_i[19];
      \nz.mem_366_sv2v_reg  <= w_data_i[18];
      \nz.mem_365_sv2v_reg  <= w_data_i[17];
      \nz.mem_364_sv2v_reg  <= w_data_i[16];
      \nz.mem_363_sv2v_reg  <= w_data_i[15];
      \nz.mem_362_sv2v_reg  <= w_data_i[14];
      \nz.mem_361_sv2v_reg  <= w_data_i[13];
      \nz.mem_360_sv2v_reg  <= w_data_i[12];
      \nz.mem_359_sv2v_reg  <= w_data_i[11];
      \nz.mem_358_sv2v_reg  <= w_data_i[10];
      \nz.mem_357_sv2v_reg  <= w_data_i[9];
      \nz.mem_356_sv2v_reg  <= w_data_i[8];
      \nz.mem_355_sv2v_reg  <= w_data_i[7];
      \nz.mem_354_sv2v_reg  <= w_data_i[6];
      \nz.mem_353_sv2v_reg  <= w_data_i[5];
      \nz.mem_352_sv2v_reg  <= w_data_i[4];
      \nz.mem_351_sv2v_reg  <= w_data_i[3];
      \nz.mem_350_sv2v_reg  <= w_data_i[2];
      \nz.mem_349_sv2v_reg  <= w_data_i[1];
    end 
    if(N36) begin
      \nz.mem_347_sv2v_reg  <= w_data_i[173];
      \nz.mem_346_sv2v_reg  <= w_data_i[172];
      \nz.mem_345_sv2v_reg  <= w_data_i[171];
      \nz.mem_344_sv2v_reg  <= w_data_i[170];
      \nz.mem_343_sv2v_reg  <= w_data_i[169];
      \nz.mem_342_sv2v_reg  <= w_data_i[168];
      \nz.mem_341_sv2v_reg  <= w_data_i[167];
      \nz.mem_340_sv2v_reg  <= w_data_i[166];
      \nz.mem_339_sv2v_reg  <= w_data_i[165];
      \nz.mem_338_sv2v_reg  <= w_data_i[164];
      \nz.mem_337_sv2v_reg  <= w_data_i[163];
      \nz.mem_336_sv2v_reg  <= w_data_i[162];
      \nz.mem_335_sv2v_reg  <= w_data_i[161];
      \nz.mem_334_sv2v_reg  <= w_data_i[160];
      \nz.mem_333_sv2v_reg  <= w_data_i[159];
      \nz.mem_332_sv2v_reg  <= w_data_i[158];
      \nz.mem_331_sv2v_reg  <= w_data_i[157];
      \nz.mem_330_sv2v_reg  <= w_data_i[156];
      \nz.mem_329_sv2v_reg  <= w_data_i[155];
      \nz.mem_328_sv2v_reg  <= w_data_i[154];
      \nz.mem_327_sv2v_reg  <= w_data_i[153];
      \nz.mem_326_sv2v_reg  <= w_data_i[152];
      \nz.mem_325_sv2v_reg  <= w_data_i[151];
      \nz.mem_324_sv2v_reg  <= w_data_i[150];
      \nz.mem_323_sv2v_reg  <= w_data_i[149];
      \nz.mem_322_sv2v_reg  <= w_data_i[148];
      \nz.mem_321_sv2v_reg  <= w_data_i[147];
      \nz.mem_320_sv2v_reg  <= w_data_i[146];
      \nz.mem_319_sv2v_reg  <= w_data_i[145];
      \nz.mem_318_sv2v_reg  <= w_data_i[144];
      \nz.mem_317_sv2v_reg  <= w_data_i[143];
      \nz.mem_316_sv2v_reg  <= w_data_i[142];
      \nz.mem_315_sv2v_reg  <= w_data_i[141];
      \nz.mem_314_sv2v_reg  <= w_data_i[140];
      \nz.mem_313_sv2v_reg  <= w_data_i[139];
      \nz.mem_312_sv2v_reg  <= w_data_i[138];
      \nz.mem_311_sv2v_reg  <= w_data_i[137];
      \nz.mem_310_sv2v_reg  <= w_data_i[136];
      \nz.mem_309_sv2v_reg  <= w_data_i[135];
      \nz.mem_308_sv2v_reg  <= w_data_i[134];
      \nz.mem_307_sv2v_reg  <= w_data_i[133];
      \nz.mem_306_sv2v_reg  <= w_data_i[132];
      \nz.mem_305_sv2v_reg  <= w_data_i[131];
      \nz.mem_304_sv2v_reg  <= w_data_i[130];
      \nz.mem_303_sv2v_reg  <= w_data_i[129];
      \nz.mem_302_sv2v_reg  <= w_data_i[128];
      \nz.mem_301_sv2v_reg  <= w_data_i[127];
      \nz.mem_300_sv2v_reg  <= w_data_i[126];
      \nz.mem_299_sv2v_reg  <= w_data_i[125];
      \nz.mem_298_sv2v_reg  <= w_data_i[124];
      \nz.mem_297_sv2v_reg  <= w_data_i[123];
      \nz.mem_296_sv2v_reg  <= w_data_i[122];
      \nz.mem_295_sv2v_reg  <= w_data_i[121];
      \nz.mem_294_sv2v_reg  <= w_data_i[120];
      \nz.mem_293_sv2v_reg  <= w_data_i[119];
      \nz.mem_292_sv2v_reg  <= w_data_i[118];
      \nz.mem_291_sv2v_reg  <= w_data_i[117];
      \nz.mem_290_sv2v_reg  <= w_data_i[116];
      \nz.mem_289_sv2v_reg  <= w_data_i[115];
      \nz.mem_288_sv2v_reg  <= w_data_i[114];
      \nz.mem_287_sv2v_reg  <= w_data_i[113];
      \nz.mem_286_sv2v_reg  <= w_data_i[112];
      \nz.mem_285_sv2v_reg  <= w_data_i[111];
      \nz.mem_284_sv2v_reg  <= w_data_i[110];
      \nz.mem_283_sv2v_reg  <= w_data_i[109];
      \nz.mem_282_sv2v_reg  <= w_data_i[108];
      \nz.mem_281_sv2v_reg  <= w_data_i[107];
      \nz.mem_280_sv2v_reg  <= w_data_i[106];
      \nz.mem_279_sv2v_reg  <= w_data_i[105];
      \nz.mem_278_sv2v_reg  <= w_data_i[104];
      \nz.mem_277_sv2v_reg  <= w_data_i[103];
      \nz.mem_276_sv2v_reg  <= w_data_i[102];
      \nz.mem_275_sv2v_reg  <= w_data_i[101];
      \nz.mem_274_sv2v_reg  <= w_data_i[100];
      \nz.mem_273_sv2v_reg  <= w_data_i[99];
      \nz.mem_272_sv2v_reg  <= w_data_i[98];
      \nz.mem_271_sv2v_reg  <= w_data_i[97];
      \nz.mem_270_sv2v_reg  <= w_data_i[96];
      \nz.mem_269_sv2v_reg  <= w_data_i[95];
      \nz.mem_268_sv2v_reg  <= w_data_i[94];
      \nz.mem_267_sv2v_reg  <= w_data_i[93];
      \nz.mem_266_sv2v_reg  <= w_data_i[92];
      \nz.mem_265_sv2v_reg  <= w_data_i[91];
      \nz.mem_264_sv2v_reg  <= w_data_i[90];
      \nz.mem_263_sv2v_reg  <= w_data_i[89];
      \nz.mem_262_sv2v_reg  <= w_data_i[88];
      \nz.mem_261_sv2v_reg  <= w_data_i[87];
      \nz.mem_260_sv2v_reg  <= w_data_i[86];
      \nz.mem_259_sv2v_reg  <= w_data_i[85];
      \nz.mem_258_sv2v_reg  <= w_data_i[84];
      \nz.mem_257_sv2v_reg  <= w_data_i[83];
      \nz.mem_256_sv2v_reg  <= w_data_i[82];
      \nz.mem_255_sv2v_reg  <= w_data_i[81];
      \nz.mem_254_sv2v_reg  <= w_data_i[80];
      \nz.mem_253_sv2v_reg  <= w_data_i[79];
      \nz.mem_252_sv2v_reg  <= w_data_i[78];
      \nz.mem_251_sv2v_reg  <= w_data_i[77];
      \nz.mem_250_sv2v_reg  <= w_data_i[76];
      \nz.mem_249_sv2v_reg  <= w_data_i[75];
      \nz.mem_174_sv2v_reg  <= w_data_i[0];
    end 
    if(N37) begin
      \nz.mem_248_sv2v_reg  <= w_data_i[74];
      \nz.mem_247_sv2v_reg  <= w_data_i[73];
      \nz.mem_246_sv2v_reg  <= w_data_i[72];
      \nz.mem_245_sv2v_reg  <= w_data_i[71];
      \nz.mem_244_sv2v_reg  <= w_data_i[70];
      \nz.mem_243_sv2v_reg  <= w_data_i[69];
      \nz.mem_242_sv2v_reg  <= w_data_i[68];
      \nz.mem_241_sv2v_reg  <= w_data_i[67];
      \nz.mem_240_sv2v_reg  <= w_data_i[66];
      \nz.mem_239_sv2v_reg  <= w_data_i[65];
      \nz.mem_238_sv2v_reg  <= w_data_i[64];
      \nz.mem_237_sv2v_reg  <= w_data_i[63];
      \nz.mem_236_sv2v_reg  <= w_data_i[62];
      \nz.mem_235_sv2v_reg  <= w_data_i[61];
      \nz.mem_234_sv2v_reg  <= w_data_i[60];
      \nz.mem_233_sv2v_reg  <= w_data_i[59];
      \nz.mem_232_sv2v_reg  <= w_data_i[58];
      \nz.mem_231_sv2v_reg  <= w_data_i[57];
      \nz.mem_230_sv2v_reg  <= w_data_i[56];
      \nz.mem_229_sv2v_reg  <= w_data_i[55];
      \nz.mem_228_sv2v_reg  <= w_data_i[54];
      \nz.mem_227_sv2v_reg  <= w_data_i[53];
      \nz.mem_226_sv2v_reg  <= w_data_i[52];
      \nz.mem_225_sv2v_reg  <= w_data_i[51];
      \nz.mem_224_sv2v_reg  <= w_data_i[50];
      \nz.mem_223_sv2v_reg  <= w_data_i[49];
      \nz.mem_222_sv2v_reg  <= w_data_i[48];
      \nz.mem_221_sv2v_reg  <= w_data_i[47];
      \nz.mem_220_sv2v_reg  <= w_data_i[46];
      \nz.mem_219_sv2v_reg  <= w_data_i[45];
      \nz.mem_218_sv2v_reg  <= w_data_i[44];
      \nz.mem_217_sv2v_reg  <= w_data_i[43];
      \nz.mem_216_sv2v_reg  <= w_data_i[42];
      \nz.mem_215_sv2v_reg  <= w_data_i[41];
      \nz.mem_214_sv2v_reg  <= w_data_i[40];
      \nz.mem_213_sv2v_reg  <= w_data_i[39];
      \nz.mem_212_sv2v_reg  <= w_data_i[38];
      \nz.mem_211_sv2v_reg  <= w_data_i[37];
      \nz.mem_210_sv2v_reg  <= w_data_i[36];
      \nz.mem_209_sv2v_reg  <= w_data_i[35];
      \nz.mem_208_sv2v_reg  <= w_data_i[34];
      \nz.mem_207_sv2v_reg  <= w_data_i[33];
      \nz.mem_206_sv2v_reg  <= w_data_i[32];
      \nz.mem_205_sv2v_reg  <= w_data_i[31];
      \nz.mem_204_sv2v_reg  <= w_data_i[30];
      \nz.mem_203_sv2v_reg  <= w_data_i[29];
      \nz.mem_202_sv2v_reg  <= w_data_i[28];
      \nz.mem_201_sv2v_reg  <= w_data_i[27];
      \nz.mem_200_sv2v_reg  <= w_data_i[26];
      \nz.mem_199_sv2v_reg  <= w_data_i[25];
      \nz.mem_198_sv2v_reg  <= w_data_i[24];
      \nz.mem_197_sv2v_reg  <= w_data_i[23];
      \nz.mem_196_sv2v_reg  <= w_data_i[22];
      \nz.mem_195_sv2v_reg  <= w_data_i[21];
      \nz.mem_194_sv2v_reg  <= w_data_i[20];
      \nz.mem_193_sv2v_reg  <= w_data_i[19];
      \nz.mem_192_sv2v_reg  <= w_data_i[18];
      \nz.mem_191_sv2v_reg  <= w_data_i[17];
      \nz.mem_190_sv2v_reg  <= w_data_i[16];
      \nz.mem_189_sv2v_reg  <= w_data_i[15];
      \nz.mem_188_sv2v_reg  <= w_data_i[14];
      \nz.mem_187_sv2v_reg  <= w_data_i[13];
      \nz.mem_186_sv2v_reg  <= w_data_i[12];
      \nz.mem_185_sv2v_reg  <= w_data_i[11];
      \nz.mem_184_sv2v_reg  <= w_data_i[10];
      \nz.mem_183_sv2v_reg  <= w_data_i[9];
      \nz.mem_182_sv2v_reg  <= w_data_i[8];
      \nz.mem_181_sv2v_reg  <= w_data_i[7];
      \nz.mem_180_sv2v_reg  <= w_data_i[6];
      \nz.mem_179_sv2v_reg  <= w_data_i[5];
      \nz.mem_178_sv2v_reg  <= w_data_i[4];
      \nz.mem_177_sv2v_reg  <= w_data_i[3];
      \nz.mem_176_sv2v_reg  <= w_data_i[2];
      \nz.mem_175_sv2v_reg  <= w_data_i[1];
    end 
    if(N34) begin
      \nz.mem_173_sv2v_reg  <= w_data_i[173];
      \nz.mem_172_sv2v_reg  <= w_data_i[172];
      \nz.mem_171_sv2v_reg  <= w_data_i[171];
      \nz.mem_170_sv2v_reg  <= w_data_i[170];
      \nz.mem_169_sv2v_reg  <= w_data_i[169];
      \nz.mem_168_sv2v_reg  <= w_data_i[168];
      \nz.mem_167_sv2v_reg  <= w_data_i[167];
      \nz.mem_166_sv2v_reg  <= w_data_i[166];
      \nz.mem_165_sv2v_reg  <= w_data_i[165];
      \nz.mem_164_sv2v_reg  <= w_data_i[164];
      \nz.mem_163_sv2v_reg  <= w_data_i[163];
      \nz.mem_162_sv2v_reg  <= w_data_i[162];
      \nz.mem_161_sv2v_reg  <= w_data_i[161];
      \nz.mem_160_sv2v_reg  <= w_data_i[160];
      \nz.mem_159_sv2v_reg  <= w_data_i[159];
      \nz.mem_158_sv2v_reg  <= w_data_i[158];
      \nz.mem_157_sv2v_reg  <= w_data_i[157];
      \nz.mem_156_sv2v_reg  <= w_data_i[156];
      \nz.mem_155_sv2v_reg  <= w_data_i[155];
      \nz.mem_154_sv2v_reg  <= w_data_i[154];
      \nz.mem_153_sv2v_reg  <= w_data_i[153];
      \nz.mem_152_sv2v_reg  <= w_data_i[152];
      \nz.mem_151_sv2v_reg  <= w_data_i[151];
      \nz.mem_150_sv2v_reg  <= w_data_i[150];
      \nz.mem_149_sv2v_reg  <= w_data_i[149];
      \nz.mem_148_sv2v_reg  <= w_data_i[148];
      \nz.mem_147_sv2v_reg  <= w_data_i[147];
      \nz.mem_146_sv2v_reg  <= w_data_i[146];
      \nz.mem_145_sv2v_reg  <= w_data_i[145];
      \nz.mem_144_sv2v_reg  <= w_data_i[144];
      \nz.mem_143_sv2v_reg  <= w_data_i[143];
      \nz.mem_142_sv2v_reg  <= w_data_i[142];
      \nz.mem_141_sv2v_reg  <= w_data_i[141];
      \nz.mem_140_sv2v_reg  <= w_data_i[140];
      \nz.mem_139_sv2v_reg  <= w_data_i[139];
      \nz.mem_138_sv2v_reg  <= w_data_i[138];
      \nz.mem_137_sv2v_reg  <= w_data_i[137];
      \nz.mem_136_sv2v_reg  <= w_data_i[136];
      \nz.mem_135_sv2v_reg  <= w_data_i[135];
      \nz.mem_134_sv2v_reg  <= w_data_i[134];
      \nz.mem_133_sv2v_reg  <= w_data_i[133];
      \nz.mem_132_sv2v_reg  <= w_data_i[132];
      \nz.mem_131_sv2v_reg  <= w_data_i[131];
      \nz.mem_130_sv2v_reg  <= w_data_i[130];
      \nz.mem_129_sv2v_reg  <= w_data_i[129];
      \nz.mem_128_sv2v_reg  <= w_data_i[128];
      \nz.mem_127_sv2v_reg  <= w_data_i[127];
      \nz.mem_126_sv2v_reg  <= w_data_i[126];
      \nz.mem_125_sv2v_reg  <= w_data_i[125];
      \nz.mem_124_sv2v_reg  <= w_data_i[124];
      \nz.mem_123_sv2v_reg  <= w_data_i[123];
      \nz.mem_122_sv2v_reg  <= w_data_i[122];
      \nz.mem_121_sv2v_reg  <= w_data_i[121];
      \nz.mem_120_sv2v_reg  <= w_data_i[120];
      \nz.mem_119_sv2v_reg  <= w_data_i[119];
      \nz.mem_118_sv2v_reg  <= w_data_i[118];
      \nz.mem_117_sv2v_reg  <= w_data_i[117];
      \nz.mem_116_sv2v_reg  <= w_data_i[116];
      \nz.mem_115_sv2v_reg  <= w_data_i[115];
      \nz.mem_114_sv2v_reg  <= w_data_i[114];
      \nz.mem_113_sv2v_reg  <= w_data_i[113];
      \nz.mem_112_sv2v_reg  <= w_data_i[112];
      \nz.mem_111_sv2v_reg  <= w_data_i[111];
      \nz.mem_110_sv2v_reg  <= w_data_i[110];
      \nz.mem_109_sv2v_reg  <= w_data_i[109];
      \nz.mem_108_sv2v_reg  <= w_data_i[108];
      \nz.mem_107_sv2v_reg  <= w_data_i[107];
      \nz.mem_106_sv2v_reg  <= w_data_i[106];
      \nz.mem_105_sv2v_reg  <= w_data_i[105];
      \nz.mem_104_sv2v_reg  <= w_data_i[104];
      \nz.mem_103_sv2v_reg  <= w_data_i[103];
      \nz.mem_102_sv2v_reg  <= w_data_i[102];
      \nz.mem_101_sv2v_reg  <= w_data_i[101];
      \nz.mem_100_sv2v_reg  <= w_data_i[100];
      \nz.mem_99_sv2v_reg  <= w_data_i[99];
      \nz.mem_98_sv2v_reg  <= w_data_i[98];
      \nz.mem_97_sv2v_reg  <= w_data_i[97];
      \nz.mem_96_sv2v_reg  <= w_data_i[96];
      \nz.mem_95_sv2v_reg  <= w_data_i[95];
      \nz.mem_94_sv2v_reg  <= w_data_i[94];
      \nz.mem_93_sv2v_reg  <= w_data_i[93];
      \nz.mem_92_sv2v_reg  <= w_data_i[92];
      \nz.mem_91_sv2v_reg  <= w_data_i[91];
      \nz.mem_90_sv2v_reg  <= w_data_i[90];
      \nz.mem_89_sv2v_reg  <= w_data_i[89];
      \nz.mem_88_sv2v_reg  <= w_data_i[88];
      \nz.mem_87_sv2v_reg  <= w_data_i[87];
      \nz.mem_86_sv2v_reg  <= w_data_i[86];
      \nz.mem_85_sv2v_reg  <= w_data_i[85];
      \nz.mem_84_sv2v_reg  <= w_data_i[84];
      \nz.mem_83_sv2v_reg  <= w_data_i[83];
      \nz.mem_82_sv2v_reg  <= w_data_i[82];
      \nz.mem_81_sv2v_reg  <= w_data_i[81];
      \nz.mem_80_sv2v_reg  <= w_data_i[80];
      \nz.mem_79_sv2v_reg  <= w_data_i[79];
      \nz.mem_78_sv2v_reg  <= w_data_i[78];
      \nz.mem_77_sv2v_reg  <= w_data_i[77];
      \nz.mem_76_sv2v_reg  <= w_data_i[76];
      \nz.mem_75_sv2v_reg  <= w_data_i[75];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
    if(N35) begin
      \nz.mem_74_sv2v_reg  <= w_data_i[74];
      \nz.mem_73_sv2v_reg  <= w_data_i[73];
      \nz.mem_72_sv2v_reg  <= w_data_i[72];
      \nz.mem_71_sv2v_reg  <= w_data_i[71];
      \nz.mem_70_sv2v_reg  <= w_data_i[70];
      \nz.mem_69_sv2v_reg  <= w_data_i[69];
      \nz.mem_68_sv2v_reg  <= w_data_i[68];
      \nz.mem_67_sv2v_reg  <= w_data_i[67];
      \nz.mem_66_sv2v_reg  <= w_data_i[66];
      \nz.mem_65_sv2v_reg  <= w_data_i[65];
      \nz.mem_64_sv2v_reg  <= w_data_i[64];
      \nz.mem_63_sv2v_reg  <= w_data_i[63];
      \nz.mem_62_sv2v_reg  <= w_data_i[62];
      \nz.mem_61_sv2v_reg  <= w_data_i[61];
      \nz.mem_60_sv2v_reg  <= w_data_i[60];
      \nz.mem_59_sv2v_reg  <= w_data_i[59];
      \nz.mem_58_sv2v_reg  <= w_data_i[58];
      \nz.mem_57_sv2v_reg  <= w_data_i[57];
      \nz.mem_56_sv2v_reg  <= w_data_i[56];
      \nz.mem_55_sv2v_reg  <= w_data_i[55];
      \nz.mem_54_sv2v_reg  <= w_data_i[54];
      \nz.mem_53_sv2v_reg  <= w_data_i[53];
      \nz.mem_52_sv2v_reg  <= w_data_i[52];
      \nz.mem_51_sv2v_reg  <= w_data_i[51];
      \nz.mem_50_sv2v_reg  <= w_data_i[50];
      \nz.mem_49_sv2v_reg  <= w_data_i[49];
      \nz.mem_48_sv2v_reg  <= w_data_i[48];
      \nz.mem_47_sv2v_reg  <= w_data_i[47];
      \nz.mem_46_sv2v_reg  <= w_data_i[46];
      \nz.mem_45_sv2v_reg  <= w_data_i[45];
      \nz.mem_44_sv2v_reg  <= w_data_i[44];
      \nz.mem_43_sv2v_reg  <= w_data_i[43];
      \nz.mem_42_sv2v_reg  <= w_data_i[42];
      \nz.mem_41_sv2v_reg  <= w_data_i[41];
      \nz.mem_40_sv2v_reg  <= w_data_i[40];
      \nz.mem_39_sv2v_reg  <= w_data_i[39];
      \nz.mem_38_sv2v_reg  <= w_data_i[38];
      \nz.mem_37_sv2v_reg  <= w_data_i[37];
      \nz.mem_36_sv2v_reg  <= w_data_i[36];
      \nz.mem_35_sv2v_reg  <= w_data_i[35];
      \nz.mem_34_sv2v_reg  <= w_data_i[34];
      \nz.mem_33_sv2v_reg  <= w_data_i[33];
      \nz.mem_32_sv2v_reg  <= w_data_i[32];
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
    end 
  end


endmodule



module bsg_mem_1r1w_000000ae_00000008
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [2:0] w_addr_i;
  input [173:0] w_data_i;
  input [2:0] r_addr_i;
  output [173:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [173:0] r_data_o;

  bsg_mem_1r1w_synth_000000ae_00000008_0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bp_be_instr_decoder_00
(
  preissue_pkt_i,
  decode_info_i,
  decode_o,
  illegal_instr_o,
  ecall_m_o,
  ecall_s_o,
  ecall_u_o,
  ebreak_o,
  dbreak_o,
  dret_o,
  mret_o,
  sret_o,
  wfi_o,
  sfence_vma_o,
  fencei_o,
  csrw_o,
  imm_o
);

  input [38:0] preissue_pkt_i;
  input [12:0] decode_info_i;
  output [53:0] decode_o;
  output [63:0] imm_o;
  output illegal_instr_o;
  output ecall_m_o;
  output ecall_s_o;
  output ecall_u_o;
  output ebreak_o;
  output dbreak_o;
  output dret_o;
  output mret_o;
  output sret_o;
  output wfi_o;
  output sfence_vma_o;
  output fencei_o;
  output csrw_o;
  wire [53:0] decode_o;
  wire [63:0] imm_o;
  wire illegal_instr_o,ecall_m_o,ecall_s_o,ecall_u_o,ebreak_o,dbreak_o,dret_o,mret_o,
  sret_o,wfi_o,sfence_vma_o,fencei_o,csrw_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,
  N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,
  N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,
  N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,
  N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,
  N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,
  N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,
  N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,
  N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,
  N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,
  decode_o_45_,decode_o_44_,decode_o_43_,decode_o_42_,decode_o_41_,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,
  N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,
  N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,
  N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,
  N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,
  N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,
  N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,
  N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
  N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,
  N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
  N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,
  N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,
  N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,
  N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,
  N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,
  N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,
  N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,
  N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,
  N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,
  N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,
  N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,
  N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,
  N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,
  N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,
  N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,
  N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,
  N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,
  N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,
  N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,
  N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,
  N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,
  N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,
  N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,
  N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
  N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,
  N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,
  N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,
  N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,
  N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,
  N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,
  N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,
  N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,
  N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,
  N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,
  N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,
  N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,
  N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,
  N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,
  N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,
  N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,
  N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,
  N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,
  N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,
  N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,
  N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,
  N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,
  N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,
  N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,
  N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,
  N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,
  N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,
  N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,
  N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,
  N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,
  N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,
  N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,
  N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,
  N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,
  N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,
  N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,
  N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,
  N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,
  N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,
  N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,
  N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,
  N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,
  N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,
  N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,
  N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,
  N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,
  N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,
  N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,
  N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,
  N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
  N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,
  N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,
  N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,
  N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,
  N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,
  N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,
  N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,
  N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,
  N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,
  N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,
  N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,
  N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,
  N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,
  N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,
  N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,
  N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,
  N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,
  N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,
  N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,
  N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,
  N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,
  N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,
  N1754,N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,
  N1767,N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,
  N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,
  N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,
  N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,
  N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,
  N1834,N1835,N1836,N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,
  N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,
  N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,
  N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,
  N1887,N1888,N1889,N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,
  N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,
  N1914,N1915,N1916,N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,
  N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,
  N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,
  N1954,N1955,N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,
  N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,
  N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,
  N1994,N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,
  N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,
  N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,
  N2034,N2035,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,
  N2047,N2048,N2049,N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,
  N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,
  N2074,N2075,N2076,N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,
  N2087,N2088,N2089,N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,
  N2100,N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,
  N2114,N2115,N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,
  N2127,N2128,N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,
  N2140,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,
  N2154,N2155,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,
  N2167,N2168,N2169,N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,
  N2180,N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,
  N2194,N2195,N2196,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,
  N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,
  N2220,N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,
  N2234,N2235,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,
  N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,
  N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,
  N2274,N2275,N2276,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,
  N2287,N2288,N2289,N2290,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,
  N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,
  N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,
  N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,
  N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,
  N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,
  N2367,N2368,N2369,N2370,N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,
  N2380,N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,
  N2394,N2395,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,
  N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,
  N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,
  N2434,N2435,N2436,N2437,N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,
  N2447,N2448,N2449,N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,
  N2460,N2461,N2462,N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,
  N2474,N2475,N2476,N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,
  N2487,N2488,N2489,N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,
  N2500,N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,
  N2514,N2515,N2516,N2517,N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,
  N2527,N2528,N2529,N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,
  N2540,N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,
  N2554,N2555,N2556,N2557,N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,
  N2567,N2568,N2569,N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,
  N2580,N2581,N2582,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,
  N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,
  N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,
  N2620,N2621,N2622,N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,
  N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,
  N2647,N2648,N2649,N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,
  N2660,N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,
  N2674,N2675,N2676,N2677,N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,
  N2687,N2688,N2689,N2690,N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,
  N2700,N2701,N2702,N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,
  N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,
  N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,
  N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,
  N2754,N2755,N2756,N2757,N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,
  N2767,N2768,N2769,N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,
  N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,
  N2794,N2795,N2796,N2797,N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,
  N2807,N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,N2819,
  N2820,N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,
  N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,
  N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,N2859,
  N2860,N2861,N2862,N2863,N2864,N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,
  N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,
  N2887,N2888,N2889,N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,
  N2900,N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908;
  assign decode_o[7] = 1'b0;
  assign decode_o[19] = 1'b0;
  assign decode_o[31] = 1'b0;
  assign decode_o_45_ = preissue_pkt_i[38];
  assign decode_o[45] = decode_o_45_;
  assign decode_o_44_ = preissue_pkt_i[37];
  assign decode_o[44] = decode_o_44_;
  assign decode_o_43_ = preissue_pkt_i[36];
  assign decode_o[43] = decode_o_43_;
  assign decode_o_42_ = preissue_pkt_i[35];
  assign decode_o[42] = decode_o_42_;
  assign decode_o_41_ = preissue_pkt_i[34];
  assign decode_o[41] = decode_o_41_;
  assign N173 = preissue_pkt_i[3] & preissue_pkt_i[2];
  assign N175 = N188 | preissue_pkt_i[4];
  assign N176 = N187 | N183;
  assign N177 = N176 | preissue_pkt_i[4];
  assign N179 = preissue_pkt_i[8] | preissue_pkt_i[7];
  assign N180 = N203 | preissue_pkt_i[5];
  assign N181 = N179 | N180;
  assign N182 = N181 | preissue_pkt_i[4];
  assign N183 = N203 | N204;
  assign N184 = N179 | N183;
  assign N185 = N184 | preissue_pkt_i[4];
  assign N187 = preissue_pkt_i[8] | N202;
  assign N188 = N187 | N180;
  assign N189 = N188 | N205;
  assign N191 = N181 | N205;
  assign N193 = N197 | N235;
  assign N194 = N193 | N205;
  assign N195 = N198 | N205;
  assign N197 = N201 | N202;
  assign N198 = N197 | N212;
  assign N199 = N198 | preissue_pkt_i[4];
  assign N206 = N201 & N202;
  assign N207 = N203 & N204;
  assign N208 = N206 & N207;
  assign N209 = N208 & N205;
  assign N210 = N2568 | N205;
  assign N212 = preissue_pkt_i[6] | preissue_pkt_i[5];
  assign N213 = N187 | N212;
  assign N214 = N213 | preissue_pkt_i[4];
  assign N216 = N213 | N205;
  assign N218 = N179 | N235;
  assign N219 = N218 | N205;
  assign N221 = N197 | N180;
  assign N222 = N221 | preissue_pkt_i[4];
  assign N224 = N201 | preissue_pkt_i[7];
  assign N225 = N224 | N180;
  assign N226 = N225 | preissue_pkt_i[4];
  assign N228 = N224 | N212;
  assign N229 = N228 | preissue_pkt_i[4];
  assign N230 = N228 | N205;
  assign N231 = N224 | N235;
  assign N232 = N231 | preissue_pkt_i[4];
  assign N233 = N231 | N205;
  assign N235 = preissue_pkt_i[6] | N204;
  assign N236 = N187 | N235;
  assign N237 = N236 | N205;
  assign N239 = preissue_pkt_i[6] & preissue_pkt_i[5];
  assign N240 = N239 & preissue_pkt_i[4];
  assign N241 = preissue_pkt_i[8] & preissue_pkt_i[6];
  assign N242 = N241 & preissue_pkt_i[4];
  assign N243 = N241 & preissue_pkt_i[5];
  assign N244 = preissue_pkt_i[7] & N203;
  assign N245 = preissue_pkt_i[5] & N205;
  assign N246 = N244 & N245;
  assign N247 = N201 & N203;
  assign N248 = N247 & N245;
  assign N250 = preissue_pkt_i[16] | N526;
  assign N251 = preissue_pkt_i[15] | N250;
  assign N252 = preissue_pkt_i[14] | N251;
  assign N253 = preissue_pkt_i[8] | N252;
  assign N254 = N1328 | N253;
  assign N255 = N394 | N254;
  assign N256 = preissue_pkt_i[5] | N255;
  assign N257 = preissue_pkt_i[4] | N256;
  assign N258 = N395 | N257;
  assign N259 = N396 | N258;
  assign N260 = ~N259;
  assign N261 = N1329 | N255;
  assign N262 = preissue_pkt_i[4] | N261;
  assign N263 = N395 | N262;
  assign N264 = N396 | N263;
  assign N265 = ~N264;
  assign N266 = N260 | N265;
  assign N267 = N2305 | N251;
  assign N268 = preissue_pkt_i[8] | N267;
  assign N269 = N1328 | N268;
  assign N270 = N394 | N269;
  assign N271 = preissue_pkt_i[5] | N270;
  assign N272 = preissue_pkt_i[4] | N271;
  assign N273 = N395 | N272;
  assign N274 = N396 | N273;
  assign N275 = ~N274;
  assign N276 = N394 | N483;
  assign N277 = preissue_pkt_i[5] | N276;
  assign N278 = preissue_pkt_i[4] | N277;
  assign N279 = N395 | N278;
  assign N280 = N396 | N279;
  assign N281 = ~N280;
  assign N282 = N275 | N281;
  assign N283 = N394 | N492;
  assign N284 = preissue_pkt_i[5] | N283;
  assign N285 = preissue_pkt_i[4] | N284;
  assign N286 = N395 | N285;
  assign N287 = N396 | N286;
  assign N288 = ~N287;
  assign N289 = N282 | N288;
  assign N290 = preissue_pkt_i[5] | N305;
  assign N291 = preissue_pkt_i[4] | N290;
  assign N292 = N395 | N291;
  assign N293 = N396 | N292;
  assign N294 = ~N293;
  assign N295 = N289 | N294;
  assign N296 = preissue_pkt_i[5] | N312;
  assign N297 = preissue_pkt_i[4] | N296;
  assign N298 = N395 | N297;
  assign N299 = N396 | N298;
  assign N300 = ~N299;
  assign N301 = N295 | N300;
  assign N302 = preissue_pkt_i[14] | N506;
  assign N303 = preissue_pkt_i[8] | N302;
  assign N304 = N1328 | N303;
  assign N305 = N394 | N304;
  assign N306 = N1329 | N305;
  assign N307 = preissue_pkt_i[4] | N306;
  assign N308 = N395 | N307;
  assign N309 = N396 | N308;
  assign N310 = ~N309;
  assign N311 = N301 | N310;
  assign N312 = N394 | N509;
  assign N313 = N1329 | N312;
  assign N314 = preissue_pkt_i[4] | N313;
  assign N315 = N395 | N314;
  assign N316 = N396 | N315;
  assign N317 = ~N316;
  assign N318 = N311 | N317;
  assign N319 = preissue_pkt_i[5] | N334;
  assign N320 = preissue_pkt_i[4] | N319;
  assign N321 = N395 | N320;
  assign N322 = N396 | N321;
  assign N323 = ~N322;
  assign N324 = N318 | N323;
  assign N325 = preissue_pkt_i[5] | N341;
  assign N326 = preissue_pkt_i[4] | N325;
  assign N327 = N395 | N326;
  assign N328 = N396 | N327;
  assign N329 = ~N328;
  assign N330 = N324 | N329;
  assign N331 = preissue_pkt_i[14] | N528;
  assign N332 = preissue_pkt_i[8] | N331;
  assign N333 = N1328 | N332;
  assign N334 = N394 | N333;
  assign N335 = N1329 | N334;
  assign N336 = preissue_pkt_i[4] | N335;
  assign N337 = N395 | N336;
  assign N338 = N396 | N337;
  assign N339 = ~N338;
  assign N340 = N330 | N339;
  assign N341 = N394 | N531;
  assign N342 = N1329 | N341;
  assign N343 = preissue_pkt_i[4] | N342;
  assign N344 = N395 | N343;
  assign N345 = N396 | N344;
  assign N346 = ~N345;
  assign N347 = N340 | N346;
  assign N350 = preissue_pkt_i[16] | N402;
  assign N351 = preissue_pkt_i[15] | N350;
  assign N352 = preissue_pkt_i[14] | N351;
  assign N353 = preissue_pkt_i[8] | N352;
  assign N354 = N1328 | N353;
  assign N355 = N394 | N354;
  assign N356 = N1329 | N355;
  assign N357 = preissue_pkt_i[4] | N356;
  assign N358 = N395 | N357;
  assign N359 = N396 | N358;
  assign N360 = ~N359;
  assign N361 = preissue_pkt_i[16] | N974;
  assign N362 = N2304 | N361;
  assign N363 = preissue_pkt_i[14] | N362;
  assign N364 = preissue_pkt_i[8] | N363;
  assign N365 = N1328 | N364;
  assign N366 = N394 | N365;
  assign N367 = N1329 | N366;
  assign N368 = preissue_pkt_i[4] | N367;
  assign N369 = N395 | N368;
  assign N370 = N396 | N369;
  assign N371 = ~N370;
  assign N372 = N360 | N371;
  assign N373 = preissue_pkt_i[15] | N975;
  assign N374 = preissue_pkt_i[14] | N373;
  assign N375 = preissue_pkt_i[8] | N374;
  assign N376 = N1328 | N375;
  assign N377 = N394 | N376;
  assign N378 = N1329 | N377;
  assign N379 = preissue_pkt_i[4] | N378;
  assign N380 = N395 | N379;
  assign N381 = N396 | N380;
  assign N382 = ~N381;
  assign N383 = N372 | N382;
  assign N384 = N394 | N979;
  assign N385 = N1329 | N384;
  assign N386 = preissue_pkt_i[4] | N385;
  assign N387 = N395 | N386;
  assign N388 = N396 | N387;
  assign N389 = ~N388;
  assign N390 = N383 | N389;
  assign N393 = ~preissue_pkt_i[29];
  assign N394 = ~preissue_pkt_i[6];
  assign N395 = ~preissue_pkt_i[3];
  assign N396 = ~preissue_pkt_i[2];
  assign N397 = preissue_pkt_i[32] | preissue_pkt_i[33];
  assign N398 = preissue_pkt_i[31] | N397;
  assign N399 = preissue_pkt_i[30] | N398;
  assign N400 = N393 | N399;
  assign N401 = preissue_pkt_i[28] | N400;
  assign N402 = preissue_pkt_i[27] | N401;
  assign N403 = N1631 | N402;
  assign N404 = preissue_pkt_i[15] | N403;
  assign N405 = preissue_pkt_i[14] | N404;
  assign N406 = preissue_pkt_i[8] | N405;
  assign N407 = N1328 | N406;
  assign N408 = N394 | N407;
  assign N409 = N1329 | N408;
  assign N410 = preissue_pkt_i[4] | N409;
  assign N411 = N395 | N410;
  assign N412 = N396 | N411;
  assign N413 = ~N412;
  assign N415 = N288 | N300;
  assign N416 = N415 | N317;
  assign N417 = N416 | N329;
  assign N418 = N417 | N346;
  assign N419 = preissue_pkt_i[5] | N425;
  assign N420 = preissue_pkt_i[4] | N419;
  assign N421 = N395 | N420;
  assign N422 = N396 | N421;
  assign N423 = ~N422;
  assign N424 = N418 | N423;
  assign N425 = N394 | N860;
  assign N426 = N1329 | N425;
  assign N427 = preissue_pkt_i[4] | N426;
  assign N428 = N395 | N427;
  assign N429 = N396 | N428;
  assign N430 = ~N429;
  assign N431 = N424 | N430;
  assign N432 = N431 | N360;
  assign N433 = N432 | N371;
  assign N434 = N433 | N382;
  assign N435 = N434 | N389;
  assign N436 = N394 | N407;
  assign N437 = N1329 | N436;
  assign N438 = preissue_pkt_i[4] | N437;
  assign N439 = N395 | N438;
  assign N440 = N396 | N439;
  assign N441 = ~N440;
  assign N442 = N435 | N441;
  assign N443 = preissue_pkt_i[5] | N449;
  assign N444 = preissue_pkt_i[4] | N443;
  assign N445 = N395 | N444;
  assign N446 = N396 | N445;
  assign N447 = ~N446;
  assign N448 = N442 | N447;
  assign N449 = N394 | N914;
  assign N450 = N1329 | N449;
  assign N451 = preissue_pkt_i[4] | N450;
  assign N452 = N395 | N451;
  assign N453 = N396 | N452;
  assign N454 = ~N453;
  assign N455 = N448 | N454;
  assign N456 = preissue_pkt_i[5] | N473;
  assign N457 = preissue_pkt_i[4] | N456;
  assign N458 = N395 | N457;
  assign N459 = N396 | N458;
  assign N460 = ~N459;
  assign N461 = N455 | N460;
  assign N462 = ~preissue_pkt_i[31];
  assign N463 = N462 | N1288;
  assign N464 = preissue_pkt_i[30] | N463;
  assign N465 = preissue_pkt_i[29] | N464;
  assign N466 = preissue_pkt_i[28] | N465;
  assign N467 = preissue_pkt_i[27] | N466;
  assign N468 = preissue_pkt_i[16] | N467;
  assign N469 = preissue_pkt_i[15] | N468;
  assign N470 = N2305 | N469;
  assign N471 = preissue_pkt_i[8] | N470;
  assign N472 = N1328 | N471;
  assign N473 = N394 | N472;
  assign N474 = N1329 | N473;
  assign N475 = preissue_pkt_i[4] | N474;
  assign N476 = N395 | N475;
  assign N477 = N396 | N476;
  assign N478 = ~N477;
  assign N479 = N461 | N478;
  assign N480 = N2304 | N250;
  assign N481 = preissue_pkt_i[14] | N480;
  assign N482 = preissue_pkt_i[8] | N481;
  assign N483 = N1328 | N482;
  assign N484 = N394 | N483;
  assign N485 = preissue_pkt_i[5] | N484;
  assign N486 = preissue_pkt_i[4] | N485;
  assign N487 = N395 | N486;
  assign N488 = N396 | N487;
  assign N489 = ~N488;
  assign N490 = N2305 | N480;
  assign N491 = preissue_pkt_i[8] | N490;
  assign N492 = N1328 | N491;
  assign N493 = N394 | N492;
  assign N494 = preissue_pkt_i[5] | N493;
  assign N495 = preissue_pkt_i[4] | N494;
  assign N496 = N395 | N495;
  assign N497 = N396 | N496;
  assign N498 = ~N497;
  assign N499 = N489 | N498;
  assign N500 = preissue_pkt_i[5] | N510;
  assign N501 = preissue_pkt_i[4] | N500;
  assign N502 = N395 | N501;
  assign N503 = N396 | N502;
  assign N504 = ~N503;
  assign N505 = N499 | N504;
  assign N506 = preissue_pkt_i[15] | N527;
  assign N507 = N2305 | N506;
  assign N508 = preissue_pkt_i[8] | N507;
  assign N509 = N1328 | N508;
  assign N510 = N394 | N509;
  assign N511 = N1329 | N510;
  assign N512 = preissue_pkt_i[4] | N511;
  assign N513 = N395 | N512;
  assign N514 = N396 | N513;
  assign N515 = ~N514;
  assign N516 = N505 | N515;
  assign N517 = preissue_pkt_i[5] | N532;
  assign N518 = preissue_pkt_i[4] | N517;
  assign N519 = N395 | N518;
  assign N520 = N396 | N519;
  assign N521 = ~N520;
  assign N522 = N516 | N521;
  assign N523 = ~preissue_pkt_i[27];
  assign N524 = preissue_pkt_i[29] | N399;
  assign N525 = preissue_pkt_i[28] | N524;
  assign N526 = N523 | N525;
  assign N527 = N1631 | N526;
  assign N528 = N2304 | N527;
  assign N529 = N2305 | N528;
  assign N530 = preissue_pkt_i[8] | N529;
  assign N531 = N1328 | N530;
  assign N532 = N394 | N531;
  assign N533 = N1329 | N532;
  assign N534 = preissue_pkt_i[4] | N533;
  assign N535 = N395 | N534;
  assign N536 = N396 | N535;
  assign N537 = ~N536;
  assign N538 = N522 | N537;
  assign N539 = N2135 & N2303;
  assign N540 = N2684 & N1327;
  assign N541 = N1330 & preissue_pkt_i[3];
  assign N542 = N539 & N540;
  assign N543 = N2573 & N541;
  assign N544 = N542 & N543;
  assign N545 = N544 & preissue_pkt_i[2];
  assign N547 = N2305 & N1329;
  assign N548 = N617 & N547;
  assign N549 = N585 & N548;
  assign N550 = N2305 & preissue_pkt_i[5];
  assign N551 = N617 & N550;
  assign N552 = N585 & N551;
  assign N553 = N581 & N616;
  assign N554 = N553 & N551;
  assign N555 = preissue_pkt_i[32] & N462;
  assign N556 = N555 & N582;
  assign N557 = N617 & N584;
  assign N558 = N556 & N557;
  assign N559 = N617 & N697;
  assign N560 = N556 & N559;
  assign N561 = N585 & N619;
  assign N562 = N617 & N651;
  assign N563 = N585 & N562;
  assign N564 = N585 & N595;
  assign N565 = N1357 & N651;
  assign N566 = N585 & N565;
  assign N567 = N625 & N582;
  assign N568 = N567 & N586;
  assign N569 = N583 & N697;
  assign N570 = N567 & N569;
  assign N571 = N567 & N593;
  assign N572 = N1357 & N697;
  assign N573 = N567 & N572;
  assign N574 = N567 & N597;
  assign N575 = N1360 & N697;
  assign N576 = N567 & N575;
  assign N577 = N553 & N572;
  assign N578 = N556 & N595;
  assign N579 = N556 & N565;
  assign N581 = N1287 & N462;
  assign N582 = N393 & N523;
  assign N583 = N1631 & preissue_pkt_i[15];
  assign N584 = N2305 & N1329;
  assign N585 = N581 & N582;
  assign N586 = N583 & N584;
  assign N587 = N585 & N586;
  assign N588 = preissue_pkt_i[14] & N1329;
  assign N589 = N583 & N588;
  assign N590 = N585 & N589;
  assign N591 = preissue_pkt_i[29] & preissue_pkt_i[27];
  assign N592 = N581 & N591;
  assign N593 = N1357 & N584;
  assign N594 = N592 & N593;
  assign N595 = N1357 & N588;
  assign N596 = N592 & N595;
  assign N597 = N1360 & N584;
  assign N598 = N592 & N597;
  assign N599 = N1360 & N588;
  assign N600 = N592 & N599;
  assign N601 = N585 & N593;
  assign N602 = N556 & N593;
  assign N604 = N622 & N582;
  assign N605 = N604 & N619;
  assign N606 = N604 & N562;
  assign N607 = N604 & N595;
  assign N608 = N604 & N565;
  assign N609 = N585 & N597;
  assign N610 = N556 & N597;
  assign N612 = N585 & N599;
  assign N613 = N556 & N599;
  assign N615 = preissue_pkt_i[32] & N462;
  assign N616 = preissue_pkt_i[29] & N523;
  assign N617 = N1631 & N2304;
  assign N618 = N615 & N616;
  assign N619 = N617 & N588;
  assign N620 = N618 & N619;
  assign N621 = N618 & N595;
  assign N622 = preissue_pkt_i[32] & preissue_pkt_i[31];
  assign N623 = N622 & N616;
  assign N624 = N623 & N619;
  assign N625 = N1287 & preissue_pkt_i[31];
  assign N626 = N625 & N616;
  assign N627 = N626 & N619;
  assign N628 = N633 & N557;
  assign N629 = N633 & N559;
  assign N631 = N1287 & N462;
  assign N632 = N393 & preissue_pkt_i[27];
  assign N633 = N631 & N632;
  assign N634 = N633 & N619;
  assign N635 = N633 & N586;
  assign N636 = N633 & N589;
  assign N637 = N633 & N593;
  assign N638 = N633 & N572;
  assign N640 = N633 & N595;
  assign N641 = N633 & N565;
  assign N643 = N633 & N597;
  assign N644 = N633 & N575;
  assign N646 = N633 & N599;
  assign N647 = N1360 & N651;
  assign N648 = N633 & N647;
  assign N650 = N523 & preissue_pkt_i[15];
  assign N651 = preissue_pkt_i[14] & preissue_pkt_i[5];
  assign N652 = N650 & N651;
  assign N653 = N1287 & preissue_pkt_i[29];
  assign N654 = N523 & preissue_pkt_i[16];
  assign N655 = N653 & N654;
  assign N656 = N655 & preissue_pkt_i[14];
  assign N657 = preissue_pkt_i[16] & preissue_pkt_i[14];
  assign N658 = N2458 & N657;
  assign N659 = N1287 & preissue_pkt_i[31];
  assign N660 = N659 & N657;
  assign N661 = preissue_pkt_i[31] & preissue_pkt_i[15];
  assign N662 = N661 & preissue_pkt_i[14];
  assign N663 = N393 & preissue_pkt_i[14];
  assign N664 = N659 & N663;
  assign N665 = N583 & N651;
  assign N666 = N615 & N672;
  assign N667 = N666 & preissue_pkt_i[5];
  assign N668 = preissue_pkt_i[29] & preissue_pkt_i[14];
  assign N669 = N668 & preissue_pkt_i[5];
  assign N670 = preissue_pkt_i[27] & N1631;
  assign N671 = N670 & N651;
  assign N672 = N1631 & preissue_pkt_i[14];
  assign N673 = N591 & N672;
  assign N674 = N631 & N688;
  assign N675 = N674 & preissue_pkt_i[14];
  assign N676 = N393 & N1631;
  assign N677 = N615 & N676;
  assign N678 = N677 & preissue_pkt_i[14];
  assign N679 = preissue_pkt_i[29] & preissue_pkt_i[15];
  assign N680 = N679 & preissue_pkt_i[5];
  assign N681 = N616 & preissue_pkt_i[15];
  assign N682 = N622 & preissue_pkt_i[15];
  assign N683 = N462 & N523;
  assign N684 = preissue_pkt_i[15] & preissue_pkt_i[5];
  assign N685 = N683 & N684;
  assign N686 = preissue_pkt_i[32] & N1631;
  assign N687 = N686 & preissue_pkt_i[15];
  assign N688 = preissue_pkt_i[29] & N1631;
  assign N689 = N688 & preissue_pkt_i[15];
  assign N690 = N462 & N1631;
  assign N691 = N690 & N684;
  assign N692 = preissue_pkt_i[32] & preissue_pkt_i[16];
  assign N693 = N692 & N1410;
  assign N694 = N693 & preissue_pkt_i[5];
  assign N695 = N2458 & preissue_pkt_i[5];
  assign N696 = N462 & N393;
  assign N697 = N2305 & preissue_pkt_i[5];
  assign N698 = N696 & N654;
  assign N699 = N698 & N697;
  assign N700 = N591 & preissue_pkt_i[5];
  assign N701 = N2460 & preissue_pkt_i[5];
  assign N702 = preissue_pkt_i[31] & preissue_pkt_i[27];
  assign N703 = N616 & N584;
  assign N704 = N622 & N584;
  assign N705 = preissue_pkt_i[31] & N1631;
  assign N706 = N705 & N1410;
  assign N707 = N688 & N584;
  assign N708 = preissue_pkt_i[32] & preissue_pkt_i[27];
  assign N722 = preissue_pkt_i[16] | N2036;
  assign N723 = preissue_pkt_i[15] | N722;
  assign N724 = preissue_pkt_i[14] | N723;
  assign N725 = preissue_pkt_i[8] | N724;
  assign N726 = N1328 | N725;
  assign N727 = N394 | N726;
  assign N728 = preissue_pkt_i[5] | N727;
  assign N729 = preissue_pkt_i[4] | N728;
  assign N730 = N395 | N729;
  assign N731 = N396 | N730;
  assign N732 = ~N731;
  assign N733 = N1329 | N727;
  assign N734 = preissue_pkt_i[4] | N733;
  assign N735 = N395 | N734;
  assign N736 = N396 | N735;
  assign N737 = ~N736;
  assign N738 = N732 | N737;
  assign N739 = preissue_pkt_i[14] | N749;
  assign N740 = preissue_pkt_i[8] | N739;
  assign N741 = N1328 | N740;
  assign N742 = N394 | N741;
  assign N743 = preissue_pkt_i[5] | N742;
  assign N744 = preissue_pkt_i[4] | N743;
  assign N745 = N395 | N744;
  assign N746 = N396 | N745;
  assign N747 = ~N746;
  assign N748 = N738 | N747;
  assign N749 = N2304 | N836;
  assign N750 = N2305 | N749;
  assign N751 = preissue_pkt_i[8] | N750;
  assign N752 = N1328 | N751;
  assign N753 = N394 | N752;
  assign N754 = preissue_pkt_i[5] | N753;
  assign N755 = preissue_pkt_i[4] | N754;
  assign N756 = N395 | N755;
  assign N757 = N396 | N756;
  assign N758 = ~N757;
  assign N759 = N748 | N758;
  assign N760 = preissue_pkt_i[14] | N770;
  assign N761 = preissue_pkt_i[8] | N760;
  assign N762 = N1328 | N761;
  assign N763 = N394 | N762;
  assign N764 = preissue_pkt_i[5] | N763;
  assign N765 = preissue_pkt_i[4] | N764;
  assign N766 = N395 | N765;
  assign N767 = N396 | N766;
  assign N768 = ~N767;
  assign N769 = N759 | N768;
  assign N770 = preissue_pkt_i[15] | N792;
  assign N771 = N2305 | N770;
  assign N772 = preissue_pkt_i[8] | N771;
  assign N773 = N1328 | N772;
  assign N774 = N394 | N773;
  assign N775 = preissue_pkt_i[5] | N774;
  assign N776 = preissue_pkt_i[4] | N775;
  assign N777 = N395 | N776;
  assign N778 = N396 | N777;
  assign N779 = ~N778;
  assign N780 = N769 | N779;
  assign N781 = preissue_pkt_i[14] | N793;
  assign N782 = preissue_pkt_i[8] | N781;
  assign N783 = N1328 | N782;
  assign N784 = N394 | N783;
  assign N785 = preissue_pkt_i[5] | N784;
  assign N786 = preissue_pkt_i[4] | N785;
  assign N787 = N395 | N786;
  assign N788 = N396 | N787;
  assign N789 = ~N788;
  assign N790 = N780 | N789;
  assign N791 = N523 | N401;
  assign N792 = N1631 | N791;
  assign N793 = N2304 | N792;
  assign N794 = N2305 | N793;
  assign N795 = preissue_pkt_i[8] | N794;
  assign N796 = N1328 | N795;
  assign N797 = N394 | N796;
  assign N798 = preissue_pkt_i[5] | N797;
  assign N799 = preissue_pkt_i[4] | N798;
  assign N800 = N395 | N799;
  assign N801 = N396 | N800;
  assign N802 = ~N801;
  assign N803 = N790 | N802;
  assign N804 = N2304 | N879;
  assign N805 = N2305 | N804;
  assign N806 = preissue_pkt_i[8] | N805;
  assign N807 = N1328 | N806;
  assign N808 = N394 | N807;
  assign N809 = preissue_pkt_i[5] | N808;
  assign N810 = preissue_pkt_i[4] | N809;
  assign N811 = N395 | N810;
  assign N812 = N396 | N811;
  assign N813 = ~N812;
  assign N814 = preissue_pkt_i[14] | N804;
  assign N815 = preissue_pkt_i[8] | N814;
  assign N816 = N1328 | N815;
  assign N817 = N394 | N816;
  assign N818 = preissue_pkt_i[5] | N817;
  assign N819 = preissue_pkt_i[4] | N818;
  assign N820 = N395 | N819;
  assign N821 = N396 | N820;
  assign N822 = ~N821;
  assign N823 = N813 | N822;
  assign N824 = preissue_pkt_i[14] | N880;
  assign N825 = preissue_pkt_i[8] | N824;
  assign N826 = N1328 | N825;
  assign N827 = N394 | N826;
  assign N828 = preissue_pkt_i[5] | N827;
  assign N829 = preissue_pkt_i[4] | N828;
  assign N830 = N395 | N829;
  assign N831 = N396 | N830;
  assign N832 = ~N831;
  assign N833 = N823 | N832;
  assign N836 = preissue_pkt_i[16] | N1809;
  assign N837 = preissue_pkt_i[15] | N836;
  assign N838 = N2305 | N837;
  assign N839 = preissue_pkt_i[8] | N838;
  assign N840 = N1328 | N839;
  assign N841 = N394 | N840;
  assign N842 = preissue_pkt_i[5] | N841;
  assign N843 = preissue_pkt_i[4] | N842;
  assign N844 = N395 | N843;
  assign N845 = N396 | N844;
  assign N846 = ~N845;
  assign N847 = N1329 | N841;
  assign N848 = preissue_pkt_i[4] | N847;
  assign N849 = N395 | N848;
  assign N850 = N396 | N849;
  assign N851 = ~N850;
  assign N852 = N846 | N851;
  assign N856 = N1631 | N1809;
  assign N857 = preissue_pkt_i[15] | N856;
  assign N858 = N2305 | N857;
  assign N859 = preissue_pkt_i[8] | N858;
  assign N860 = N1328 | N859;
  assign N861 = N394 | N860;
  assign N862 = preissue_pkt_i[5] | N861;
  assign N863 = preissue_pkt_i[4] | N862;
  assign N864 = N395 | N863;
  assign N865 = N396 | N864;
  assign N866 = ~N865;
  assign N867 = N1329 | N861;
  assign N868 = preissue_pkt_i[4] | N867;
  assign N869 = N395 | N868;
  assign N870 = N396 | N869;
  assign N871 = ~N870;
  assign N872 = N866 | N871;
  assign N873 = preissue_pkt_i[5] | N884;
  assign N874 = preissue_pkt_i[4] | N873;
  assign N875 = N395 | N874;
  assign N876 = N396 | N875;
  assign N877 = ~N876;
  assign N878 = N872 | N877;
  assign N879 = N1631 | N2036;
  assign N880 = preissue_pkt_i[15] | N879;
  assign N881 = N2305 | N880;
  assign N882 = preissue_pkt_i[8] | N881;
  assign N883 = N1328 | N882;
  assign N884 = N394 | N883;
  assign N885 = N1329 | N884;
  assign N886 = preissue_pkt_i[4] | N885;
  assign N887 = N395 | N886;
  assign N888 = N396 | N887;
  assign N889 = ~N888;
  assign N890 = N878 | N889;
  assign N896 = N394 | N472;
  assign N897 = preissue_pkt_i[5] | N896;
  assign N898 = preissue_pkt_i[4] | N897;
  assign N899 = N395 | N898;
  assign N900 = N396 | N899;
  assign N901 = ~N900;
  assign N902 = N1329 | N896;
  assign N903 = preissue_pkt_i[4] | N902;
  assign N904 = N395 | N903;
  assign N905 = N396 | N904;
  assign N906 = ~N905;
  assign N907 = N901 | N906;
  assign N914 = N1328 | N1249;
  assign N915 = N394 | N914;
  assign N916 = preissue_pkt_i[5] | N915;
  assign N917 = preissue_pkt_i[4] | N916;
  assign N918 = N395 | N917;
  assign N919 = N396 | N918;
  assign N920 = ~N919;
  assign N921 = N1329 | N915;
  assign N922 = preissue_pkt_i[4] | N921;
  assign N923 = N395 | N922;
  assign N924 = N396 | N923;
  assign N925 = ~N924;
  assign N926 = N920 | N925;
  assign N933 = N395 | N410;
  assign N934 = N396 | N933;
  assign N935 = ~N934;
  assign N939 = N394 | N365;
  assign N940 = preissue_pkt_i[5] | N939;
  assign N941 = preissue_pkt_i[4] | N940;
  assign N942 = N395 | N941;
  assign N943 = N396 | N942;
  assign N944 = ~N943;
  assign N945 = N1329 | N939;
  assign N946 = preissue_pkt_i[4] | N945;
  assign N947 = N395 | N946;
  assign N948 = N396 | N947;
  assign N949 = ~N948;
  assign N950 = N944 | N949;
  assign N951 = preissue_pkt_i[5] | N957;
  assign N952 = preissue_pkt_i[4] | N951;
  assign N953 = N395 | N952;
  assign N954 = N396 | N953;
  assign N955 = ~N954;
  assign N956 = N950 | N955;
  assign N957 = N394 | N376;
  assign N958 = N1329 | N957;
  assign N959 = preissue_pkt_i[4] | N958;
  assign N960 = N395 | N959;
  assign N961 = N396 | N960;
  assign N962 = ~N961;
  assign N963 = N956 | N962;
  assign N964 = preissue_pkt_i[5] | N980;
  assign N965 = preissue_pkt_i[4] | N964;
  assign N966 = N395 | N965;
  assign N967 = N396 | N966;
  assign N968 = ~N967;
  assign N969 = N963 | N968;
  assign N970 = N462 | N397;
  assign N971 = preissue_pkt_i[30] | N970;
  assign N972 = preissue_pkt_i[29] | N971;
  assign N973 = preissue_pkt_i[28] | N972;
  assign N974 = preissue_pkt_i[27] | N973;
  assign N975 = N1631 | N974;
  assign N976 = N2304 | N975;
  assign N977 = preissue_pkt_i[14] | N976;
  assign N978 = preissue_pkt_i[8] | N977;
  assign N979 = N1328 | N978;
  assign N980 = N394 | N979;
  assign N981 = N1329 | N980;
  assign N982 = preissue_pkt_i[4] | N981;
  assign N983 = N395 | N982;
  assign N984 = N396 | N983;
  assign N985 = ~N984;
  assign N986 = N969 | N985;
  assign N991 = preissue_pkt_i[16] | N401;
  assign N992 = preissue_pkt_i[15] | N991;
  assign N993 = N2305 | N992;
  assign N994 = preissue_pkt_i[8] | N993;
  assign N995 = preissue_pkt_i[7] | N994;
  assign N996 = N394 | N995;
  assign N997 = N1329 | N996;
  assign N998 = preissue_pkt_i[4] | N997;
  assign N999 = N395 | N998;
  assign N1000 = N396 | N999;
  assign N1001 = ~N1000;
  assign N1003 = N1011 & N2339;
  assign N1004 = N1003 & N1016;
  assign N1005 = N1018 & N1004;
  assign N1006 = N1005 & N1020;
  assign N1007 = N2135 & preissue_pkt_i[32];
  assign N1008 = preissue_pkt_i[31] & N2303;
  assign N1009 = N393 & N2684;
  assign N1010 = N523 & N2685;
  assign N1011 = N2686 & preissue_pkt_i[24];
  assign N1012 = N2079 & preissue_pkt_i[22];
  assign N1013 = N1007 & N1008;
  assign N1014 = N1009 & N1010;
  assign N1015 = N1011 & N1012;
  assign N1016 = N1354 & N2384;
  assign N1017 = N1870 & N2290;
  assign N1018 = N1013 & N1014;
  assign N1019 = N1015 & N1016;
  assign N1020 = N1017 & N173;
  assign N1021 = N1018 & N1019;
  assign N1022 = N1021 & N1020;
  assign N1027 = preissue_pkt_i[6] & N1330;
  assign N1028 = N1426 & N1027;
  assign N1029 = N1028 & N173;
  assign N1031 = N1354 & N584;
  assign N1032 = N1354 & N697;
  assign N1033 = N462 & N2303;
  assign N1034 = N1973 & N1033;
  assign N1035 = N1009 & N1354;
  assign N1036 = N1034 & N1035;
  assign N1037 = N1036 & N588;
  assign N1038 = N1036 & N651;
  assign N1039 = N1034 & N1103;
  assign N1040 = N1039 & N651;
  assign N1041 = N1034 & N1055;
  assign N1042 = N1041 & N588;
  assign N1043 = N1041 & N651;
  assign N1044 = N1003 & N1069;
  assign N1045 = N1018 & N1044;
  assign N1046 = N1015 & N1069;
  assign N1047 = N1018 & N1046;
  assign N1048 = N1007 & N1033;
  assign N1049 = N1048 & N1055;
  assign N1050 = N1049 & N588;
  assign N1051 = N1049 & N651;
  assign N1053 = N1363 & N584;
  assign N1054 = N1363 & N588;
  assign N1055 = N1009 & N1357;
  assign N1056 = N1013 & N1055;
  assign N1057 = N1056 & N588;
  assign N1058 = N1009 & N654;
  assign N1059 = N1411 & preissue_pkt_i[5];
  assign N1060 = N1013 & N1058;
  assign N1061 = N1060 & N1059;
  assign N1063 = N1461 & N1069;
  assign N1064 = N1018 & N1063;
  assign N1065 = N1461 & N1072;
  assign N1066 = N1018 & N1065;
  assign N1068 = N2383 & N1012;
  assign N1069 = N1354 & N588;
  assign N1070 = N1068 & N1069;
  assign N1071 = N1018 & N1070;
  assign N1072 = N1354 & N651;
  assign N1073 = N1068 & N1072;
  assign N1074 = N1018 & N1073;
  assign N1075 = N2383 & N2339;
  assign N1076 = N1075 & N1069;
  assign N1077 = N1018 & N1076;
  assign N1078 = N1075 & N1072;
  assign N1079 = N1018 & N1078;
  assign N1081 = preissue_pkt_i[23] & preissue_pkt_i[22];
  assign N1082 = N1102 & N1010;
  assign N1083 = N1011 & N1081;
  assign N1084 = N1928 & N1082;
  assign N1085 = N1083 & N595;
  assign N1086 = N1084 & N1085;
  assign N1087 = preissue_pkt_i[27] & preissue_pkt_i[26];
  assign N1088 = preissue_pkt_i[25] & N1183;
  assign N1089 = N1102 & N1087;
  assign N1090 = N1088 & N2339;
  assign N1091 = N1099 & N1089;
  assign N1092 = N1090 & N595;
  assign N1093 = N1091 & N1092;
  assign N1094 = N1874 & N1103;
  assign N1095 = N1094 & N588;
  assign N1096 = N1102 & N1357;
  assign N1097 = N1874 & N1096;
  assign N1098 = N1097 & N588;
  assign N1099 = N1007 & N2005;
  assign N1100 = N1099 & N1103;
  assign N1101 = N1100 & N588;
  assign N1102 = preissue_pkt_i[29] & N2684;
  assign N1103 = N1102 & N1354;
  assign N1104 = N1928 & N1103;
  assign N1105 = N1104 & N588;
  assign N1132 = preissue_pkt_i[26] | N467;
  assign N1133 = preissue_pkt_i[25] | N1132;
  assign N1134 = preissue_pkt_i[24] | N1133;
  assign N1135 = preissue_pkt_i[23] | N1134;
  assign N1136 = N2035 | N1135;
  assign N1137 = preissue_pkt_i[16] | N1136;
  assign N1138 = preissue_pkt_i[15] | N1137;
  assign N1139 = N2305 | N1138;
  assign N1140 = preissue_pkt_i[8] | N1139;
  assign N1141 = preissue_pkt_i[7] | N1140;
  assign N1142 = N394 | N1141;
  assign N1143 = preissue_pkt_i[5] | N1142;
  assign N1144 = preissue_pkt_i[4] | N1143;
  assign N1145 = N395 | N1144;
  assign N1146 = N396 | N1145;
  assign N1147 = ~N1146;
  assign N1148 = N1329 | N1142;
  assign N1149 = preissue_pkt_i[4] | N1148;
  assign N1150 = N395 | N1149;
  assign N1151 = N396 | N1150;
  assign N1152 = ~N1151;
  assign N1153 = N1147 | N1152;
  assign N1154 = N1280 | N1001;
  assign N1155 = N2079 | N1134;
  assign N1156 = preissue_pkt_i[22] | N1155;
  assign N1157 = preissue_pkt_i[16] | N1156;
  assign N1158 = preissue_pkt_i[15] | N1157;
  assign N1159 = N2305 | N1158;
  assign N1160 = preissue_pkt_i[8] | N1159;
  assign N1161 = preissue_pkt_i[7] | N1160;
  assign N1162 = N394 | N1161;
  assign N1163 = N1329 | N1162;
  assign N1164 = preissue_pkt_i[4] | N1163;
  assign N1165 = N395 | N1164;
  assign N1166 = N396 | N1165;
  assign N1167 = ~N1166;
  assign N1168 = N1154 | N1167;
  assign N1169 = preissue_pkt_i[22] | N1135;
  assign N1170 = preissue_pkt_i[16] | N1169;
  assign N1171 = preissue_pkt_i[15] | N1170;
  assign N1172 = N2305 | N1171;
  assign N1173 = preissue_pkt_i[8] | N1172;
  assign N1174 = preissue_pkt_i[7] | N1173;
  assign N1175 = N394 | N1174;
  assign N1176 = N1329 | N1175;
  assign N1177 = preissue_pkt_i[4] | N1176;
  assign N1178 = N395 | N1177;
  assign N1179 = N396 | N1178;
  assign N1180 = ~N1179;
  assign N1181 = N1168 | N1180;
  assign N1182 = N1181 | N1152;
  assign N1183 = ~preissue_pkt_i[24];
  assign N1184 = N1183 | N1133;
  assign N1185 = preissue_pkt_i[23] | N1184;
  assign N1186 = preissue_pkt_i[22] | N1185;
  assign N1187 = preissue_pkt_i[16] | N1186;
  assign N1188 = preissue_pkt_i[15] | N1187;
  assign N1189 = N2305 | N1188;
  assign N1190 = preissue_pkt_i[8] | N1189;
  assign N1191 = preissue_pkt_i[7] | N1190;
  assign N1192 = N394 | N1191;
  assign N1193 = preissue_pkt_i[5] | N1192;
  assign N1194 = preissue_pkt_i[4] | N1193;
  assign N1195 = N395 | N1194;
  assign N1196 = N396 | N1195;
  assign N1197 = ~N1196;
  assign N1198 = N2035 | N1185;
  assign N1199 = preissue_pkt_i[16] | N1198;
  assign N1200 = preissue_pkt_i[15] | N1199;
  assign N1201 = N2305 | N1200;
  assign N1202 = preissue_pkt_i[8] | N1201;
  assign N1203 = preissue_pkt_i[7] | N1202;
  assign N1204 = N394 | N1203;
  assign N1205 = preissue_pkt_i[5] | N1204;
  assign N1206 = preissue_pkt_i[4] | N1205;
  assign N1207 = N395 | N1206;
  assign N1208 = N396 | N1207;
  assign N1209 = ~N1208;
  assign N1210 = N1197 | N1209;
  assign N1213 = preissue_pkt_i[16] | N525;
  assign N1214 = preissue_pkt_i[15] | N1213;
  assign N1215 = N2305 | N1214;
  assign N1216 = preissue_pkt_i[8] | N1215;
  assign N1217 = preissue_pkt_i[7] | N1216;
  assign N1218 = N394 | N1217;
  assign N1219 = preissue_pkt_i[5] | N1218;
  assign N1220 = preissue_pkt_i[4] | N1219;
  assign N1221 = N395 | N1220;
  assign N1222 = N396 | N1221;
  assign N1223 = ~N1222;
  assign N1224 = N1329 | N1218;
  assign N1225 = preissue_pkt_i[4] | N1224;
  assign N1226 = N395 | N1225;
  assign N1227 = N396 | N1226;
  assign N1228 = ~N1227;
  assign N1229 = N1223 | N1228;
  assign N1230 = N1229 | N1001;
  assign N1235 = N1631 | N466;
  assign N1236 = preissue_pkt_i[15] | N1235;
  assign N1237 = N2305 | N1236;
  assign N1238 = preissue_pkt_i[8] | N1237;
  assign N1239 = preissue_pkt_i[7] | N1238;
  assign N1240 = N394 | N1239;
  assign N1241 = preissue_pkt_i[5] | N1240;
  assign N1242 = preissue_pkt_i[4] | N1241;
  assign N1243 = N395 | N1242;
  assign N1244 = N396 | N1243;
  assign N1245 = ~N1244;
  assign N1246 = N1631 | N467;
  assign N1247 = preissue_pkt_i[15] | N1246;
  assign N1248 = N2305 | N1247;
  assign N1249 = preissue_pkt_i[8] | N1248;
  assign N1250 = preissue_pkt_i[7] | N1249;
  assign N1251 = N394 | N1250;
  assign N1252 = N1329 | N1251;
  assign N1253 = preissue_pkt_i[4] | N1252;
  assign N1254 = N395 | N1253;
  assign N1255 = N396 | N1254;
  assign N1256 = ~N1255;
  assign N1257 = N1245 | N1256;
  assign N1264 = N1631 | N525;
  assign N1265 = preissue_pkt_i[15] | N1264;
  assign N1266 = N2305 | N1265;
  assign N1267 = preissue_pkt_i[8] | N1266;
  assign N1268 = preissue_pkt_i[7] | N1267;
  assign N1269 = N394 | N1268;
  assign N1270 = preissue_pkt_i[5] | N1269;
  assign N1271 = preissue_pkt_i[4] | N1270;
  assign N1272 = N395 | N1271;
  assign N1273 = N396 | N1272;
  assign N1274 = ~N1273;
  assign N1275 = N1329 | N1269;
  assign N1276 = preissue_pkt_i[4] | N1275;
  assign N1277 = N395 | N1276;
  assign N1278 = N396 | N1277;
  assign N1279 = ~N1278;
  assign N1280 = N1274 | N1279;
  assign N1281 = preissue_pkt_i[5] | N1298;
  assign N1282 = preissue_pkt_i[4] | N1281;
  assign N1283 = N395 | N1282;
  assign N1284 = N396 | N1283;
  assign N1285 = ~N1284;
  assign N1286 = N1280 | N1285;
  assign N1287 = ~preissue_pkt_i[32];
  assign N1288 = N1287 | preissue_pkt_i[33];
  assign N1289 = preissue_pkt_i[31] | N1288;
  assign N1290 = preissue_pkt_i[30] | N1289;
  assign N1291 = preissue_pkt_i[29] | N1290;
  assign N1292 = preissue_pkt_i[28] | N1291;
  assign N1293 = N1631 | N1292;
  assign N1294 = preissue_pkt_i[15] | N1293;
  assign N1295 = N2305 | N1294;
  assign N1296 = preissue_pkt_i[8] | N1295;
  assign N1297 = preissue_pkt_i[7] | N1296;
  assign N1298 = N394 | N1297;
  assign N1299 = N1329 | N1298;
  assign N1300 = preissue_pkt_i[4] | N1299;
  assign N1301 = N395 | N1300;
  assign N1302 = N396 | N1301;
  assign N1303 = ~N1302;
  assign N1304 = N1286 | N1303;
  assign N1311 = N394 | N1389;
  assign N1312 = preissue_pkt_i[5] | N1311;
  assign N1313 = preissue_pkt_i[4] | N1312;
  assign N1314 = N395 | N1313;
  assign N1315 = N396 | N1314;
  assign N1316 = ~N1315;
  assign N1317 = N2305 | N1386;
  assign N1318 = preissue_pkt_i[8] | N1317;
  assign N1319 = preissue_pkt_i[7] | N1318;
  assign N1320 = N394 | N1319;
  assign N1321 = preissue_pkt_i[5] | N1320;
  assign N1322 = preissue_pkt_i[4] | N1321;
  assign N1323 = N395 | N1322;
  assign N1324 = N396 | N1323;
  assign N1325 = ~N1324;
  assign N1326 = N1316 | N1325;
  assign N1327 = ~preissue_pkt_i[8];
  assign N1328 = ~preissue_pkt_i[7];
  assign N1329 = ~preissue_pkt_i[5];
  assign N1330 = ~preissue_pkt_i[4];
  assign N1331 = N1328 | N1327;
  assign N1332 = preissue_pkt_i[6] | N1331;
  assign N1333 = N1329 | N1332;
  assign N1334 = N1330 | N1333;
  assign N1335 = N395 | N1334;
  assign N1336 = N396 | N1335;
  assign N1337 = ~N1336;
  assign N1338 = preissue_pkt_i[15] | preissue_pkt_i[16];
  assign N1339 = preissue_pkt_i[14] | N1338;
  assign N1340 = N1327 | N1339;
  assign N1341 = N1328 | N1340;
  assign N1342 = preissue_pkt_i[6] | N1341;
  assign N1343 = preissue_pkt_i[5] | N1342;
  assign N1344 = N1330 | N1343;
  assign N1345 = N395 | N1344;
  assign N1346 = N396 | N1345;
  assign N1347 = ~N1346;
  assign N1348 = N1337 | N1347;
  assign N1350 = preissue_pkt_i[4] | N395;
  assign N1351 = N1350 | N396;
  assign N1352 = N2553 | N1351;
  assign N1354 = N1631 & N2304;
  assign N1355 = N1354 & N2305;
  assign N1356 = N1354 & preissue_pkt_i[14];
  assign N1357 = preissue_pkt_i[16] & N2304;
  assign N1358 = N1357 & N2305;
  assign N1359 = N1357 & preissue_pkt_i[14];
  assign N1360 = preissue_pkt_i[16] & preissue_pkt_i[15];
  assign N1361 = N1360 & N2305;
  assign N1362 = N1360 & preissue_pkt_i[14];
  assign N1363 = N1631 & preissue_pkt_i[15];
  assign N1374 = N2568 | N1351;
  assign N1376 = N1363 & N2305;
  assign N1377 = N1363 & preissue_pkt_i[14];
  assign N1386 = N2304 | preissue_pkt_i[16];
  assign N1387 = preissue_pkt_i[14] | N1386;
  assign N1388 = preissue_pkt_i[8] | N1387;
  assign N1389 = preissue_pkt_i[7] | N1388;
  assign N1390 = preissue_pkt_i[6] | N1389;
  assign N1391 = preissue_pkt_i[5] | N1390;
  assign N1392 = N1330 | N1391;
  assign N1393 = N395 | N1392;
  assign N1394 = N396 | N1393;
  assign N1395 = ~N1394;
  assign N1396 = preissue_pkt_i[4] & preissue_pkt_i[3];
  assign N1397 = N1363 & N1426;
  assign N1398 = N2561 & N1396;
  assign N1399 = N1397 & N1398;
  assign N1400 = N1399 & preissue_pkt_i[2];
  assign N1404 = N1631 & N1327;
  assign N1405 = preissue_pkt_i[7] & N394;
  assign N1406 = N1404 & N1405;
  assign N1407 = N2290 & N173;
  assign N1408 = N1406 & N1407;
  assign N1410 = N2304 & N2305;
  assign N1411 = N2304 & preissue_pkt_i[14];
  assign N1412 = preissue_pkt_i[15] & N2305;
  assign N1413 = preissue_pkt_i[15] & preissue_pkt_i[14];
  assign N1419 = N1327 & preissue_pkt_i[7];
  assign N1420 = N1363 & N1419;
  assign N1421 = N1420 & N1398;
  assign N1422 = N1421 & preissue_pkt_i[2];
  assign N1426 = N1327 & N1328;
  assign N1427 = N1426 & N173;
  assign N1429 = N2305 & N394;
  assign N1430 = N1354 & N1429;
  assign N1431 = N1430 & N2295;
  assign N1432 = preissue_pkt_i[14] & N394;
  assign N1433 = N1354 & N1432;
  assign N1434 = N1433 & N2295;
  assign N1435 = N1075 & N1442;
  assign N1436 = N1449 & N1435;
  assign N1437 = N1436 & N1467;
  assign N1438 = N1068 & N1442;
  assign N1439 = N1449 & N1438;
  assign N1440 = N1439 & N1467;
  assign N1441 = preissue_pkt_i[14] & N1589;
  assign N1442 = N1360 & N1441;
  assign N1443 = N1461 & N1442;
  assign N1444 = N1449 & N1443;
  assign N1445 = N1444 & N1467;
  assign N1446 = N1003 & N1462;
  assign N1447 = N1449 & N1446;
  assign N1448 = N1447 & N1467;
  assign N1449 = N1976 & N1014;
  assign N1450 = N1068 & N1462;
  assign N1451 = N1449 & N1450;
  assign N1452 = N1451 & N1467;
  assign N1453 = N1075 & N1462;
  assign N1454 = N1465 & N1453;
  assign N1455 = N1454 & N1467;
  assign N1456 = preissue_pkt_i[23] & N2035;
  assign N1457 = N2305 & N1589;
  assign N1458 = N1590 & N1591;
  assign N1459 = N1592 & N1593;
  assign N1460 = N2666 & N1010;
  assign N1461 = N2383 & N1456;
  assign N1462 = N1363 & N1457;
  assign N1463 = N1458 & N1459;
  assign N1464 = N2575 & preissue_pkt_i[4];
  assign N1465 = N1976 & N1460;
  assign N1466 = N1461 & N1462;
  assign N1467 = N1463 & N1464;
  assign N1468 = N1465 & N1466;
  assign N1469 = N1468 & N1467;
  assign N1470 = N2035 & preissue_pkt_i[16];
  assign N1471 = N1470 & N1412;
  assign N1472 = N1474 & N1471;
  assign N1473 = N1472 & N1484;
  assign N1474 = N1880 & N1881;
  assign N1475 = N1474 & N1480;
  assign N1476 = N1475 & N1484;
  assign N1477 = preissue_pkt_i[22] & preissue_pkt_i[16];
  assign N1478 = N1593 & preissue_pkt_i[6];
  assign N1479 = N1880 & N1886;
  assign N1480 = N1477 & N1412;
  assign N1481 = N1594 & N1595;
  assign N1482 = N1478 & N2290;
  assign N1483 = N1479 & N1480;
  assign N1484 = N1481 & N1482;
  assign N1485 = N1483 & N1484;
  assign N1516 = N2548 | N2542;
  assign N1517 = N1516 | N1351;
  assign N1524 = N1519 & N1520;
  assign N1525 = N1521 & N1522;
  assign N1526 = N1523 & N1631;
  assign N1527 = N1524 & N1525;
  assign N1528 = N1526 & N1410;
  assign N1529 = N1075 & N1527;
  assign N1530 = N1528 & N1481;
  assign N1531 = N1465 & N1529;
  assign N1532 = N1530 & N1593;
  assign N1533 = N1531 & N1532;
  assign N1534 = preissue_pkt_i[31] | preissue_pkt_i[30];
  assign N1535 = N1564 | N1534;
  assign N1536 = N1557 | N1569;
  assign N1537 = N1535 | N1577;
  assign N1538 = N1536 | N1579;
  assign N1539 = N1537 | N1538;
  assign N1540 = N1539 | N1586;
  assign N1542 = preissue_pkt_i[33] | N1287;
  assign N1543 = N393 | preissue_pkt_i[28];
  assign N1544 = N523 | N2685;
  assign N1545 = N1542 | N1551;
  assign N1546 = N1543 | N1544;
  assign N1547 = N1545 | N1546;
  assign N1548 = N1547 | N1560;
  assign N1549 = N1548 | N1586;
  assign N1551 = N462 | N2303;
  assign N1552 = N1564 | N1551;
  assign N1553 = N1552 | N1577;
  assign N1554 = N1553 | N1560;
  assign N1555 = N1554 | N1586;
  assign N1557 = preissue_pkt_i[25] | preissue_pkt_i[24];
  assign N1558 = N2079 | preissue_pkt_i[22];
  assign N1559 = N1557 | N1558;
  assign N1560 = N1559 | N1579;
  assign N1561 = N1582 | N1560;
  assign N1562 = N1561 | N1586;
  assign N1564 = preissue_pkt_i[33] | preissue_pkt_i[32];
  assign N1565 = preissue_pkt_i[31] | N2303;
  assign N1566 = preissue_pkt_i[29] | preissue_pkt_i[28];
  assign N1567 = preissue_pkt_i[27] | preissue_pkt_i[26];
  assign N1568 = preissue_pkt_i[25] | N1183;
  assign N1569 = preissue_pkt_i[23] | N2035;
  assign N1570 = preissue_pkt_i[21] | preissue_pkt_i[20];
  assign N1571 = preissue_pkt_i[19] | preissue_pkt_i[18];
  assign N1572 = preissue_pkt_i[17] | preissue_pkt_i[16];
  assign N1573 = preissue_pkt_i[15] | preissue_pkt_i[14];
  assign N1574 = preissue_pkt_i[13] | preissue_pkt_i[12];
  assign N1575 = preissue_pkt_i[11] | preissue_pkt_i[10];
  assign N1576 = N1564 | N1565;
  assign N1577 = N1566 | N1567;
  assign N1578 = N1568 | N1569;
  assign N1579 = N1570 | N1571;
  assign N1580 = N1572 | N1573;
  assign N1581 = N1574 | N1575;
  assign N1582 = N1576 | N1577;
  assign N1583 = N1578 | N1579;
  assign N1584 = N1580 | N1581;
  assign N1585 = N1582 | N1583;
  assign N1586 = N1584 | preissue_pkt_i[9];
  assign N1587 = N1585 | N1586;
  assign N1594 = N1589 & N1590;
  assign N1595 = N1591 & N1592;
  assign N1596 = N1973 & N1986;
  assign N1597 = N2666 & N670;
  assign N1598 = N1410 & N1594;
  assign N1599 = N1595 & N1593;
  assign N1600 = N1596 & N1597;
  assign N1601 = N1598 & N1599;
  assign N1602 = N1600 & N1601;
  assign N1622 = N2305 | N1338;
  assign N1623 = N1327 | N1622;
  assign N1624 = N1328 | N1623;
  assign N1625 = N394 | N1624;
  assign N1626 = preissue_pkt_i[5] | N1625;
  assign N1627 = preissue_pkt_i[4] | N1626;
  assign N1628 = N395 | N1627;
  assign N1629 = N396 | N1628;
  assign N1630 = ~N1629;
  assign N1631 = ~preissue_pkt_i[16];
  assign N1632 = preissue_pkt_i[15] | N1631;
  assign N1633 = N2305 | N1632;
  assign N1634 = N1327 | N1633;
  assign N1635 = N1328 | N1634;
  assign N1636 = N394 | N1635;
  assign N1637 = preissue_pkt_i[5] | N1636;
  assign N1638 = preissue_pkt_i[4] | N1637;
  assign N1639 = N395 | N1638;
  assign N1640 = N396 | N1639;
  assign N1641 = ~N1640;
  assign N1642 = N1630 | N1641;
  assign N1644 = N2079 | N2035;
  assign N1645 = N1557 | N1644;
  assign N1646 = N1537 | N1645;
  assign N1647 = N1537 | N1536;
  assign N1648 = N1537 | N1559;
  assign N1650 = N1654 | N1659;
  assign N1652 = N2135 | N1287;
  assign N1653 = N1652 | N1534;
  assign N1654 = N1653 | N1577;
  assign N1655 = N1654 | N1559;
  assign N1657 = preissue_pkt_i[23] | preissue_pkt_i[22];
  assign N1658 = N1543 | N1567;
  assign N1659 = N1557 | N1657;
  assign N1660 = N1576 | N1658;
  assign N1661 = N1660 | N1659;
  assign N1706 = preissue_pkt_i[15] | N361;
  assign N1707 = preissue_pkt_i[14] | N1706;
  assign N1708 = N1327 | N1707;
  assign N1709 = preissue_pkt_i[7] | N1708;
  assign N1710 = N394 | N1709;
  assign N1711 = preissue_pkt_i[5] | N1710;
  assign N1712 = preissue_pkt_i[4] | N1711;
  assign N1713 = N395 | N1712;
  assign N1714 = N396 | N1713;
  assign N1715 = ~N1714;
  assign N1716 = N2305 | N1706;
  assign N1717 = N1327 | N1716;
  assign N1718 = preissue_pkt_i[7] | N1717;
  assign N1719 = N394 | N1718;
  assign N1720 = preissue_pkt_i[5] | N1719;
  assign N1721 = preissue_pkt_i[4] | N1720;
  assign N1722 = N395 | N1721;
  assign N1723 = N396 | N1722;
  assign N1724 = ~N1723;
  assign N1725 = N1715 | N1724;
  assign N1726 = N1327 | N363;
  assign N1727 = preissue_pkt_i[7] | N1726;
  assign N1728 = N394 | N1727;
  assign N1729 = preissue_pkt_i[5] | N1728;
  assign N1730 = preissue_pkt_i[4] | N1729;
  assign N1731 = N395 | N1730;
  assign N1732 = N396 | N1731;
  assign N1733 = ~N1732;
  assign N1734 = N1725 | N1733;
  assign N1735 = preissue_pkt_i[14] | N1749;
  assign N1736 = N1327 | N1735;
  assign N1737 = preissue_pkt_i[7] | N1736;
  assign N1738 = N394 | N1737;
  assign N1739 = preissue_pkt_i[5] | N1738;
  assign N1740 = preissue_pkt_i[4] | N1739;
  assign N1741 = N395 | N1740;
  assign N1742 = N396 | N1741;
  assign N1743 = ~N1742;
  assign N1744 = N1734 | N1743;
  assign N1745 = N393 | N971;
  assign N1746 = preissue_pkt_i[28] | N1745;
  assign N1747 = preissue_pkt_i[27] | N1746;
  assign N1748 = preissue_pkt_i[16] | N1747;
  assign N1749 = preissue_pkt_i[15] | N1748;
  assign N1750 = N2305 | N1749;
  assign N1751 = N1327 | N1750;
  assign N1752 = preissue_pkt_i[7] | N1751;
  assign N1753 = N394 | N1752;
  assign N1754 = preissue_pkt_i[5] | N1753;
  assign N1755 = preissue_pkt_i[4] | N1754;
  assign N1756 = N395 | N1755;
  assign N1757 = N396 | N1756;
  assign N1758 = ~N1757;
  assign N1759 = N1744 | N1758;
  assign N1760 = N2304 | N1787;
  assign N1761 = preissue_pkt_i[14] | N1760;
  assign N1762 = N1327 | N1761;
  assign N1763 = preissue_pkt_i[7] | N1762;
  assign N1764 = N394 | N1763;
  assign N1765 = preissue_pkt_i[5] | N1764;
  assign N1766 = preissue_pkt_i[4] | N1765;
  assign N1767 = N395 | N1766;
  assign N1768 = N396 | N1767;
  assign N1769 = ~N1768;
  assign N1770 = N1759 | N1769;
  assign N1771 = N2305 | N1788;
  assign N1772 = N1327 | N1771;
  assign N1773 = preissue_pkt_i[7] | N1772;
  assign N1774 = N394 | N1773;
  assign N1775 = preissue_pkt_i[5] | N1774;
  assign N1776 = preissue_pkt_i[4] | N1775;
  assign N1777 = N395 | N1776;
  assign N1778 = N396 | N1777;
  assign N1779 = ~N1778;
  assign N1780 = N1770 | N1779;
  assign N1781 = preissue_pkt_i[32] | N2135;
  assign N1782 = N462 | N1781;
  assign N1783 = preissue_pkt_i[30] | N1782;
  assign N1784 = preissue_pkt_i[29] | N1783;
  assign N1785 = preissue_pkt_i[28] | N1784;
  assign N1786 = preissue_pkt_i[27] | N1785;
  assign N1787 = preissue_pkt_i[16] | N1786;
  assign N1788 = preissue_pkt_i[15] | N1787;
  assign N1789 = preissue_pkt_i[14] | N1788;
  assign N1790 = N1327 | N1789;
  assign N1791 = preissue_pkt_i[7] | N1790;
  assign N1792 = N394 | N1791;
  assign N1793 = preissue_pkt_i[5] | N1792;
  assign N1794 = preissue_pkt_i[4] | N1793;
  assign N1795 = N395 | N1794;
  assign N1796 = N396 | N1795;
  assign N1797 = ~N1796;
  assign N1798 = N1780 | N1797;
  assign N1799 = N2305 | N2220;
  assign N1800 = N1327 | N1799;
  assign N1801 = preissue_pkt_i[7] | N1800;
  assign N1802 = N394 | N1801;
  assign N1803 = preissue_pkt_i[5] | N1802;
  assign N1804 = preissue_pkt_i[4] | N1803;
  assign N1805 = N395 | N1804;
  assign N1806 = N396 | N1805;
  assign N1807 = ~N1806;
  assign N1808 = N1798 | N1807;
  assign N1809 = preissue_pkt_i[27] | N525;
  assign N1810 = N1327 | N1809;
  assign N1811 = preissue_pkt_i[7] | N1810;
  assign N1812 = N394 | N1811;
  assign N1813 = preissue_pkt_i[5] | N1812;
  assign N1814 = preissue_pkt_i[4] | N1813;
  assign N1815 = N395 | N1814;
  assign N1816 = N396 | N1815;
  assign N1817 = ~N1816;
  assign N1818 = N1808 | N1817;
  assign N1819 = N1327 | N402;
  assign N1820 = preissue_pkt_i[7] | N1819;
  assign N1821 = N394 | N1820;
  assign N1822 = preissue_pkt_i[5] | N1821;
  assign N1823 = preissue_pkt_i[4] | N1822;
  assign N1824 = N395 | N1823;
  assign N1825 = N396 | N1824;
  assign N1826 = ~N1825;
  assign N1827 = N1818 | N1826;
  assign N1828 = preissue_pkt_i[28] | N2307;
  assign N1829 = preissue_pkt_i[27] | N1828;
  assign N1830 = N1327 | N1829;
  assign N1831 = preissue_pkt_i[7] | N1830;
  assign N1832 = N394 | N1831;
  assign N1833 = preissue_pkt_i[5] | N1832;
  assign N1834 = preissue_pkt_i[4] | N1833;
  assign N1835 = N395 | N1834;
  assign N1836 = N396 | N1835;
  assign N1837 = ~N1836;
  assign N1838 = N1827 | N1837;
  assign N1839 = N393 | N2306;
  assign N1840 = preissue_pkt_i[28] | N1839;
  assign N1841 = preissue_pkt_i[27] | N1840;
  assign N1842 = N1327 | N1841;
  assign N1843 = preissue_pkt_i[7] | N1842;
  assign N1844 = N394 | N1843;
  assign N1845 = preissue_pkt_i[5] | N1844;
  assign N1846 = preissue_pkt_i[4] | N1845;
  assign N1847 = N395 | N1846;
  assign N1848 = N396 | N1847;
  assign N1849 = ~N1848;
  assign N1850 = N1838 | N1849;
  assign N1851 = N2303 | N1289;
  assign N1852 = N393 | N1851;
  assign N1853 = preissue_pkt_i[28] | N1852;
  assign N1854 = preissue_pkt_i[27] | N1853;
  assign N1855 = preissue_pkt_i[26] | N1854;
  assign N1856 = preissue_pkt_i[25] | N1855;
  assign N1857 = preissue_pkt_i[24] | N1856;
  assign N1858 = preissue_pkt_i[23] | N1857;
  assign N1859 = preissue_pkt_i[22] | N1858;
  assign N1860 = N1327 | N1859;
  assign N1861 = preissue_pkt_i[7] | N1860;
  assign N1862 = N394 | N1861;
  assign N1863 = preissue_pkt_i[5] | N1862;
  assign N1864 = preissue_pkt_i[4] | N1863;
  assign N1865 = N395 | N1864;
  assign N1866 = N396 | N1865;
  assign N1867 = ~N1866;
  assign N1868 = N1850 | N1867;
  assign N1869 = N2684 & preissue_pkt_i[8];
  assign N1870 = N1328 & preissue_pkt_i[6];
  assign N1871 = N1869 & N1870;
  assign N1872 = N1871 & N1407;
  assign N1874 = N1007 & N1974;
  assign N1875 = N1874 & N1882;
  assign N1876 = N1875 & N1894;
  assign N1877 = N1874 & N1889;
  assign N1878 = N1877 & N1883;
  assign N1880 = N2685 & N2686;
  assign N1881 = N1183 & N2079;
  assign N1882 = N1975 & N1880;
  assign N1883 = N1881 & N2035;
  assign N1884 = N2446 & N1882;
  assign N1885 = N1884 & N1883;
  assign N1886 = N1183 & preissue_pkt_i[23];
  assign N1887 = N1886 & N2035;
  assign N1888 = N1884 & N1887;
  assign N1889 = N1978 & N1880;
  assign N1890 = N2446 & N1889;
  assign N1891 = N1890 & N1883;
  assign N1892 = N1890 & N1887;
  assign N1894 = N1881 & preissue_pkt_i[22];
  assign N1895 = N1884 & N1894;
  assign N1896 = N1886 & preissue_pkt_i[22];
  assign N1897 = N1884 & N1896;
  assign N1898 = N1890 & N1894;
  assign N1899 = N1890 & N1896;
  assign N1901 = N2445 & N1986;
  assign N1902 = N1901 & N1882;
  assign N1903 = N1902 & N1883;
  assign N1904 = N1902 & N1887;
  assign N1905 = N1901 & N1889;
  assign N1906 = N1905 & N1883;
  assign N1907 = N1905 & N1887;
  assign N1909 = N1902 & N1894;
  assign N1910 = N1902 & N1896;
  assign N1911 = N1905 & N1894;
  assign N1912 = N1905 & N1896;
  assign N1914 = N2035 & N1631;
  assign N1915 = N1881 & N1914;
  assign N1916 = N2451 & N1882;
  assign N1917 = N1915 & N1410;
  assign N1918 = N1916 & N1917;
  assign N1919 = N2451 & N1889;
  assign N1920 = N1919 & N1917;
  assign N1922 = N2445 & N2457;
  assign N1923 = N1922 & N1882;
  assign N1924 = N1923 & N1917;
  assign N1925 = N1922 & N1889;
  assign N1926 = N1925 & N1917;
  assign N1928 = N1973 & N2005;
  assign N1929 = N1975 & N1354;
  assign N1930 = N1928 & N1929;
  assign N1931 = N1930 & N2305;
  assign N1932 = N1978 & N1354;
  assign N1933 = N1928 & N1932;
  assign N1934 = N1933 & N2305;
  assign N1936 = N1930 & preissue_pkt_i[14];
  assign N1937 = N1933 & preissue_pkt_i[14];
  assign N1939 = N1975 & N1363;
  assign N1940 = N1928 & N1939;
  assign N1941 = N1940 & N2305;
  assign N1942 = N1978 & N1363;
  assign N1943 = N1928 & N1942;
  assign N1944 = N1943 & N2305;
  assign N1946 = N616 & N1354;
  assign N1947 = N1928 & N1946;
  assign N1948 = N1947 & N2305;
  assign N1949 = N591 & N1354;
  assign N1950 = N1928 & N1949;
  assign N1951 = N1950 & N2305;
  assign N1953 = N1947 & preissue_pkt_i[14];
  assign N1954 = N1950 & preissue_pkt_i[14];
  assign N1956 = N2440 & N1939;
  assign N1957 = N1956 & N2305;
  assign N1958 = N2440 & N1942;
  assign N1959 = N1958 & N2305;
  assign N1961 = N2440 & N1929;
  assign N1962 = N1961 & preissue_pkt_i[14];
  assign N1963 = N2440 & N1932;
  assign N1964 = N1963 & preissue_pkt_i[14];
  assign N1966 = N1961 & N2305;
  assign N1967 = N1963 & N2305;
  assign N1969 = N1915 & N1411;
  assign N1970 = N1916 & N1969;
  assign N1971 = N1919 & N1969;
  assign N1973 = N2135 & N1287;
  assign N1974 = N462 & N2303;
  assign N1975 = N393 & N523;
  assign N1976 = N1973 & N1974;
  assign N1977 = N1976 & N1975;
  assign N1978 = N393 & preissue_pkt_i[27];
  assign N1979 = N1976 & N1978;
  assign N1981 = N1976 & N616;
  assign N1982 = N2135 & N1287;
  assign N1983 = N1982 & N1974;
  assign N1984 = N1983 & N591;
  assign N1986 = N462 & preissue_pkt_i[30];
  assign N1987 = N1982 & N1986;
  assign N1988 = N1987 & N1975;
  assign N1989 = N1987 & N1978;
  assign N1991 = N1987 & N616;
  assign N1992 = N1987 & N591;
  assign N1994 = N2002 & N1986;
  assign N1995 = N616 & N1880;
  assign N1996 = N1994 & N1995;
  assign N1997 = N1996 & N1883;
  assign N1998 = N591 & N1880;
  assign N1999 = N1994 & N1998;
  assign N2000 = N1999 & N1883;
  assign N2002 = N2135 & preissue_pkt_i[32];
  assign N2003 = preissue_pkt_i[27] & preissue_pkt_i[22];
  assign N2004 = N2002 & N2003;
  assign N2005 = preissue_pkt_i[31] & N2303;
  assign N2006 = N2002 & N2005;
  assign N2007 = N2006 & preissue_pkt_i[27];
  assign N2008 = preissue_pkt_i[32] & preissue_pkt_i[26];
  assign N2009 = preissue_pkt_i[32] & preissue_pkt_i[25];
  assign N2010 = preissue_pkt_i[32] & preissue_pkt_i[24];
  assign N2011 = preissue_pkt_i[30] & preissue_pkt_i[22];
  assign N2012 = N2002 & N2011;
  assign N2013 = N2460 & preissue_pkt_i[22];
  assign N2014 = N2460 & preissue_pkt_i[23];
  assign N2015 = N622 & preissue_pkt_i[29];
  assign N2016 = N2002 & N2463;
  assign N2017 = N2457 & preissue_pkt_i[14];
  assign N2018 = preissue_pkt_i[32] & N2303;
  assign N2019 = N2018 & preissue_pkt_i[29];
  assign N2020 = N622 & preissue_pkt_i[22];
  assign N2021 = N2002 & preissue_pkt_i[23];
  assign N2022 = N2303 & N523;
  assign N2023 = N2002 & N2022;
  assign N2024 = N2023 & N2035;
  assign N2025 = N622 & preissue_pkt_i[23];
  assign N2026 = N2458 & preissue_pkt_i[15];
  assign N2027 = preissue_pkt_i[33] & N1287;
  assign N2028 = N2027 & N462;
  assign N2029 = N2027 & preissue_pkt_i[30];
  assign N2030 = N2027 & preissue_pkt_i[16];
  assign N2031 = N2027 & N1413;
  assign N2032 = N659 & preissue_pkt_i[30];
  assign N2033 = preissue_pkt_i[31] & preissue_pkt_i[16];
  assign N2035 = ~preissue_pkt_i[22];
  assign N2036 = preissue_pkt_i[27] | N1292;
  assign N2037 = preissue_pkt_i[26] | N2036;
  assign N2038 = preissue_pkt_i[25] | N2037;
  assign N2039 = preissue_pkt_i[24] | N2038;
  assign N2040 = preissue_pkt_i[23] | N2039;
  assign N2041 = N2035 | N2040;
  assign N2042 = N1327 | N2041;
  assign N2043 = preissue_pkt_i[7] | N2042;
  assign N2044 = N394 | N2043;
  assign N2045 = preissue_pkt_i[5] | N2044;
  assign N2046 = preissue_pkt_i[4] | N2045;
  assign N2047 = N395 | N2046;
  assign N2048 = N396 | N2047;
  assign N2049 = N523 | N1292;
  assign N2050 = preissue_pkt_i[26] | N2049;
  assign N2051 = preissue_pkt_i[25] | N2050;
  assign N2052 = preissue_pkt_i[24] | N2051;
  assign N2053 = preissue_pkt_i[23] | N2052;
  assign N2054 = preissue_pkt_i[22] | N2053;
  assign N2055 = N1327 | N2054;
  assign N2056 = preissue_pkt_i[7] | N2055;
  assign N2057 = N394 | N2056;
  assign N2058 = preissue_pkt_i[5] | N2057;
  assign N2059 = preissue_pkt_i[4] | N2058;
  assign N2060 = N395 | N2059;
  assign N2061 = N396 | N2060;
  assign N2062 = preissue_pkt_i[30] | N2137;
  assign N2063 = preissue_pkt_i[29] | N2062;
  assign N2064 = preissue_pkt_i[28] | N2063;
  assign N2065 = preissue_pkt_i[27] | N2064;
  assign N2066 = preissue_pkt_i[26] | N2065;
  assign N2067 = preissue_pkt_i[25] | N2066;
  assign N2068 = preissue_pkt_i[24] | N2067;
  assign N2069 = preissue_pkt_i[23] | N2068;
  assign N2070 = preissue_pkt_i[22] | N2069;
  assign N2071 = N1327 | N2070;
  assign N2072 = preissue_pkt_i[7] | N2071;
  assign N2073 = N394 | N2072;
  assign N2074 = preissue_pkt_i[5] | N2073;
  assign N2075 = preissue_pkt_i[4] | N2074;
  assign N2076 = N395 | N2075;
  assign N2077 = N396 | N2076;
  assign N2078 = ~N2077;
  assign N2079 = ~preissue_pkt_i[23];
  assign N2080 = N2079 | N2068;
  assign N2081 = preissue_pkt_i[22] | N2080;
  assign N2082 = N1327 | N2081;
  assign N2083 = preissue_pkt_i[7] | N2082;
  assign N2084 = N394 | N2083;
  assign N2085 = preissue_pkt_i[5] | N2084;
  assign N2086 = preissue_pkt_i[4] | N2085;
  assign N2087 = N395 | N2086;
  assign N2088 = N396 | N2087;
  assign N2089 = ~N2088;
  assign N2090 = N2078 | N2089;
  assign N2091 = N523 | N2064;
  assign N2092 = preissue_pkt_i[26] | N2091;
  assign N2093 = preissue_pkt_i[25] | N2092;
  assign N2094 = preissue_pkt_i[24] | N2093;
  assign N2095 = preissue_pkt_i[23] | N2094;
  assign N2096 = preissue_pkt_i[22] | N2095;
  assign N2097 = N1327 | N2096;
  assign N2098 = preissue_pkt_i[7] | N2097;
  assign N2099 = N394 | N2098;
  assign N2100 = preissue_pkt_i[5] | N2099;
  assign N2101 = preissue_pkt_i[4] | N2100;
  assign N2102 = N395 | N2101;
  assign N2103 = N396 | N2102;
  assign N2104 = ~N2103;
  assign N2105 = N2078 | N2104;
  assign N2106 = N2035 | N2069;
  assign N2107 = N1327 | N2106;
  assign N2108 = preissue_pkt_i[7] | N2107;
  assign N2109 = N394 | N2108;
  assign N2110 = preissue_pkt_i[5] | N2109;
  assign N2111 = preissue_pkt_i[4] | N2110;
  assign N2112 = N395 | N2111;
  assign N2113 = N396 | N2112;
  assign N2114 = ~N2113;
  assign N2115 = N2035 | N2080;
  assign N2116 = N1327 | N2115;
  assign N2117 = preissue_pkt_i[7] | N2116;
  assign N2118 = N394 | N2117;
  assign N2119 = preissue_pkt_i[5] | N2118;
  assign N2120 = preissue_pkt_i[4] | N2119;
  assign N2121 = N395 | N2120;
  assign N2122 = N396 | N2121;
  assign N2123 = ~N2122;
  assign N2124 = N2114 | N2123;
  assign N2125 = N2035 | N2095;
  assign N2126 = N1327 | N2125;
  assign N2127 = preissue_pkt_i[7] | N2126;
  assign N2128 = N394 | N2127;
  assign N2129 = preissue_pkt_i[5] | N2128;
  assign N2130 = preissue_pkt_i[4] | N2129;
  assign N2131 = N395 | N2130;
  assign N2132 = N396 | N2131;
  assign N2133 = ~N2132;
  assign N2134 = N2114 | N2133;
  assign N2135 = ~preissue_pkt_i[33];
  assign N2136 = N1287 | N2135;
  assign N2137 = preissue_pkt_i[31] | N2136;
  assign N2138 = N2303 | N2137;
  assign N2139 = preissue_pkt_i[29] | N2138;
  assign N2140 = preissue_pkt_i[28] | N2139;
  assign N2141 = preissue_pkt_i[27] | N2140;
  assign N2142 = preissue_pkt_i[26] | N2141;
  assign N2143 = preissue_pkt_i[25] | N2142;
  assign N2144 = preissue_pkt_i[24] | N2143;
  assign N2145 = preissue_pkt_i[23] | N2144;
  assign N2146 = preissue_pkt_i[22] | N2145;
  assign N2147 = N1327 | N2146;
  assign N2148 = preissue_pkt_i[7] | N2147;
  assign N2149 = N394 | N2148;
  assign N2150 = preissue_pkt_i[5] | N2149;
  assign N2151 = preissue_pkt_i[4] | N2150;
  assign N2152 = N395 | N2151;
  assign N2153 = N396 | N2152;
  assign N2154 = ~N2153;
  assign N2155 = N523 | N2140;
  assign N2156 = preissue_pkt_i[26] | N2155;
  assign N2157 = preissue_pkt_i[25] | N2156;
  assign N2158 = preissue_pkt_i[24] | N2157;
  assign N2159 = preissue_pkt_i[23] | N2158;
  assign N2160 = preissue_pkt_i[22] | N2159;
  assign N2161 = N1327 | N2160;
  assign N2162 = preissue_pkt_i[7] | N2161;
  assign N2163 = N394 | N2162;
  assign N2164 = preissue_pkt_i[5] | N2163;
  assign N2165 = preissue_pkt_i[4] | N2164;
  assign N2166 = N395 | N2165;
  assign N2167 = N396 | N2166;
  assign N2168 = ~N2167;
  assign N2169 = N2154 | N2168;
  assign N2170 = N2079 | N2144;
  assign N2171 = preissue_pkt_i[22] | N2170;
  assign N2172 = N1327 | N2171;
  assign N2173 = preissue_pkt_i[7] | N2172;
  assign N2174 = N394 | N2173;
  assign N2175 = preissue_pkt_i[5] | N2174;
  assign N2176 = preissue_pkt_i[4] | N2175;
  assign N2177 = N395 | N2176;
  assign N2178 = N396 | N2177;
  assign N2179 = ~N2178;
  assign N2180 = N2154 | N2179;
  assign N2181 = N2035 | N2145;
  assign N2182 = N1327 | N2181;
  assign N2183 = preissue_pkt_i[7] | N2182;
  assign N2184 = N394 | N2183;
  assign N2185 = preissue_pkt_i[5] | N2184;
  assign N2186 = preissue_pkt_i[4] | N2185;
  assign N2187 = N395 | N2186;
  assign N2188 = N396 | N2187;
  assign N2189 = ~N2188;
  assign N2190 = N2035 | N2159;
  assign N2191 = N1327 | N2190;
  assign N2192 = preissue_pkt_i[7] | N2191;
  assign N2193 = N394 | N2192;
  assign N2194 = preissue_pkt_i[5] | N2193;
  assign N2195 = preissue_pkt_i[4] | N2194;
  assign N2196 = N395 | N2195;
  assign N2197 = N396 | N2196;
  assign N2198 = ~N2197;
  assign N2199 = N2189 | N2198;
  assign N2200 = N2035 | N2170;
  assign N2201 = N1327 | N2200;
  assign N2202 = preissue_pkt_i[7] | N2201;
  assign N2203 = N394 | N2202;
  assign N2204 = preissue_pkt_i[5] | N2203;
  assign N2205 = preissue_pkt_i[4] | N2204;
  assign N2206 = N395 | N2205;
  assign N2207 = N396 | N2206;
  assign N2208 = ~N2207;
  assign N2209 = N2189 | N2208;
  assign N2210 = preissue_pkt_i[30] | N2230;
  assign N2211 = preissue_pkt_i[29] | N2210;
  assign N2212 = preissue_pkt_i[28] | N2211;
  assign N2213 = preissue_pkt_i[27] | N2212;
  assign N2214 = preissue_pkt_i[26] | N2213;
  assign N2215 = preissue_pkt_i[25] | N2214;
  assign N2216 = preissue_pkt_i[24] | N2215;
  assign N2217 = preissue_pkt_i[23] | N2216;
  assign N2218 = preissue_pkt_i[22] | N2217;
  assign N2219 = preissue_pkt_i[16] | N2218;
  assign N2220 = preissue_pkt_i[15] | N2219;
  assign N2221 = preissue_pkt_i[14] | N2220;
  assign N2222 = N1327 | N2221;
  assign N2223 = preissue_pkt_i[7] | N2222;
  assign N2224 = N394 | N2223;
  assign N2225 = preissue_pkt_i[5] | N2224;
  assign N2226 = preissue_pkt_i[4] | N2225;
  assign N2227 = N395 | N2226;
  assign N2228 = N396 | N2227;
  assign N2229 = ~N2228;
  assign N2230 = N462 | N2136;
  assign N2231 = N2303 | N2230;
  assign N2232 = preissue_pkt_i[29] | N2231;
  assign N2233 = preissue_pkt_i[28] | N2232;
  assign N2234 = preissue_pkt_i[27] | N2233;
  assign N2235 = preissue_pkt_i[26] | N2234;
  assign N2236 = preissue_pkt_i[25] | N2235;
  assign N2237 = preissue_pkt_i[24] | N2236;
  assign N2238 = preissue_pkt_i[23] | N2237;
  assign N2239 = preissue_pkt_i[22] | N2238;
  assign N2240 = preissue_pkt_i[16] | N2239;
  assign N2241 = preissue_pkt_i[15] | N2240;
  assign N2242 = preissue_pkt_i[14] | N2241;
  assign N2243 = N1327 | N2242;
  assign N2244 = preissue_pkt_i[7] | N2243;
  assign N2245 = N394 | N2244;
  assign N2246 = preissue_pkt_i[5] | N2245;
  assign N2247 = preissue_pkt_i[4] | N2246;
  assign N2248 = N395 | N2247;
  assign N2249 = N396 | N2248;
  assign N2250 = ~N2249;
  assign N2286 = N394 & preissue_pkt_i[3];
  assign N2287 = N2577 & N2286;
  assign N2288 = N2287 & preissue_pkt_i[2];
  assign N2290 = N1329 & N1330;
  assign N2291 = preissue_pkt_i[5] | N1330;
  assign N2293 = N1329 | preissue_pkt_i[4];
  assign N2295 = preissue_pkt_i[5] & preissue_pkt_i[4];
  assign N2303 = ~preissue_pkt_i[30];
  assign N2304 = ~preissue_pkt_i[15];
  assign N2305 = ~preissue_pkt_i[14];
  assign N2306 = N2303 | N398;
  assign N2307 = preissue_pkt_i[29] | N2306;
  assign N2308 = preissue_pkt_i[26] | N2307;
  assign N2309 = preissue_pkt_i[25] | N2308;
  assign N2310 = preissue_pkt_i[24] | N2309;
  assign N2311 = preissue_pkt_i[23] | N2310;
  assign N2312 = preissue_pkt_i[22] | N2311;
  assign N2313 = preissue_pkt_i[16] | N2312;
  assign N2314 = N2304 | N2313;
  assign N2315 = N2305 | N2314;
  assign N2316 = preissue_pkt_i[8] | N2315;
  assign N2317 = N1328 | N2316;
  assign N2318 = preissue_pkt_i[6] | N2317;
  assign N2319 = N1329 | N2318;
  assign N2320 = N1330 | N2319;
  assign N2321 = N395 | N2320;
  assign N2322 = N396 | N2321;
  assign N2323 = ~N2322;
  assign N2324 = preissue_pkt_i[14] | N2314;
  assign N2325 = preissue_pkt_i[8] | N2324;
  assign N2326 = N1328 | N2325;
  assign N2327 = preissue_pkt_i[6] | N2326;
  assign N2328 = N1329 | N2327;
  assign N2329 = N1330 | N2328;
  assign N2330 = N395 | N2329;
  assign N2331 = N396 | N2330;
  assign N2332 = ~N2331;
  assign N2333 = N2323 | N2332;
  assign N2335 = N2575 & N1396;
  assign N2336 = N1420 & N2335;
  assign N2337 = N2336 & preissue_pkt_i[2];
  assign N2339 = N2079 & N2035;
  assign N2340 = N2339 & preissue_pkt_i[14];
  assign N2341 = N2389 & N2340;
  assign N2342 = N2339 & N2305;
  assign N2343 = N2389 & N2342;
  assign N2344 = N1987 & N668;
  assign N2345 = preissue_pkt_i[29] & N2305;
  assign N2346 = N1987 & N2345;
  assign N2347 = N1983 & N668;
  assign N2348 = N1983 & N2345;
  assign N2349 = N393 & preissue_pkt_i[14];
  assign N2350 = N1983 & N2349;
  assign N2351 = N393 & N2305;
  assign N2352 = N1983 & N2351;
  assign N2353 = N2425 & N2349;
  assign N2354 = N2425 & N2351;
  assign N2355 = N2006 & N2349;
  assign N2356 = N2006 & N2351;
  assign N2357 = N2420 & N2349;
  assign N2358 = N2420 & N2351;
  assign N2359 = N2435 & N2349;
  assign N2360 = N2435 & N2351;
  assign N2361 = N2440 & N2349;
  assign N2362 = N2440 & N2351;
  assign N2363 = N2446 & N2349;
  assign N2364 = N2446 & N2351;
  assign N2365 = N2451 & N2349;
  assign N2366 = N2451 & N2351;
  assign N2382 = N393 & N2685;
  assign N2383 = N2686 & N1183;
  assign N2384 = preissue_pkt_i[14] & N1327;
  assign N2385 = N2382 & N2383;
  assign N2386 = N2339 & N1363;
  assign N2387 = N2384 & N1405;
  assign N2388 = N2295 & N173;
  assign N2389 = N1987 & N2385;
  assign N2390 = N2386 & N2387;
  assign N2391 = N2389 & N2390;
  assign N2392 = N2391 & N2388;
  assign N2393 = N2305 & N1327;
  assign N2394 = N2393 & N1405;
  assign N2395 = N2386 & N2394;
  assign N2396 = N2389 & N2395;
  assign N2397 = N2396 & N2388;
  assign N2398 = N688 & N1413;
  assign N2399 = N1419 & N2575;
  assign N2400 = N1396 & preissue_pkt_i[2];
  assign N2401 = N1987 & N2398;
  assign N2402 = N2399 & N2400;
  assign N2403 = N2401 & N2402;
  assign N2404 = N688 & N1412;
  assign N2405 = N1987 & N2404;
  assign N2406 = N2405 & N2402;
  assign N2408 = N1983 & N2398;
  assign N2409 = N2408 & N2402;
  assign N2410 = N1983 & N2404;
  assign N2411 = N2410 & N2402;
  assign N2413 = N393 & N1631;
  assign N2414 = N2413 & N1413;
  assign N2415 = N2006 & N2414;
  assign N2416 = N2415 & N2402;
  assign N2417 = N2413 & N1412;
  assign N2418 = N2006 & N2417;
  assign N2419 = N2418 & N2402;
  assign N2420 = N2002 & N1974;
  assign N2421 = N2420 & N2414;
  assign N2422 = N2421 & N2402;
  assign N2423 = N2420 & N2417;
  assign N2424 = N2423 & N2402;
  assign N2425 = N1982 & N2005;
  assign N2426 = N2425 & N2414;
  assign N2427 = N2426 & N2402;
  assign N2428 = N2425 & N2417;
  assign N2429 = N2428 & N2402;
  assign N2431 = N1983 & N2414;
  assign N2432 = N2431 & N2402;
  assign N2433 = N1983 & N2417;
  assign N2434 = N2433 & N2402;
  assign N2435 = N2027 & N1974;
  assign N2436 = N2435 & N2414;
  assign N2437 = N2436 & N2402;
  assign N2438 = N2435 & N2417;
  assign N2439 = N2438 & N2402;
  assign N2440 = N2027 & N2005;
  assign N2441 = N2440 & N2414;
  assign N2442 = N2441 & N2402;
  assign N2443 = N2440 & N2417;
  assign N2444 = N2443 & N2402;
  assign N2445 = preissue_pkt_i[33] & preissue_pkt_i[32];
  assign N2446 = N2445 & N1974;
  assign N2447 = N2446 & N2414;
  assign N2448 = N2447 & N2402;
  assign N2449 = N2446 & N2417;
  assign N2450 = N2449 & N2402;
  assign N2451 = N2445 & N2005;
  assign N2452 = N2451 & N2414;
  assign N2453 = N2452 & N2402;
  assign N2454 = N2451 & N2417;
  assign N2455 = N2454 & N2402;
  assign N2457 = preissue_pkt_i[31] & preissue_pkt_i[30];
  assign N2458 = preissue_pkt_i[31] & preissue_pkt_i[29];
  assign N2459 = preissue_pkt_i[33] & preissue_pkt_i[29];
  assign N2460 = preissue_pkt_i[32] & preissue_pkt_i[29];
  assign N2461 = preissue_pkt_i[32] & preissue_pkt_i[30];
  assign N2462 = preissue_pkt_i[33] & preissue_pkt_i[30];
  assign N2463 = preissue_pkt_i[30] & N393;
  assign N2464 = N2463 & preissue_pkt_i[26];
  assign N2465 = N2463 & preissue_pkt_i[25];
  assign N2466 = N2463 & preissue_pkt_i[24];
  assign N2467 = N2463 & preissue_pkt_i[23];
  assign N2468 = N2463 & preissue_pkt_i[22];
  assign N2541 = preissue_pkt_i[8] | N1328;
  assign N2542 = N394 | preissue_pkt_i[5];
  assign N2543 = N2541 | N2542;
  assign N2544 = N2543 | N1330;
  assign N2545 = N179 | N2542;
  assign N2546 = N2545 | N1330;
  assign N2548 = N1327 | N1328;
  assign N2549 = preissue_pkt_i[6] | N1329;
  assign N2550 = N2548 | N2549;
  assign N2551 = N2550 | N1330;
  assign N2553 = N2548 | N212;
  assign N2554 = N2553 | preissue_pkt_i[4];
  assign N2556 = N2541 | N212;
  assign N2557 = N2556 | preissue_pkt_i[4];
  assign N2558 = N2556 | N1330;
  assign N2560 = N2553 | N1330;
  assign N2561 = N394 & N1329;
  assign N2562 = N1426 & N2561;
  assign N2563 = N2562 & N1330;
  assign N2564 = N2545 | preissue_pkt_i[4];
  assign N2565 = N394 | N1329;
  assign N2566 = N179 | N2565;
  assign N2567 = N2566 | preissue_pkt_i[4];
  assign N2568 = N179 | N212;
  assign N2569 = N2568 | N1330;
  assign N2571 = N1327 & preissue_pkt_i[5];
  assign N2572 = N2571 & preissue_pkt_i[4];
  assign N2573 = preissue_pkt_i[7] & preissue_pkt_i[6];
  assign N2574 = N2573 & N1330;
  assign N2575 = N394 & preissue_pkt_i[5];
  assign N2576 = N2575 & N1330;
  assign N2577 = preissue_pkt_i[8] & N1328;
  assign N2643 = N1363 & N2393;
  assign N2644 = N2643 & N1017;
  assign N2645 = N2644 & N173;
  assign N2646 = N1363 & N2384;
  assign N2647 = N2646 & N1017;
  assign N2648 = N2647 & N173;
  assign N2650 = N523 & N1631;
  assign N2651 = N2666 & N2650;
  assign N2652 = N2425 & N2651;
  assign N2653 = N2652 & N2672;
  assign N2654 = N2653 & preissue_pkt_i[2];
  assign N2655 = N2652 & N2676;
  assign N2656 = N2655 & preissue_pkt_i[2];
  assign N2658 = N1410 & N1419;
  assign N2659 = N2658 & N2670;
  assign N2660 = N2671 & N2659;
  assign N2661 = N2660 & preissue_pkt_i[2];
  assign N2662 = N2658 & N2675;
  assign N2663 = N2671 & N2662;
  assign N2664 = N2663 & preissue_pkt_i[2];
  assign N2666 = N393 & N2684;
  assign N2667 = preissue_pkt_i[6] & N1329;
  assign N2668 = N2666 & N654;
  assign N2669 = N1412 & N1419;
  assign N2670 = N2667 & N541;
  assign N2671 = N2425 & N2668;
  assign N2672 = N2669 & N2670;
  assign N2673 = N2671 & N2672;
  assign N2674 = N2673 & preissue_pkt_i[2];
  assign N2675 = N239 & N541;
  assign N2676 = N2669 & N2675;
  assign N2677 = N2671 & N2676;
  assign N2678 = N2677 & preissue_pkt_i[2];
  assign N2704 = preissue_pkt_i[12] | preissue_pkt_i[13];
  assign N2705 = preissue_pkt_i[11] | N2704;
  assign N2706 = preissue_pkt_i[10] | N2705;
  assign N2707 = preissue_pkt_i[9] | N2706;
  assign N2708 = preissue_pkt_i[27] | preissue_pkt_i[28];
  assign N2709 = ~N2708;
  assign N2710 = N1328 | preissue_pkt_i[8];
  assign N2711 = N394 | N2710;
  assign N2712 = N1329 | N2711;
  assign N2713 = preissue_pkt_i[4] | N2712;
  assign N2714 = N395 | N2713;
  assign N2715 = N396 | N2714;
  assign N2716 = ~N2715;
  assign N2717 = preissue_pkt_i[7] | preissue_pkt_i[8];
  assign N2718 = N394 | N2717;
  assign N2719 = N1329 | N2718;
  assign N2720 = preissue_pkt_i[4] | N2719;
  assign N2721 = N395 | N2720;
  assign N2722 = N396 | N2721;
  assign N2723 = ~N2722;
  assign N2724 = preissue_pkt_i[20] | preissue_pkt_i[21];
  assign N2725 = preissue_pkt_i[19] | N2724;
  assign N2726 = preissue_pkt_i[18] | N2725;
  assign N2727 = preissue_pkt_i[17] | N2726;
  assign N349 = ~N348;
  assign N391 = ~N390;
  assign N392 = (N0)? N391 : 
                (N1)? 1'b0 : 1'b0;
  assign N0 = N2716;
  assign N1 = N2715;
  assign N414 = (N2)? 1'b0 : 
                (N3)? N2716 : 1'b0;
  assign N2 = N413;
  assign N3 = N412;
  assign { N714, N713, N712, N711, N710 } = (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                            (N5)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                            (N6)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                            (N7)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                                            (N8)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                            (N9)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                                            (N10)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                                            (N11)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                            (N12)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                            (N13)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                            (N14)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                            (N15)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                            (N16)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                            (N17)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                            (N18)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                            (N19)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                            (N20)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                            (N21)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                            (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                            (N23)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                            (N24)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                            (N25)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                            (N26)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N4 = N580;
  assign N5 = N587;
  assign N6 = N590;
  assign N7 = N594;
  assign N8 = N596;
  assign N9 = N598;
  assign N10 = N600;
  assign N11 = N603;
  assign N12 = N611;
  assign N13 = N614;
  assign N14 = N620;
  assign N15 = N621;
  assign N16 = N624;
  assign N17 = N627;
  assign N18 = N630;
  assign N19 = N634;
  assign N20 = N635;
  assign N21 = N636;
  assign N22 = N639;
  assign N23 = N642;
  assign N24 = N645;
  assign N25 = N649;
  assign N26 = N709;
  assign N715 = (N4)? 1'b0 : 
                (N5)? 1'b0 : 
                (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N8)? 1'b0 : 
                (N9)? 1'b0 : 
                (N10)? 1'b0 : 
                (N11)? 1'b0 : 
                (N12)? 1'b0 : 
                (N13)? 1'b0 : 
                (N14)? 1'b0 : 
                (N15)? 1'b0 : 
                (N16)? 1'b0 : 
                (N17)? 1'b0 : 
                (N18)? 1'b0 : 
                (N19)? 1'b0 : 
                (N20)? 1'b0 : 
                (N21)? 1'b0 : 
                (N22)? 1'b0 : 
                (N23)? 1'b0 : 
                (N24)? 1'b0 : 
                (N25)? 1'b0 : 
                (N26)? 1'b1 : 1'b0;
  assign { N720, N719, N718, N717, N716 } = (N27)? { N714, N713, N712, N711, N710 } : 
                                            (N546)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N27 = N545;
  assign N721 = (N27)? N715 : 
                (N546)? 1'b1 : 1'b0;
  assign N835 = (N28)? 1'b1 : 
                (N834)? N803 : 1'b0;
  assign N28 = N833;
  assign { N855, N854 } = (N29)? { 1'b1, 1'b0 } : 
                          (N853)? { N835, N835 } : 1'b0;
  assign N29 = N852;
  assign { N895, N894, N893, N892 } = (N30)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                      (N891)? { N852, N852, N855, N854 } : 1'b0;
  assign N30 = N890;
  assign { N913, N912, N911, N910, N909 } = (N31)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                            (N908)? { N895, N894, N890, N893, N892 } : 1'b0;
  assign N31 = N907;
  assign { N932, N931, N930, N929, N928 } = (N32)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                            (N927)? { N913, N912, N911, N910, N909 } : 1'b0;
  assign N32 = N926;
  assign { N938, N937, N936 } = (N33)? { 1'b0, 1'b1, 1'b0 } : 
                                (N34)? { N930, N929, N928 } : 1'b0;
  assign N33 = N935;
  assign N34 = N934;
  assign { N990, N989, N988 } = (N35)? { 1'b0, 1'b1, 1'b1 } : 
                                (N987)? { N926, N932, N931 } : 1'b0;
  assign N35 = N986;
  assign N1002 = (N36)? N1000 : 
                 (N37)? 1'b0 : 1'b0;
  assign N36 = N2723;
  assign N37 = N2722;
  assign { N1026, N1025 } = (N38)? { 1'b1, 1'b1 } : 
                            (N39)? { 1'b1, 1'b0 } : 
                            (N1024)? { 1'b0, N2723 } : 1'b0;
  assign N38 = N1006;
  assign N39 = N1022;
  assign { N1124, N1123, N1122, N1121, N1120 } = (N40)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                 (N41)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                                 (N42)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                 (N43)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                                 (N44)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                                 (N45)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                 (N46)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                                 (N47)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                                                 (N48)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                                 (N49)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                 (N50)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                 (N51)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                                 (N52)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                                 (N53)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                                 (N1119)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N40 = N1052;
  assign N41 = N1053;
  assign N42 = N1054;
  assign N43 = N593;
  assign N44 = N1062;
  assign N45 = N599;
  assign N46 = N1067;
  assign N47 = N1080;
  assign N48 = N1086;
  assign N49 = N1093;
  assign N50 = N1095;
  assign N51 = N1098;
  assign N52 = N1101;
  assign N53 = N1105;
  assign N1125 = (N40)? 1'b0 : 
                 (N41)? 1'b0 : 
                 (N42)? 1'b0 : 
                 (N43)? 1'b0 : 
                 (N44)? 1'b0 : 
                 (N45)? 1'b0 : 
                 (N46)? 1'b0 : 
                 (N47)? 1'b0 : 
                 (N48)? 1'b0 : 
                 (N49)? 1'b0 : 
                 (N50)? 1'b0 : 
                 (N51)? 1'b0 : 
                 (N52)? 1'b0 : 
                 (N53)? 1'b0 : 
                 (N1119)? 1'b1 : 1'b0;
  assign { N1130, N1129, N1128, N1127, N1126 } = (N54)? { N1124, N1123, N1122, N1121, N1120 } : 
                                                 (N1030)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N54 = N1029;
  assign N1131 = (N54)? N1125 : 
                 (N1030)? 1'b1 : 1'b0;
  assign N1212 = (N55)? 1'b1 : 
                 (N1211)? N1182 : 1'b0;
  assign N55 = N1210;
  assign { N1234, N1233, N1232 } = (N56)? { 1'b0, 1'b1, 1'b1 } : 
                                   (N1231)? { N1153, N1153, N1212 } : 1'b0;
  assign N56 = N1230;
  assign { N1263, N1262, N1261, N1260, N1259 } = (N57)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                                 (N1258)? { N1182, N1234, N1230, N1233, N1232 } : 1'b0;
  assign N57 = N1257;
  assign { N1310, N1309, N1308, N1307, N1306 } = (N58)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                                                 (N1305)? { N1262, N1261, N1260, N1257, N1259 } : 1'b0;
  assign N58 = N1304;
  assign { N1367, N1366, N1365, N1364 } = (N59)? { 1'b1, 1'b1, 1'b0, 1'b0 } : 
                                          (N60)? { 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                          (N61)? { 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                          (N62)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                                          (N63)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                          (N64)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                          (N65)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N59 = N1355;
  assign N60 = N1356;
  assign N61 = N1358;
  assign N62 = N1359;
  assign N63 = N1361;
  assign N64 = N1362;
  assign N65 = N1363;
  assign N1368 = (N59)? 1'b0 : 
                 (N60)? 1'b0 : 
                 (N61)? 1'b0 : 
                 (N62)? 1'b0 : 
                 (N63)? 1'b0 : 
                 (N64)? 1'b0 : 
                 (N65)? 1'b1 : 1'b0;
  assign { N1372, N1371, N1370, N1369 } = (N66)? { N1367, N1366, N1365, N1364 } : 
                                          (N67)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N66 = N1353;
  assign N67 = N1352;
  assign N1373 = (N66)? N1368 : 
                 (N67)? 1'b1 : 1'b0;
  assign { N1380, N1379, N1378 } = (N59)? { 1'b0, 1'b0, 1'b0 } : 
                                   (N60)? { 1'b0, 1'b0, 1'b1 } : 
                                   (N68)? { 1'b0, 1'b1, 1'b0 } : 
                                   (N61)? { 1'b1, 1'b0, 1'b0 } : 
                                   (N62)? { 1'b1, 1'b0, 1'b1 } : 
                                   (N63)? { 1'b1, 1'b1, 1'b0 } : 
                                   (N69)? { 1'b0, 1'b1, 1'b1 } : 
                                   (N64)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N68 = N1376;
  assign N69 = N1377;
  assign N1381 = (N59)? 1'b0 : 
                 (N60)? 1'b0 : 
                 (N68)? 1'b0 : 
                 (N61)? 1'b0 : 
                 (N62)? 1'b0 : 
                 (N63)? 1'b0 : 
                 (N69)? 1'b0 : 
                 (N64)? 1'b1 : 1'b0;
  assign { N1384, N1383, N1382 } = (N70)? { N1380, N1379, N1378 } : 
                                   (N71)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N70 = N1375;
  assign N71 = N1374;
  assign N1385 = (N70)? N1381 : 
                 (N71)? 1'b1 : 1'b0;
  assign N1402 = (N72)? preissue_pkt_i[14] : 
                 (N1401)? 1'b0 : 1'b0;
  assign N72 = N1400;
  assign N1403 = (N72)? N2302 : 
                 (N1401)? 1'b1 : 1'b0;
  assign { N1415, N1414 } = (N73)? { 1'b0, 1'b0 } : 
                            (N74)? { 1'b0, 1'b1 } : 
                            (N75)? { 1'b1, 1'b0 } : 
                            (N76)? { 1'b1, 1'b1 } : 1'b0;
  assign N73 = N1410;
  assign N74 = N1411;
  assign N75 = N1412;
  assign N76 = N1413;
  assign { N1417, N1416 } = (N77)? { N1415, N1414 } : 
                            (N1409)? { 1'b0, 1'b0 } : 1'b0;
  assign N77 = N1408;
  assign N1418 = ~N1408;
  assign N1424 = (N78)? preissue_pkt_i[14] : 
                 (N1423)? 1'b0 : 1'b0;
  assign N78 = N1422;
  assign N1425 = (N78)? N2302 : 
                 (N1423)? 1'b1 : 1'b0;
  assign { N1503, N1502, N1501, N1500, N1499, N1498, N1497 } = (N79)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N80)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                                               (N81)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                                                               (N82)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                                               (N83)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                               (N84)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N85)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                                               (N86)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                                               (N87)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                                               (N88)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N89)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N90)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N91)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N79 = N1431;
  assign N80 = N1434;
  assign N81 = N1437;
  assign N82 = N1440;
  assign N83 = N1445;
  assign N84 = N1448;
  assign N85 = N1452;
  assign N86 = N1455;
  assign N87 = N1469;
  assign N88 = N1473;
  assign N89 = N1476;
  assign N90 = N1485;
  assign N91 = N1505;
  assign N1504 = (N79)? 1'b0 : 
                 (N80)? 1'b1 : 
                 (N81)? 1'b0 : 
                 (N82)? 1'b0 : 
                 (N83)? 1'b0 : 
                 (N84)? 1'b0 : 
                 (N85)? 1'b0 : 
                 (N86)? 1'b0 : 
                 (N87)? 1'b0 : 
                 (N88)? 1'b0 : 
                 (N89)? 1'b0 : 
                 (N90)? 1'b0 : 
                 (N91)? 1'b0 : 1'b0;
  assign N1505 = ~N1496;
  assign N1506 = (N92)? N1504 : 
                 (N1428)? 1'b0 : 1'b0;
  assign N92 = N1427;
  assign N1507 = (N92)? N1505 : 
                 (N1428)? 1'b1 : 1'b0;
  assign { N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508 } = (N92)? { N1503, N1448, N1502, N1501, N1500, N1499, N1498, N1497 } : 
                                                                      (N1428)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1675 = (N93)? N2302 : 
                 (N2688)? N1663 : 
                 (N2690)? N1664 : 
                 (N2692)? N1665 : 
                 (N2694)? N1621 : 
                 (N2697)? decode_info_i[12] : 
                 (N2700)? N1666 : 
                 (N2703)? N1666 : 
                 (N1674)? 1'b0 : 1'b0;
  assign N93 = N1649;
  assign N1676 = (N94)? decode_info_i[10] : 
                 (N95)? 1'b0 : 
                 (N96)? 1'b0 : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N94 = N1533;
  assign N95 = N1541;
  assign N96 = N1550;
  assign N97 = N1556;
  assign N98 = N1563;
  assign N99 = N1588;
  assign N100 = N1602;
  assign N101 = N1603;
  assign N1677 = (N94)? decode_info_i[11] : 
                 (N95)? 1'b0 : 
                 (N96)? 1'b0 : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N1678 = (N94)? decode_info_i[12] : 
                 (N95)? 1'b0 : 
                 (N96)? 1'b0 : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N1679 = (N94)? 1'b0 : 
                 (N95)? N1612 : 
                 (N96)? 1'b0 : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N1680 = (N94)? 1'b0 : 
                 (N95)? N1613 : 
                 (N96)? 1'b0 : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N1681 = (N94)? 1'b0 : 
                 (N95)? 1'b0 : 
                 (N96)? N1614 : 
                 (N97)? N1666 : 
                 (N98)? N1616 : 
                 (N99)? decode_info_i[7] : 
                 (N100)? N1619 : 
                 (N101)? N1675 : 
                 (N1611)? 1'b1 : 1'b0;
  assign N1682 = (N94)? 1'b0 : 
                 (N95)? 1'b0 : 
                 (N96)? decode_info_i[9] : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N1683 = (N94)? 1'b0 : 
                 (N95)? 1'b0 : 
                 (N96)? 1'b0 : 
                 (N97)? N1615 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N1684 = (N94)? 1'b0 : 
                 (N95)? 1'b0 : 
                 (N96)? 1'b0 : 
                 (N97)? 1'b0 : 
                 (N98)? N1617 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N1685 = (N94)? 1'b0 : 
                 (N95)? 1'b0 : 
                 (N96)? 1'b0 : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? N1618 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign { N1689, N1688, N1687, N1686 } = (N94)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                          (N95)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                          (N96)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                          (N97)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                          (N98)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                          (N99)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                          (N100)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                          (N101)? { N2707, 1'b0, N1621, N1643 } : 
                                          (N1611)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1690 = (N94)? 1'b0 : 
                 (N95)? 1'b0 : 
                 (N96)? 1'b0 : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? N1620 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N1691 = (N102)? N1690 : 
                 (N103)? 1'b0 : 1'b0;
  assign N102 = N1518;
  assign N103 = N1517;
  assign N1692 = (N102)? N1676 : 
                 (N103)? 1'b0 : 1'b0;
  assign N1693 = (N102)? N1677 : 
                 (N103)? 1'b0 : 1'b0;
  assign N1694 = (N102)? N1678 : 
                 (N103)? 1'b0 : 1'b0;
  assign N1695 = (N102)? N1679 : 
                 (N103)? 1'b0 : 1'b0;
  assign N1696 = (N102)? N1680 : 
                 (N103)? 1'b0 : 1'b0;
  assign N1697 = (N102)? N1681 : 
                 (N103)? 1'b1 : 1'b0;
  assign N1698 = (N102)? N1682 : 
                 (N103)? 1'b0 : 1'b0;
  assign N1699 = (N102)? N1683 : 
                 (N103)? 1'b0 : 1'b0;
  assign N1700 = (N102)? N1684 : 
                 (N103)? 1'b0 : 1'b0;
  assign N1701 = (N102)? N1685 : 
                 (N103)? 1'b0 : 1'b0;
  assign { N1705, N1704, N1703, N1702 } = (N102)? { N1689, N1688, N1687, N1686 } : 
                                          (N103)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2256, N2255, N2254, N2253, N2252, N2251 } = (N104)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, N2048, 1'b0, 1'b0, 1'b0, 1'b0, N2061, 1'b0 } : 
                                                                                                                (N105)? { 1'b1, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, N2090, 1'b0, 1'b0, 1'b0, 1'b1, N1868, N2105 } : 
                                                                                                                (N106)? { 1'b1, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, N2124, 1'b0, 1'b0, 1'b1, 1'b1, N1868, N2134 } : 
                                                                                                                (N107)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, N2169, N1868, 1'b0, 1'b0, 1'b1, 1'b0, N2180, 1'b0 } : 
                                                                                                                (N108)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, N2199, N1868, 1'b0, 1'b1, 1'b0, 1'b0, N2209, 1'b0 } : 
                                                                                                                (N109)? { 1'b1, 1'b0, N2707, 1'b0, 1'b0, 1'b1, 1'b0, N2229, 1'b0, 1'b1, 1'b1, 1'b0, N1868, N2229 } : 
                                                                                                                (N110)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, N2250, N1868, 1'b0, 1'b1, 1'b0, 1'b1, N2250, 1'b0 } : 
                                                                                                                (N111)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, N1868, 1'b0, 1'b1, 1'b1, 1'b1, N1868, 1'b0 } : 
                                                                                                                (N112)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, N1868, 1'b1, 1'b0, 1'b0, 1'b0, N1868, 1'b0 } : 
                                                                                                                (N113)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, N1868, 1'b1, 1'b0, 1'b0, 1'b1, N1868, 1'b0 } : 
                                                                                                                (N114)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, N1868, 1'b1, 1'b1, 1'b1, 1'b0, N1868, 1'b0 } : 
                                                                                                                (N115)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, N1868, 1'b1, 1'b1, 1'b0, 1'b1, N1868, 1'b0 } : 
                                                                                                                (N116)? { 1'b1, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, N1868, 1'b1, 1'b0, 1'b1, 1'b0, N1868, 1'b0 } : 
                                                                                                                (N117)? { 1'b1, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, N1868, 1'b1, 1'b0, 1'b1, 1'b1, N1868, 1'b0 } : 
                                                                                                                (N118)? { 1'b1, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, N1868, 1'b1, 1'b1, 1'b0, 1'b0, N1868, 1'b0 } : 
                                                                                                                (N119)? { 1'b1, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, N1868, 1'b1, 1'b1, 1'b1, 1'b1, N1868, 1'b0 } : 
                                                                                                                (N120)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, N1868, 1'b0, 1'b0, 1'b0, 1'b0, N1868, 1'b0 } : 
                                                                                                                (N121)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, N1868, 1'b0, 1'b0, 1'b0, 1'b1, N1868, 1'b0 } : 
                                                                                                                (N122)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, N1868, 1'b0, 1'b0, 1'b1, 1'b0, N1868, 1'b0 } : 
                                                                                                                (N123)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, N1868, 1'b1, 1'b0, 1'b0, 1'b0, N1868, 1'b0 } : 
                                                                                                                (N124)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, N1868, 1'b1, 1'b0, 1'b0, 1'b1, N1868, 1'b0 } : 
                                                                                                                (N125)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1868, 1'b0, 1'b0, 1'b0, 1'b0, N1868, 1'b0 } : 1'b0;
  assign N104 = N1879;
  assign N105 = N1893;
  assign N106 = N1900;
  assign N107 = N1908;
  assign N108 = N1913;
  assign N109 = N1921;
  assign N110 = N1927;
  assign N111 = N1935;
  assign N112 = N1938;
  assign N113 = N1945;
  assign N114 = N1952;
  assign N115 = N1955;
  assign N116 = N1960;
  assign N117 = N1965;
  assign N118 = N1968;
  assign N119 = N1972;
  assign N120 = N1980;
  assign N121 = N1985;
  assign N122 = N1990;
  assign N123 = N1993;
  assign N124 = N2001;
  assign N125 = N2034;
  assign N2259 = (N104)? N2048 : 
                 (N2258)? N1868 : 1'b0;
  assign N2268 = (N104)? N2302 : 
                 (N105)? N2302 : 
                 (N106)? N2302 : 
                 (N107)? N2302 : 
                 (N108)? N2302 : 
                 (N109)? N2302 : 
                 (N110)? N2302 : 
                 (N111)? N2302 : 
                 (N112)? N2302 : 
                 (N113)? N2302 : 
                 (N114)? N2302 : 
                 (N115)? N2302 : 
                 (N116)? N2302 : 
                 (N117)? N2302 : 
                 (N118)? N2302 : 
                 (N119)? N2302 : 
                 (N120)? N2302 : 
                 (N121)? N2302 : 
                 (N122)? N2302 : 
                 (N123)? N2302 : 
                 (N124)? N2302 : 
                 (N125)? 1'b1 : 1'b0;
  assign { N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269 } = (N126)? { N2267, N2266, N2265, N2264, N2263, N2262, N1913, N2261, N2260, N2259, N2256, N2255, N2254, N2253, N2252, N2251 } : 
                                                                                                                              (N1873)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1868, N1868, 1'b0, 1'b0, 1'b0, 1'b0, N1868, 1'b0 } : 1'b0;
  assign N126 = N1872;
  assign N2285 = (N126)? N2268 : 
                 (N1873)? 1'b1 : 1'b0;
  assign { N2298, N2297, N2296 } = (N127)? { 1'b0, 1'b1, 1'b1 } : 
                                   (N128)? { 1'b1, 1'b0, 1'b0 } : 
                                   (N129)? { 1'b1, 1'b0, 1'b1 } : 
                                   (N130)? { 1'b1, 1'b1, 1'b0 } : 1'b0;
  assign N127 = N2290;
  assign N128 = N2292;
  assign N129 = N2294;
  assign N130 = N2295;
  assign { N2301, N2300, N2299 } = (N131)? { N2298, N2297, N2296 } : 
                                   (N2289)? { 1'b0, 1'b1, 1'b1 } : 1'b0;
  assign N131 = N2288;
  assign { N2373, N2372, N2371, N2370, N2369, N2368 } = (N132)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                                                        (N133)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                        (N134)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                                        (N135)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                                                        (N136)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                                                        (N137)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N138)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                                                        (N139)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                                        (N140)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                                        (N141)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                                        (N142)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                                                        (N143)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                        (N144)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                                                        (N145)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                                        (N146)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                                        (N147)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                                        (N148)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                        (N149)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                                        (N150)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N151)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                        (N152)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                                        (N153)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                                        (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N132 = N2341;
  assign N133 = N2343;
  assign N134 = N2344;
  assign N135 = N2346;
  assign N136 = N2347;
  assign N137 = N2348;
  assign N138 = N2350;
  assign N139 = N2352;
  assign N140 = N2353;
  assign N141 = N2354;
  assign N142 = N2355;
  assign N143 = N2356;
  assign N144 = N2357;
  assign N145 = N2358;
  assign N146 = N2359;
  assign N147 = N2360;
  assign N148 = N2361;
  assign N149 = N2362;
  assign N150 = N2363;
  assign N151 = N2364;
  assign N152 = N2365;
  assign N153 = N2366;
  assign N154 = N2367;
  assign N2374 = (N132)? 1'b0 : 
                 (N133)? 1'b0 : 
                 (N134)? 1'b0 : 
                 (N135)? 1'b0 : 
                 (N136)? 1'b0 : 
                 (N137)? 1'b0 : 
                 (N138)? 1'b0 : 
                 (N139)? 1'b0 : 
                 (N140)? 1'b0 : 
                 (N141)? 1'b0 : 
                 (N142)? 1'b0 : 
                 (N143)? 1'b0 : 
                 (N144)? 1'b0 : 
                 (N145)? 1'b0 : 
                 (N146)? 1'b0 : 
                 (N147)? 1'b0 : 
                 (N148)? 1'b0 : 
                 (N149)? 1'b0 : 
                 (N150)? 1'b0 : 
                 (N151)? 1'b0 : 
                 (N152)? 1'b0 : 
                 (N153)? 1'b0 : 
                 (N154)? 1'b1 : 1'b0;
  assign { N2380, N2379, N2378, N2377, N2376, N2375 } = (N155)? { N2373, N2372, N2371, N2370, N2369, N2368 } : 
                                                        (N2338)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N155 = N2337;
  assign N2381 = (N155)? N2374 : 
                 (N2338)? 1'b1 : 1'b0;
  assign N2470 = (N156)? 1'b0 : 
                 (N157)? 1'b0 : 
                 (N158)? 1'b0 : 
                 (N159)? 1'b0 : 
                 (N160)? N2381 : 1'b0;
  assign N156 = N2407;
  assign N157 = N2412;
  assign N158 = N2430;
  assign N159 = N2456;
  assign N160 = N2469;
  assign { N2527, N2526, N2519, N2518, N2517, N2516, N2509, N2508, N2507, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2489, N2488, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471 } = (N178)? { N349, 1'b0, 1'b0, N347, N2707, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N347, 1'b0, 1'b0, N803, N479, N413, N414, 1'b0, 1'b0, N720, N719, 1'b0, N718, N717, N716, 1'b0, N392, N990, N989, N988, N938, N937, N936 } : 
                                                                                                                                                                                                                                                     (N186)? { 1'b1, 1'b0, 1'b0, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1326, N1263, N1026, N1025, 1'b0, 1'b0, N1130, N1129, 1'b0, N1128, N1127, N1126, 1'b0, N1002, N1310, N1309, N1308, N1307, N1306, 1'b0 } : 
                                                                                                                                                                                                                                                     (N190)? { 1'b1, 1'b0, 1'b0, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N192)? { 1'b1, 1'b0, 1'b0, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N196)? { 1'b1, 1'b0, 1'b0, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N200)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1372, N1371, N1370, N1369, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                                                                     (N161)? { 1'b0, 1'b1, 1'b0, 1'b0, N2707, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1384, N1383, N1382, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N211)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1400, 1'b0, 1'b0, 1'b0, N1400, N1402, N1395, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N215)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1408, 1'b0, N1417, N1416, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N217)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1422, 1'b0, 1'b0, N1422, 1'b0, N1424, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N220)? { 1'b0, N1512, 1'b0, 1'b0, 1'b0, 1'b0, N1515, 1'b0, N1514, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1512, N1512, N1511, N1510, N1509, N1508, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N223)? { 1'b0, 1'b0, 1'b0, 1'b0, N1705, 1'b0, N1704, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N227)? { 1'b0, 1'b0, N2283, N2280, N2282, N2281, 1'b0, 1'b0, 1'b0, 1'b0, N2280, 1'b0, N2279, 1'b0, N2278, 1'b0, N2277, N2276, N2275, 1'b0, 1'b0, N2274, N2273, N2272, N2271, N2270, N2269, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N234)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N2709, N2709, 1'b0, 1'b0, 1'b0, N2301, N2300, N2299, N2709, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N238)? { 1'b0, 1'b1, 1'b0, 1'b0, N2707, 1'b0, 1'b0, N2333, N2334, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N2380, N2379, N2378, N2377, N2376, N2375, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N249)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N161 = N209;
  assign N2487 = (N234)? N2709 : 
                 (N2486)? 1'b0 : 1'b0;
  assign { N2520, N2493, N2492 } = (N178)? { N266, N538, N392 } : 
                                   (N2491)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N2521, N2504, N2503 } = (N223)? { 1'b1, N1703, N1702 } : 
                                   (N2502)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2506 = (N220)? N1513 : 
                 (N2505)? 1'b0 : 1'b0;
  assign { N2513, N2512 } = (N196)? { N1337, N1347 } : 
                            (N2511)? { 1'b0, 1'b0 } : 1'b0;
  assign N2515 = (N200)? 1'b1 : 
                 (N2514)? 1'b0 : 1'b0;
  assign N2523 = (N211)? 1'b1 : 
                 (N2522)? 1'b0 : 1'b0;
  assign N2525 = (N227)? N2284 : 
                 (N2524)? 1'b0 : 1'b0;
  assign N2528 = (N178)? N721 : 
                 (N186)? N1131 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? N1349 : 
                 (N200)? N1373 : 
                 (N161)? N1385 : 
                 (N211)? N1403 : 
                 (N215)? N1418 : 
                 (N217)? N1425 : 
                 (N220)? N1507 : 
                 (N223)? N1697 : 
                 (N227)? N2285 : 
                 (N234)? N2302 : 
                 (N238)? N2470 : 
                 (N249)? 1'b1 : 1'b0;
  assign N2529 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? N1506 : 
                 (N223)? 1'b0 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2530 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1700 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2531 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1701 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2532 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1691 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2533 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1703 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2534 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1692 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2535 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1693 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2536 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1694 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2537 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1695 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2538 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1696 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2539 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1698 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2540 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1699 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign dret_o = (N162)? N2539 : 
                  (N174)? 1'b0 : 1'b0;
  assign N162 = N173;
  assign mret_o = (N162)? N2540 : 
                  (N174)? 1'b0 : 1'b0;
  assign { decode_o[53:46], decode_o[40:32], decode_o[30:20], decode_o[18:8], decode_o[6:0] } = (N162)? { N2527, N2526, N2525, N2523, N2521, N2520, N2519, N2518, N2517, N2516, N2515, N2513, N2512, N2509, N2508, N2507, N2506, N2504, N2503, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2489, N2488, N2487, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471 } : 
                                                                                                (N174)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign illegal_instr_o = (N162)? N2528 : 
                           (N174)? 1'b1 : 1'b0;
  assign fencei_o = (N162)? N2529 : 
                    (N174)? 1'b0 : 1'b0;
  assign sret_o = (N162)? N2530 : 
                  (N174)? 1'b0 : 1'b0;
  assign wfi_o = (N162)? N2531 : 
                 (N174)? 1'b0 : 1'b0;
  assign sfence_vma_o = (N162)? N2532 : 
                        (N174)? 1'b0 : 1'b0;
  assign csrw_o = (N162)? N2533 : 
                  (N174)? 1'b0 : 1'b0;
  assign ecall_m_o = (N162)? N2534 : 
                     (N174)? 1'b0 : 1'b0;
  assign ecall_s_o = (N162)? N2535 : 
                     (N174)? 1'b0 : 1'b0;
  assign ecall_u_o = (N162)? N2536 : 
                     (N174)? 1'b0 : 1'b0;
  assign dbreak_o = (N162)? N2537 : 
                    (N174)? 1'b0 : 1'b0;
  assign ebreak_o = (N162)? N2538 : 
                    (N174)? 1'b0 : 1'b0;
  assign { N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579 } = (N163)? { preissue_pkt_i[33:14], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                              (N164)? { preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[21:14], preissue_pkt_i[22:22], preissue_pkt_i[32:23], 1'b0 } : 
                                                                                                                                                                                                                                              (N165)? { preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[9:9], preissue_pkt_i[32:27], preissue_pkt_i[13:10], 1'b0 } : 
                                                                                                                                                                                                                                              (N166)? { preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:27], preissue_pkt_i[13:9] } : 
                                                                                                                                                                                                                                              (N167)? { preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:22] } : 
                                                                                                                                                                                                                                              (N168)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N163 = N2547;
  assign N164 = N2552;
  assign N165 = N2555;
  assign N166 = N2559;
  assign N167 = N2570;
  assign N168 = N2578;
  assign { N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611 } = (N162)? { N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579 } : 
                                                                                                                                                                                                                                              (N174)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign imm_o = (N169)? { N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N1287, N462, N2303, N393, N2684, N523, N2685, N2686, N1183, N2079, N2035 } : 
                 (N170)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                 (N171)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                 (N172)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                 (N2683)? { N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611 } : 1'b0;
  assign N169 = N2649;
  assign N170 = N2657;
  assign N171 = N2665;
  assign N172 = N2679;
  assign N174 = ~N173;
  assign N178 = N2728 | N2729;
  assign N2728 = ~N175;
  assign N2729 = ~N177;
  assign N186 = N2730 | N2731;
  assign N2730 = ~N182;
  assign N2731 = ~N185;
  assign N190 = ~N189;
  assign N192 = ~N191;
  assign N196 = N2732 | N2733;
  assign N2732 = ~N194;
  assign N2733 = ~N195;
  assign N200 = ~N199;
  assign N201 = ~preissue_pkt_i[8];
  assign N202 = ~preissue_pkt_i[7];
  assign N203 = ~preissue_pkt_i[6];
  assign N204 = ~preissue_pkt_i[5];
  assign N205 = ~preissue_pkt_i[4];
  assign N211 = ~N210;
  assign N215 = ~N214;
  assign N217 = ~N216;
  assign N220 = ~N219;
  assign N223 = ~N222;
  assign N227 = ~N226;
  assign N234 = N2738 | N2739;
  assign N2738 = N2736 | N2737;
  assign N2736 = N2734 | N2735;
  assign N2734 = ~N229;
  assign N2735 = ~N230;
  assign N2737 = ~N232;
  assign N2739 = ~N233;
  assign N238 = ~N237;
  assign N249 = N240 | N2742;
  assign N2742 = N242 | N2741;
  assign N2741 = N243 | N2740;
  assign N2740 = N246 | N248;
  assign N348 = N347 | N266;
  assign N546 = ~N545;
  assign N580 = N2758 | N579;
  assign N2758 = N2757 | N578;
  assign N2757 = N2756 | N577;
  assign N2756 = N2755 | N576;
  assign N2755 = N2754 | N574;
  assign N2754 = N2753 | N573;
  assign N2753 = N2752 | N571;
  assign N2752 = N2751 | N570;
  assign N2751 = N2750 | N568;
  assign N2750 = N2749 | N566;
  assign N2749 = N2748 | N564;
  assign N2748 = N2747 | N563;
  assign N2747 = N2746 | N561;
  assign N2746 = N2745 | N560;
  assign N2745 = N2744 | N558;
  assign N2744 = N2743 | N554;
  assign N2743 = N549 | N552;
  assign N603 = N601 | N602;
  assign N611 = N2762 | N610;
  assign N2762 = N2761 | N609;
  assign N2761 = N2760 | N608;
  assign N2760 = N2759 | N607;
  assign N2759 = N605 | N606;
  assign N614 = N612 | N613;
  assign N630 = N628 | N629;
  assign N639 = N637 | N638;
  assign N642 = N640 | N641;
  assign N645 = N643 | N644;
  assign N649 = N646 | N648;
  assign N709 = N652 | N2791;
  assign N2791 = N656 | N2790;
  assign N2790 = N658 | N2789;
  assign N2789 = N660 | N2788;
  assign N2788 = N662 | N2787;
  assign N2787 = N664 | N2786;
  assign N2786 = N665 | N2785;
  assign N2785 = N667 | N2784;
  assign N2784 = N669 | N2783;
  assign N2783 = N671 | N2782;
  assign N2782 = N673 | N2781;
  assign N2781 = N675 | N2780;
  assign N2780 = N678 | N2779;
  assign N2779 = N680 | N2778;
  assign N2778 = N681 | N2777;
  assign N2777 = N682 | N2776;
  assign N2776 = N685 | N2775;
  assign N2775 = N687 | N2774;
  assign N2774 = N689 | N2773;
  assign N2773 = N691 | N2772;
  assign N2772 = N694 | N2771;
  assign N2771 = N695 | N2770;
  assign N2770 = N699 | N2769;
  assign N2769 = N700 | N2768;
  assign N2768 = N701 | N2767;
  assign N2767 = N702 | N2766;
  assign N2766 = N703 | N2765;
  assign N2765 = N704 | N2764;
  assign N2764 = N706 | N2763;
  assign N2763 = N707 | N708;
  assign N834 = ~N833;
  assign N853 = ~N852;
  assign N891 = ~N890;
  assign N908 = ~N907;
  assign N927 = ~N926;
  assign N987 = ~N986;
  assign N1023 = N1022 | N1006;
  assign N1024 = ~N1023;
  assign N1030 = ~N1029;
  assign N1052 = N2800 | N1051;
  assign N2800 = N2799 | N1050;
  assign N2799 = N2798 | N1047;
  assign N2798 = N2797 | N1045;
  assign N2797 = N2796 | N1043;
  assign N2796 = N2795 | N1042;
  assign N2795 = N2794 | N1040;
  assign N2794 = N2793 | N1038;
  assign N2793 = N2792 | N1037;
  assign N2792 = N1031 | N1032;
  assign N1062 = N2801 | N597;
  assign N2801 = N1057 | N1061;
  assign N1067 = N1064 | N1066;
  assign N1080 = N2803 | N1079;
  assign N2803 = N2802 | N1077;
  assign N2802 = N1071 | N1074;
  assign N1106 = N1053 | N1052;
  assign N1107 = N1054 | N1106;
  assign N1108 = N593 | N1107;
  assign N1109 = N1062 | N1108;
  assign N1110 = N599 | N1109;
  assign N1111 = N1067 | N1110;
  assign N1112 = N1080 | N1111;
  assign N1113 = N1086 | N1112;
  assign N1114 = N1093 | N1113;
  assign N1115 = N1095 | N1114;
  assign N1116 = N1098 | N1115;
  assign N1117 = N1101 | N1116;
  assign N1118 = N1105 | N1117;
  assign N1119 = ~N1118;
  assign N1211 = ~N1210;
  assign N1231 = ~N1230;
  assign N1258 = ~N1257;
  assign N1305 = ~N1304;
  assign N1349 = ~N1348;
  assign N1353 = ~N1352;
  assign N1375 = ~N1374;
  assign N1401 = ~N1400;
  assign N1409 = ~N1408;
  assign N1423 = ~N1422;
  assign N1428 = ~N1427;
  assign N1486 = N1434 | N1431;
  assign N1487 = N1437 | N1486;
  assign N1488 = N1440 | N1487;
  assign N1489 = N1445 | N1488;
  assign N1490 = N1448 | N1489;
  assign N1491 = N1452 | N1490;
  assign N1492 = N1455 | N1491;
  assign N1493 = N1469 | N1492;
  assign N1494 = N1473 | N1493;
  assign N1495 = N1476 | N1494;
  assign N1496 = N1485 | N1495;
  assign N1518 = ~N1517;
  assign N1519 = ~preissue_pkt_i[21];
  assign N1520 = ~preissue_pkt_i[20];
  assign N1521 = ~preissue_pkt_i[19];
  assign N1522 = ~preissue_pkt_i[18];
  assign N1523 = ~preissue_pkt_i[17];
  assign N1541 = ~N1540;
  assign N1550 = ~N1549;
  assign N1556 = ~N1555;
  assign N1563 = ~N1562;
  assign N1588 = ~N1587;
  assign N1589 = ~preissue_pkt_i[13];
  assign N1590 = ~preissue_pkt_i[12];
  assign N1591 = ~preissue_pkt_i[11];
  assign N1592 = ~preissue_pkt_i[10];
  assign N1593 = ~preissue_pkt_i[9];
  assign N1603 = N2807 | N1362;
  assign N2807 = N2806 | N1377;
  assign N2806 = N2805 | N1361;
  assign N2805 = N2804 | N1376;
  assign N2804 = N1356 | N1359;
  assign N1604 = N1541 | N1533;
  assign N1605 = N1550 | N1604;
  assign N1606 = N1556 | N1605;
  assign N1607 = N1563 | N1606;
  assign N1608 = N1588 | N1607;
  assign N1609 = N1602 | N1608;
  assign N1610 = N1603 | N1609;
  assign N1611 = ~N1610;
  assign N1612 = N2811 | N2812;
  assign N2811 = N2809 | N2810;
  assign N2809 = decode_info_i[9] | N2808;
  assign N2808 = decode_info_i[5] & decode_info_i[10];
  assign N2810 = decode_info_i[4] & decode_info_i[11];
  assign N2812 = decode_info_i[3] & decode_info_i[12];
  assign N1613 = ~N1612;
  assign N1614 = ~decode_info_i[9];
  assign N1615 = ~N1666;
  assign N1616 = decode_info_i[12] | N2813;
  assign N2813 = decode_info_i[8] & decode_info_i[11];
  assign N1617 = ~N1616;
  assign N1618 = N2814 & N1614;
  assign N2814 = ~decode_info_i[7];
  assign N1619 = N2815 | decode_info_i[12];
  assign N2815 = decode_info_i[11] & decode_info_i[6];
  assign N1620 = ~N1619;
  assign N1621 = N1642 | N2727;
  assign N1643 = N2816 | N2707;
  assign N2816 = ~N1642;
  assign N1649 = N2819 | N2820;
  assign N2819 = N2817 | N2818;
  assign N2817 = ~N1646;
  assign N2818 = ~N1647;
  assign N2820 = ~N1648;
  assign N1651 = ~N1650;
  assign N1656 = ~N1655;
  assign N1662 = ~N1661;
  assign N1663 = ~decode_info_i[1];
  assign N1664 = ~decode_info_i[0];
  assign N1665 = decode_info_i[11] & decode_info_i[6];
  assign N1666 = decode_info_i[11] | decode_info_i[12];
  assign N1667 = N2688 | N1649;
  assign N1668 = N2690 | N1667;
  assign N1669 = N2692 | N1668;
  assign N1670 = N2694 | N1669;
  assign N1671 = N2697 | N1670;
  assign N1672 = N2700 | N1671;
  assign N1673 = N2703 | N1672;
  assign N1674 = ~N1673;
  assign N1873 = ~N1872;
  assign N1879 = N1876 | N1878;
  assign N1893 = N2822 | N1892;
  assign N2822 = N2821 | N1891;
  assign N2821 = N1885 | N1888;
  assign N1900 = N2824 | N1899;
  assign N2824 = N2823 | N1898;
  assign N2823 = N1895 | N1897;
  assign N1908 = N2826 | N1907;
  assign N2826 = N2825 | N1906;
  assign N2825 = N1903 | N1904;
  assign N1913 = N2828 | N1912;
  assign N2828 = N2827 | N1911;
  assign N2827 = N1909 | N1910;
  assign N1921 = N1918 | N1920;
  assign N1927 = N1924 | N1926;
  assign N1935 = N1931 | N1934;
  assign N1938 = N1936 | N1937;
  assign N1945 = N1941 | N1944;
  assign N1952 = N1948 | N1951;
  assign N1955 = N1953 | N1954;
  assign N1960 = N1957 | N1959;
  assign N1965 = N1962 | N1964;
  assign N1968 = N1966 | N1967;
  assign N1972 = N1970 | N1971;
  assign N1980 = N1977 | N1979;
  assign N1985 = N1981 | N1984;
  assign N1990 = N1988 | N1989;
  assign N1993 = N1991 | N1992;
  assign N2001 = N1997 | N2000;
  assign N2034 = N2004 | N2852;
  assign N2852 = N2007 | N2851;
  assign N2851 = N2008 | N2850;
  assign N2850 = N2009 | N2849;
  assign N2849 = N2010 | N2848;
  assign N2848 = N2012 | N2847;
  assign N2847 = N2013 | N2846;
  assign N2846 = N2014 | N2845;
  assign N2845 = N2015 | N2844;
  assign N2844 = N2016 | N2843;
  assign N2843 = N2017 | N2842;
  assign N2842 = N2019 | N2841;
  assign N2841 = N2020 | N2840;
  assign N2840 = N2021 | N2839;
  assign N2839 = N2024 | N2838;
  assign N2838 = N2025 | N2837;
  assign N2837 = N682 | N2836;
  assign N2836 = N2459 | N2835;
  assign N2835 = N2026 | N2834;
  assign N2834 = N2028 | N2833;
  assign N2833 = N2029 | N2832;
  assign N2832 = N2030 | N2831;
  assign N2831 = N2031 | N2830;
  assign N2830 = N2032 | N2829;
  assign N2829 = N2033 | N662;
  assign N2257 = ~N1879;
  assign N2258 = N2257;
  assign N2289 = ~N2288;
  assign N2292 = ~N2291;
  assign N2294 = ~N2293;
  assign N2302 = ~decode_info_i[2];
  assign N2334 = ~N2333;
  assign N2338 = ~N2337;
  assign N2367 = N2457 | N2861;
  assign N2861 = N2458 | N2860;
  assign N2860 = N2459 | N2859;
  assign N2859 = N2460 | N2858;
  assign N2858 = N2461 | N2857;
  assign N2857 = N2462 | N2856;
  assign N2856 = N2464 | N2855;
  assign N2855 = N2465 | N2854;
  assign N2854 = N2466 | N2853;
  assign N2853 = N2467 | N2468;
  assign N2407 = N2863 | N2406;
  assign N2863 = N2862 | N2403;
  assign N2862 = N2392 | N2397;
  assign N2412 = N2409 | N2411;
  assign N2430 = N2867 | N2429;
  assign N2867 = N2866 | N2427;
  assign N2866 = N2865 | N2424;
  assign N2865 = N2864 | N2422;
  assign N2864 = N2416 | N2419;
  assign N2456 = N2875 | N2455;
  assign N2875 = N2874 | N2453;
  assign N2874 = N2873 | N2450;
  assign N2873 = N2872 | N2448;
  assign N2872 = N2871 | N2444;
  assign N2871 = N2870 | N2442;
  assign N2870 = N2869 | N2439;
  assign N2869 = N2868 | N2437;
  assign N2868 = N2432 | N2434;
  assign N2469 = preissue_pkt_i[16] | N2893;
  assign N2893 = N2304 | N2892;
  assign N2892 = preissue_pkt_i[8] | N2891;
  assign N2891 = N1328 | N2890;
  assign N2890 = preissue_pkt_i[6] | N2889;
  assign N2889 = N1329 | N2888;
  assign N2888 = N1330 | N2887;
  assign N2887 = N395 | N2886;
  assign N2886 = N396 | N2885;
  assign N2885 = N2457 | N2884;
  assign N2884 = N2458 | N2883;
  assign N2883 = N2459 | N2882;
  assign N2882 = N2460 | N2881;
  assign N2881 = N2461 | N2880;
  assign N2880 = N2462 | N2879;
  assign N2879 = N2464 | N2878;
  assign N2878 = N2465 | N2877;
  assign N2877 = N2466 | N2876;
  assign N2876 = N2467 | N2468;
  assign N2485 = ~N234;
  assign N2486 = N2485;
  assign N2490 = ~N178;
  assign N2491 = N2490;
  assign N2502 = N222;
  assign N2505 = N219;
  assign N2510 = ~N196;
  assign N2511 = N2510;
  assign N2514 = N199;
  assign N2522 = N210;
  assign N2524 = N226;
  assign N2547 = N2894 | N2895;
  assign N2894 = ~N2544;
  assign N2895 = ~N2546;
  assign N2552 = ~N2551;
  assign N2555 = ~N2554;
  assign N2559 = N2896 | N2897;
  assign N2896 = ~N2557;
  assign N2897 = ~N2558;
  assign N2570 = N2903 | N2904;
  assign N2903 = N2901 | N2902;
  assign N2901 = N2899 | N2900;
  assign N2899 = N2898 | N2563;
  assign N2898 = ~N2560;
  assign N2900 = ~N2564;
  assign N2902 = ~N2567;
  assign N2904 = ~N2569;
  assign N2578 = N240 | N2908;
  assign N2908 = N2572 | N2907;
  assign N2907 = N241 | N2906;
  assign N2906 = N2574 | N2905;
  assign N2905 = N2576 | N2577;
  assign N2649 = N2645 | N2648;
  assign N2657 = N2654 | N2656;
  assign N2665 = N2661 | N2664;
  assign N2679 = N2674 | N2678;
  assign N2680 = N2657 | N2649;
  assign N2681 = N2665 | N2680;
  assign N2682 = N2679 | N2681;
  assign N2683 = ~N2682;
  assign N2684 = ~preissue_pkt_i[28];
  assign N2685 = ~preissue_pkt_i[26];
  assign N2686 = ~preissue_pkt_i[25];
  assign N2687 = ~N1649;
  assign N2688 = N1651 & N2687;
  assign N2689 = N2687 & N1650;
  assign N2690 = N1656 & N2689;
  assign N2691 = N2689 & N1655;
  assign N2692 = N1662 & N2691;
  assign N2693 = N2691 & N1661;
  assign N2694 = N2445 & N2693;
  assign N2695 = ~N2445;
  assign N2696 = N2693 & N2695;
  assign N2697 = N1986 & N2696;
  assign N2698 = ~N1986;
  assign N2699 = N2696 & N2698;
  assign N2700 = N2005 & N2699;
  assign N2701 = ~N2005;
  assign N2702 = N2699 & N2701;
  assign N2703 = N2457 & N2702;

endmodule



module bp_be_issue_queue_00
(
  clk_i,
  reset_i,
  en_i,
  clr_i,
  roll_i,
  read_i,
  read_cnt_i,
  read_size_i,
  cmt_i,
  cmt_cnt_i,
  cmt_size_i,
  fe_queue_i,
  fe_queue_v_i,
  fe_queue_ready_and_o,
  decode_info_i,
  preissue_pkt_o,
  issue_pkt_o
);

  input [3:0] read_cnt_i;
  input [3:0] read_size_i;
  input [3:0] cmt_cnt_i;
  input [3:0] cmt_size_i;
  input [173:0] fe_queue_i;
  input [12:0] decode_info_i;
  output [38:0] preissue_pkt_o;
  output [263:0] issue_pkt_o;
  input clk_i;
  input reset_i;
  input en_i;
  input clr_i;
  input roll_i;
  input read_i;
  input cmt_i;
  input fe_queue_v_i;
  output fe_queue_ready_and_o;
  wire [38:0] preissue_pkt_o;
  wire [263:0] issue_pkt_o;
  wire fe_queue_ready_and_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,
  N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,
  N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,ack,empty,empty_n,N69,N70,full,
  N71,N72,N73,N74,read_catchup,N75,N76,N77,N78,deq_catchup,N79,N80,N81,N82,N83,N84,
  N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,
  N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,
  N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,
  N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,
  N152,preissue_v,bypass_preissue,_0_net_,_2_net_,N153,queue_instr_raw_4__15_,
  queue_instr_raw_4__14_,queue_instr_raw_4__13_,queue_instr_raw_4__12_,
  queue_instr_raw_4__11_,queue_instr_raw_4__10_,queue_instr_raw_4__9_,queue_instr_raw_4__8_,
  queue_instr_raw_4__7_,queue_instr_raw_4__6_,queue_instr_raw_4__5_,
  queue_instr_raw_4__4_,queue_instr_raw_4__3_,queue_instr_raw_4__2_,queue_instr_raw_4__1_,
  queue_instr_raw_4__0_,queue_instr_raw_3__15_,queue_instr_raw_3__14_,queue_instr_raw_3__13_,
  queue_instr_raw_3__12_,queue_instr_raw_3__11_,queue_instr_raw_3__10_,
  queue_instr_raw_3__9_,queue_instr_raw_3__8_,queue_instr_raw_3__7_,queue_instr_raw_3__6_,
  queue_instr_raw_3__5_,queue_instr_raw_3__4_,queue_instr_raw_3__3_,
  queue_instr_raw_3__2_,queue_instr_raw_3__1_,queue_instr_raw_3__0_,queue_instr_raw_2__15_,
  queue_instr_raw_2__14_,queue_instr_raw_2__13_,queue_instr_raw_2__12_,
  queue_instr_raw_2__11_,queue_instr_raw_2__10_,queue_instr_raw_2__9_,queue_instr_raw_2__8_,
  queue_instr_raw_2__7_,queue_instr_raw_2__6_,queue_instr_raw_2__5_,queue_instr_raw_2__4_,
  queue_instr_raw_2__3_,queue_instr_raw_2__2_,queue_instr_raw_2__1_,
  queue_instr_raw_2__0_,queue_instr_raw_1__15_,queue_instr_raw_1__14_,queue_instr_raw_1__13_,
  queue_instr_raw_1__12_,queue_instr_raw_1__11_,queue_instr_raw_1__10_,
  queue_instr_raw_1__9_,queue_instr_raw_1__8_,queue_instr_raw_1__7_,queue_instr_raw_1__6_,
  queue_instr_raw_1__5_,queue_instr_raw_1__4_,queue_instr_raw_1__3_,queue_instr_raw_1__2_,
  queue_instr_raw_1__1_,queue_instr_raw_1__0_,queue_instr_raw_0__15_,
  queue_instr_raw_0__14_,queue_instr_raw_0__13_,queue_instr_raw_0__12_,queue_instr_raw_0__11_,
  queue_instr_raw_0__10_,queue_instr_raw_0__9_,queue_instr_raw_0__8_,
  queue_instr_raw_0__7_,queue_instr_raw_0__6_,queue_instr_raw_0__5_,queue_instr_raw_0__4_,
  queue_instr_raw_0__3_,queue_instr_raw_0__2_,queue_instr_raw_0__1_,
  queue_instr_raw_0__0_,N154,preissue_size_4__1_,preissue_size_4__0_,preissue_size_3__1_,
  preissue_size_3__0_,preissue_size_2__1_,preissue_size_2__0_,preissue_size_1__1_,
  preissue_size_1__0_,preissue_size_0__1_,preissue_size_0__0_,N155,N156,N157,N158,N159,N160,
  N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,
  N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,
  N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,
  N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,
  N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,
  N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,
  N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,
  N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
  N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,
  N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
  N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,
  N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,
  N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,
  N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,
  N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,
  N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,
  N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,
  N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,
  N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,
  N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,
  N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,
  N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,
  N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,
  N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,
  N593,N594,N595,N596,N597,N598,N599,preissue_pkt_r_irs1_v_,preissue_pkt_r_irs2_v_,
  preissue_pkt_r_frs1_v_,preissue_pkt_r_frs2_v_,preissue_pkt_r_frs3_v_,
  preissue_pkt_r_size__1_,preissue_pkt_r_size__0_,bypass_issue,_4_net_,_6_net_,
  fe_queue_lo_pc__38_,fe_queue_lo_pc__37_,fe_queue_lo_pc__36_,fe_queue_lo_pc__35_,
  fe_queue_lo_pc__34_,fe_queue_lo_pc__33_,fe_queue_lo_pc__32_,fe_queue_lo_pc__31_,
  fe_queue_lo_pc__30_,fe_queue_lo_pc__29_,fe_queue_lo_pc__28_,fe_queue_lo_pc__27_,
  fe_queue_lo_pc__26_,fe_queue_lo_pc__25_,fe_queue_lo_pc__24_,fe_queue_lo_pc__23_,
  fe_queue_lo_pc__22_,fe_queue_lo_pc__21_,fe_queue_lo_pc__20_,fe_queue_lo_pc__19_,
  fe_queue_lo_pc__18_,fe_queue_lo_pc__17_,fe_queue_lo_pc__16_,fe_queue_lo_pc__15_,
  fe_queue_lo_pc__14_,fe_queue_lo_pc__13_,fe_queue_lo_pc__12_,fe_queue_lo_pc__11_,
  fe_queue_lo_pc__10_,fe_queue_lo_pc__9_,fe_queue_lo_pc__8_,fe_queue_lo_pc__7_,fe_queue_lo_pc__6_,
  fe_queue_lo_pc__5_,fe_queue_lo_pc__4_,fe_queue_lo_pc__3_,fe_queue_lo_pc__2_,
  fe_queue_lo_pc__1_,fe_queue_lo_pc__0_,fe_queue_lo_instr__79_,fe_queue_lo_instr__78_,
  fe_queue_lo_instr__77_,fe_queue_lo_instr__76_,fe_queue_lo_instr__75_,
  fe_queue_lo_instr__74_,fe_queue_lo_instr__73_,fe_queue_lo_instr__72_,
  fe_queue_lo_instr__71_,fe_queue_lo_instr__70_,fe_queue_lo_instr__69_,fe_queue_lo_instr__68_,
  fe_queue_lo_instr__67_,fe_queue_lo_instr__66_,fe_queue_lo_instr__65_,
  fe_queue_lo_instr__64_,fe_queue_lo_instr__63_,fe_queue_lo_instr__62_,fe_queue_lo_instr__61_,
  fe_queue_lo_instr__60_,fe_queue_lo_instr__59_,fe_queue_lo_instr__58_,
  fe_queue_lo_instr__57_,fe_queue_lo_instr__56_,fe_queue_lo_instr__55_,fe_queue_lo_instr__54_,
  fe_queue_lo_instr__53_,fe_queue_lo_instr__52_,fe_queue_lo_instr__51_,
  fe_queue_lo_instr__50_,fe_queue_lo_instr__49_,fe_queue_lo_instr__48_,fe_queue_lo_instr__47_,
  fe_queue_lo_instr__46_,fe_queue_lo_instr__45_,fe_queue_lo_instr__44_,
  fe_queue_lo_instr__43_,fe_queue_lo_instr__42_,fe_queue_lo_instr__41_,fe_queue_lo_instr__40_,
  fe_queue_lo_instr__39_,fe_queue_lo_instr__38_,fe_queue_lo_instr__37_,
  fe_queue_lo_instr__36_,fe_queue_lo_instr__35_,fe_queue_lo_instr__34_,fe_queue_lo_instr__33_,
  fe_queue_lo_instr__32_,fe_queue_lo_instr__31_,fe_queue_lo_instr__30_,
  fe_queue_lo_instr__29_,fe_queue_lo_instr__28_,fe_queue_lo_instr__27_,fe_queue_lo_instr__26_,
  fe_queue_lo_instr__25_,fe_queue_lo_instr__24_,fe_queue_lo_instr__23_,
  fe_queue_lo_instr__22_,fe_queue_lo_instr__21_,fe_queue_lo_instr__20_,fe_queue_lo_instr__19_,
  fe_queue_lo_instr__18_,fe_queue_lo_instr__17_,fe_queue_lo_instr__16_,
  fe_queue_lo_instr__15_,fe_queue_lo_instr__14_,fe_queue_lo_instr__13_,fe_queue_lo_instr__12_,
  fe_queue_lo_instr__11_,fe_queue_lo_instr__10_,fe_queue_lo_instr__9_,
  fe_queue_lo_instr__8_,fe_queue_lo_instr__7_,fe_queue_lo_instr__6_,fe_queue_lo_instr__5_,
  fe_queue_lo_instr__4_,fe_queue_lo_instr__3_,fe_queue_lo_instr__2_,
  fe_queue_lo_instr__1_,fe_queue_lo_instr__0_,fe_queue_lo_msg_type__2_,fe_queue_lo_msg_type__1_,
  fe_queue_lo_msg_type__0_,N600,illegal_instr_lo,N601,N602,N604,N605,N606,N608,N609,
  N610,N612,N613,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,
  N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,
  N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,
  N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,
  N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,
  N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,
  N708,N709,N710,N711,N712,N713,N714;
  wire [6:0] rptr_r,wptr_r,rptr_n,wptr_n,cptr_r,cptr_n,rptr_jmp,wptr_jmp,cptr_jmp;
  wire [3:0] enq,read,deq;
  wire [79:0] queue_instr_n;
  wire [2:0] preissue_entry_sel;
  wire [31:0] \e_0_.instr ,\e_1_.instr ,\e_2_.instr ,\e_3_.instr ,\e_4_.instr ;
  wire [159:0] preissue_instr;
  assign issue_pkt_o[113] = 1'b0;
  assign issue_pkt_o[114] = 1'b0;
  assign empty = rptr_r == wptr_r;
  assign empty_n = rptr_n == wptr_n;
  assign N69 = cptr_r[5:3] == wptr_r[5:3];
  assign N70 = cptr_r[6] ^ wptr_r[6];
  assign read_catchup = { N74, N73, N72, N71 } >= read_cnt_i;
  assign deq_catchup = { N78, N77, N76, N75 } >= cmt_cnt_i;

  bsg_circular_ptr_slots_p128_max_add_p127
  cptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(cptr_jmp),
    .o(cptr_r),
    .n_o(cptr_n)
  );


  bsg_circular_ptr_slots_p128_max_add_p127
  wptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(wptr_jmp),
    .o(wptr_r),
    .n_o(wptr_n)
  );


  bsg_circular_ptr_slots_p128_max_add_p127
  rptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(rptr_jmp),
    .o(rptr_r),
    .n_o(rptr_n)
  );

  assign bypass_preissue = wptr_r == rptr_n;

  bsg_mem_1r1w_00000050_00000008
  preissue_fifo_mem
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(_0_net_),
    .w_addr_i(wptr_r[5:3]),
    .w_data_i(fe_queue_i[134:55]),
    .r_v_i(_2_net_),
    .r_addr_i(rptr_n[5:3]),
    .r_data_o(queue_instr_n)
  );


  bp_be_expander
  \e_0_.expander 
  (
    .cinstr_i({ queue_instr_raw_0__15_, queue_instr_raw_0__14_, queue_instr_raw_0__13_, queue_instr_raw_0__12_, queue_instr_raw_0__11_, queue_instr_raw_0__10_, queue_instr_raw_0__9_, queue_instr_raw_0__8_, queue_instr_raw_0__7_, queue_instr_raw_0__6_, queue_instr_raw_0__5_, queue_instr_raw_0__4_, queue_instr_raw_0__3_, queue_instr_raw_0__2_, queue_instr_raw_0__1_, queue_instr_raw_0__0_ }),
    .instr_o(\e_0_.instr )
  );


  bp_be_expander
  \e_1_.expander 
  (
    .cinstr_i({ queue_instr_raw_1__15_, queue_instr_raw_1__14_, queue_instr_raw_1__13_, queue_instr_raw_1__12_, queue_instr_raw_1__11_, queue_instr_raw_1__10_, queue_instr_raw_1__9_, queue_instr_raw_1__8_, queue_instr_raw_1__7_, queue_instr_raw_1__6_, queue_instr_raw_1__5_, queue_instr_raw_1__4_, queue_instr_raw_1__3_, queue_instr_raw_1__2_, queue_instr_raw_1__1_, queue_instr_raw_1__0_ }),
    .instr_o(\e_1_.instr )
  );


  bp_be_expander
  \e_2_.expander 
  (
    .cinstr_i({ queue_instr_raw_2__15_, queue_instr_raw_2__14_, queue_instr_raw_2__13_, queue_instr_raw_2__12_, queue_instr_raw_2__11_, queue_instr_raw_2__10_, queue_instr_raw_2__9_, queue_instr_raw_2__8_, queue_instr_raw_2__7_, queue_instr_raw_2__6_, queue_instr_raw_2__5_, queue_instr_raw_2__4_, queue_instr_raw_2__3_, queue_instr_raw_2__2_, queue_instr_raw_2__1_, queue_instr_raw_2__0_ }),
    .instr_o(\e_2_.instr )
  );


  bp_be_expander
  \e_3_.expander 
  (
    .cinstr_i({ queue_instr_raw_3__15_, queue_instr_raw_3__14_, queue_instr_raw_3__13_, queue_instr_raw_3__12_, queue_instr_raw_3__11_, queue_instr_raw_3__10_, queue_instr_raw_3__9_, queue_instr_raw_3__8_, queue_instr_raw_3__7_, queue_instr_raw_3__6_, queue_instr_raw_3__5_, queue_instr_raw_3__4_, queue_instr_raw_3__3_, queue_instr_raw_3__2_, queue_instr_raw_3__1_, queue_instr_raw_3__0_ }),
    .instr_o(\e_3_.instr )
  );


  bp_be_expander
  \e_4_.expander 
  (
    .cinstr_i({ queue_instr_raw_4__15_, queue_instr_raw_4__14_, queue_instr_raw_4__13_, queue_instr_raw_4__12_, queue_instr_raw_4__11_, queue_instr_raw_4__10_, queue_instr_raw_4__9_, queue_instr_raw_4__8_, queue_instr_raw_4__7_, queue_instr_raw_4__6_, queue_instr_raw_4__5_, queue_instr_raw_4__4_, queue_instr_raw_4__3_, queue_instr_raw_4__2_, queue_instr_raw_4__1_, queue_instr_raw_4__0_ }),
    .instr_o(\e_4_.instr )
  );

  assign N183 = N178 | N179;
  assign N184 = N173 | N174;
  assign N185 = N180 | N181;
  assign N186 = N183 | N184;
  assign N187 = N185 | N182;
  assign N188 = N186 | N187;
  assign N189 = N171 | N172;
  assign N190 = N175 | N181;
  assign N191 = N189 | N184;
  assign N192 = N190 | N182;
  assign N193 = N191 | N192;
  assign N195 = N194 | N174;
  assign N196 = N189 | N195;
  assign N197 = N196 | N192;
  assign N199 = N194 | N198;
  assign N200 = N189 | N199;
  assign N201 = N200 | N192;
  assign N202 = N183 | N195;
  assign N203 = N202 | N192;
  assign N205 = N186 | N192;
  assign N206 = N171 | N179;
  assign N207 = N206 | N184;
  assign N208 = N207 | N192;
  assign N209 = N206 | N195;
  assign N210 = N209 | N192;
  assign N211 = N206 | N199;
  assign N212 = N211 | N192;
  assign N213 = N173 | N198;
  assign N214 = N206 | N213;
  assign N215 = N214 | N187;
  assign N217 = N189 | N213;
  assign N218 = N217 | N187;
  assign N220 = N191 | N187;
  assign N222 = N207 | N187;
  assign N224 = N178 | N172;
  assign N225 = N224 | N195;
  assign N226 = N225 | N192;
  assign N228 = N224 | N184;
  assign N229 = N228 | N192;
  assign N230 = N228 | N187;
  assign N231 = N224 | N213;
  assign N232 = N231 | N192;
  assign N233 = N231 | N187;
  assign N235 = N171 & N172;
  assign N236 = N235 & N174;
  assign N237 = N172 & N194;
  assign N238 = N174 & N180;
  assign N239 = N237 & N238;
  assign N240 = N171 & N173;
  assign N241 = N240 & N174;
  assign N242 = N173 & N175;
  assign N243 = N178 & N194;
  assign N244 = N243 & N238;
  assign N265 = N246 & N247;
  assign N266 = N248 & N249;
  assign N267 = N250 & N251;
  assign N268 = N252 & N253;
  assign N269 = N254 & N255;
  assign N270 = preissue_pkt_o[15] & N256;
  assign N271 = N257 & N258;
  assign N272 = N259 & N260;
  assign N273 = N261 & N262;
  assign N274 = N263 & N264;
  assign N275 = preissue_pkt_o[5] & preissue_pkt_o[4];
  assign N276 = preissue_pkt_o[3] & preissue_pkt_o[2];
  assign N277 = N265 & N266;
  assign N278 = N267 & N268;
  assign N279 = N269 & N270;
  assign N280 = N271 & N272;
  assign N281 = N273 & N274;
  assign N282 = N275 & N276;
  assign N283 = N277 & N278;
  assign N284 = N279 & N280;
  assign N285 = N281 & N282;
  assign N286 = N283 & N284;
  assign N287 = N286 & N285;
  assign N290 = preissue_pkt_o[24] & N288;
  assign N291 = N290 & N289;
  assign N294 = N292 & N293;
  assign N295 = N294 & preissue_pkt_o[22];
  assign N299 = N296 & N297;
  assign N300 = N299 & N298;
  assign N303 = N301 & preissue_pkt_o[23];
  assign N304 = N303 & N302;
  assign N320 = preissue_pkt_o[32] & N312;
  assign N321 = N313 & N314;
  assign N322 = N315 & N316;
  assign N323 = preissue_pkt_o[8] & N317;
  assign N324 = preissue_pkt_o[6] & N318;
  assign N325 = N319 & preissue_pkt_o[3];
  assign N326 = N320 & N321;
  assign N327 = N322 & N323;
  assign N328 = N324 & N325;
  assign N329 = N326 & N327;
  assign N330 = N328 & preissue_pkt_o[2];
  assign N331 = N329 & N330;
  assign N338 = preissue_pkt_o[33] & N333;
  assign N339 = N334 & N335;
  assign N340 = N336 & N337;
  assign N341 = N338 & N339;
  assign N342 = N341 & N340;
  assign N347 = preissue_pkt_o[33] & N343;
  assign N348 = N344 & N345;
  assign N349 = N346 & preissue_pkt_o[22];
  assign N350 = N347 & N348;
  assign N351 = N350 & N349;
  assign N356 = preissue_pkt_o[33] & N352;
  assign N357 = N353 & N354;
  assign N358 = preissue_pkt_o[23] & N355;
  assign N359 = N356 & N357;
  assign N360 = N359 & N358;
  assign N364 = preissue_pkt_o[33] & N361;
  assign N365 = N362 & N363;
  assign N366 = preissue_pkt_o[23] & preissue_pkt_o[22];
  assign N367 = N364 & N365;
  assign N368 = N367 & N366;
  assign N373 = preissue_pkt_o[33] & N369;
  assign N374 = N370 & preissue_pkt_o[27];
  assign N375 = N371 & N372;
  assign N376 = N373 & N374;
  assign N377 = N376 & N375;
  assign N381 = preissue_pkt_o[33] & N378;
  assign N382 = N379 & preissue_pkt_o[27];
  assign N383 = N380 & preissue_pkt_o[22];
  assign N384 = N381 & N382;
  assign N385 = N384 & N383;
  assign N389 = preissue_pkt_o[33] & N386;
  assign N390 = N387 & preissue_pkt_o[27];
  assign N391 = preissue_pkt_o[23] & N388;
  assign N392 = N389 & N390;
  assign N393 = N392 & N391;
  assign N396 = preissue_pkt_o[33] & N394;
  assign N397 = N395 & preissue_pkt_o[27];
  assign N398 = preissue_pkt_o[23] & preissue_pkt_o[22];
  assign N399 = N396 & N397;
  assign N400 = N399 & N398;
  assign N406 = N401 & N402;
  assign N407 = N403 & N404;
  assign N408 = N405 & preissue_pkt_o[22];
  assign N409 = N406 & N407;
  assign N410 = N409 & N408;
  assign N416 = N411 & N412;
  assign N417 = N413 & preissue_pkt_o[27];
  assign N418 = N414 & N415;
  assign N419 = N416 & N417;
  assign N420 = N419 & N418;
  assign N428 = preissue_pkt_o[33] & preissue_pkt_o[31];
  assign N429 = N421 & N422;
  assign N430 = N423 & N424;
  assign N431 = N425 & N426;
  assign N432 = N428 & N429;
  assign N433 = N430 & N431;
  assign N434 = N432 & N433;
  assign N435 = N434 & N427;
  assign N442 = preissue_pkt_o[33] & preissue_pkt_o[31];
  assign N443 = N436 & preissue_pkt_o[27];
  assign N444 = N437 & N438;
  assign N445 = N439 & N440;
  assign N446 = N442 & N443;
  assign N447 = N444 & N445;
  assign N448 = N446 & N447;
  assign N449 = N448 & N441;
  assign N456 = preissue_pkt_o[33] & preissue_pkt_o[31];
  assign N457 = N450 & N451;
  assign N458 = N452 & N453;
  assign N459 = N454 & N455;
  assign N460 = N456 & N457;
  assign N461 = N458 & N459;
  assign N462 = N460 & N461;
  assign N463 = N462 & preissue_pkt_o[14];
  assign N469 = preissue_pkt_o[33] & preissue_pkt_o[31];
  assign N470 = N464 & preissue_pkt_o[27];
  assign N471 = N465 & N466;
  assign N472 = N467 & N468;
  assign N473 = N469 & N470;
  assign N474 = N471 & N472;
  assign N475 = N473 & N474;
  assign N476 = N475 & preissue_pkt_o[14];
  assign N482 = preissue_pkt_o[33] & N478;
  assign N483 = preissue_pkt_o[30] & N479;
  assign N484 = N480 & N481;
  assign N485 = N482 & N483;
  assign N486 = N485 & N484;
  assign N490 = preissue_pkt_o[33] & N487;
  assign N491 = preissue_pkt_o[30] & N488;
  assign N492 = N489 & preissue_pkt_o[22];
  assign N493 = N490 & N491;
  assign N494 = N493 & N492;
  assign N498 = preissue_pkt_o[33] & N495;
  assign N499 = preissue_pkt_o[30] & N496;
  assign N500 = preissue_pkt_o[23] & N497;
  assign N501 = N498 & N499;
  assign N502 = N501 & N500;
  assign N505 = preissue_pkt_o[33] & N503;
  assign N506 = preissue_pkt_o[30] & N504;
  assign N507 = preissue_pkt_o[23] & preissue_pkt_o[22];
  assign N508 = N505 & N506;
  assign N509 = N508 & N507;
  assign N513 = preissue_pkt_o[33] & N510;
  assign N514 = preissue_pkt_o[30] & preissue_pkt_o[27];
  assign N515 = N511 & N512;
  assign N516 = N513 & N514;
  assign N517 = N516 & N515;
  assign N520 = preissue_pkt_o[33] & N518;
  assign N521 = preissue_pkt_o[30] & preissue_pkt_o[27];
  assign N522 = N519 & preissue_pkt_o[22];
  assign N523 = N520 & N521;
  assign N524 = N523 & N522;
  assign N527 = preissue_pkt_o[33] & N525;
  assign N528 = preissue_pkt_o[30] & preissue_pkt_o[27];
  assign N529 = preissue_pkt_o[23] & N526;
  assign N530 = N527 & N528;
  assign N531 = N530 & N529;
  assign N533 = preissue_pkt_o[33] & N532;
  assign N534 = preissue_pkt_o[30] & preissue_pkt_o[27];
  assign N535 = preissue_pkt_o[23] & preissue_pkt_o[22];
  assign N536 = N533 & N534;
  assign N537 = N536 & N535;
  assign N544 = preissue_pkt_o[33] & preissue_pkt_o[31];
  assign N545 = preissue_pkt_o[30] & N538;
  assign N546 = N539 & N540;
  assign N547 = N541 & N542;
  assign N548 = N544 & N545;
  assign N549 = N546 & N547;
  assign N550 = N548 & N549;
  assign N551 = N550 & N543;
  assign N557 = preissue_pkt_o[33] & preissue_pkt_o[31];
  assign N558 = preissue_pkt_o[30] & preissue_pkt_o[27];
  assign N559 = N552 & N553;
  assign N560 = N554 & N555;
  assign N561 = N557 & N558;
  assign N562 = N559 & N560;
  assign N563 = N561 & N562;
  assign N564 = N563 & N556;
  assign N567 = N566 & preissue_pkt_o[27];
  assign N568 = N567 & preissue_pkt_o[22];
  assign N570 = N569 & preissue_pkt_o[31];
  assign N571 = N570 & preissue_pkt_o[27];
  assign N572 = preissue_pkt_o[31] & preissue_pkt_o[22];
  assign N574 = N573 & preissue_pkt_o[23];
  assign N576 = N575 & preissue_pkt_o[30];
  assign N580 = N577 & N578;
  assign N581 = N580 & N579;
  assign N582 = preissue_pkt_o[31] & preissue_pkt_o[30];
  assign N583 = N582 & preissue_pkt_o[14];
  assign N584 = preissue_pkt_o[31] & preissue_pkt_o[23];
  assign N585 = preissue_pkt_o[31] & preissue_pkt_o[16];
  assign N586 = preissue_pkt_o[31] & preissue_pkt_o[15];

  bsg_dff_reset_en_width_p39
  issue_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(preissue_v),
    .data_i(preissue_pkt_o),
    .data_o({ preissue_pkt_r_irs1_v_, preissue_pkt_r_irs2_v_, preissue_pkt_r_frs1_v_, preissue_pkt_r_frs2_v_, preissue_pkt_r_frs3_v_, issue_pkt_o[205:174], preissue_pkt_r_size__1_, preissue_pkt_r_size__0_ })
  );

  assign bypass_issue = wptr_r[5:3] == rptr_r[5:3];

  bsg_mem_1r1w_000000ae_00000008
  queue_fifo_mem
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(_4_net_),
    .w_addr_i(wptr_r[5:3]),
    .w_data_i(fe_queue_i),
    .r_v_i(_6_net_),
    .r_addr_i(rptr_r[5:3]),
    .r_data_o({ fe_queue_lo_pc__38_, fe_queue_lo_pc__37_, fe_queue_lo_pc__36_, fe_queue_lo_pc__35_, fe_queue_lo_pc__34_, fe_queue_lo_pc__33_, fe_queue_lo_pc__32_, fe_queue_lo_pc__31_, fe_queue_lo_pc__30_, fe_queue_lo_pc__29_, fe_queue_lo_pc__28_, fe_queue_lo_pc__27_, fe_queue_lo_pc__26_, fe_queue_lo_pc__25_, fe_queue_lo_pc__24_, fe_queue_lo_pc__23_, fe_queue_lo_pc__22_, fe_queue_lo_pc__21_, fe_queue_lo_pc__20_, fe_queue_lo_pc__19_, fe_queue_lo_pc__18_, fe_queue_lo_pc__17_, fe_queue_lo_pc__16_, fe_queue_lo_pc__15_, fe_queue_lo_pc__14_, fe_queue_lo_pc__13_, fe_queue_lo_pc__12_, fe_queue_lo_pc__11_, fe_queue_lo_pc__10_, fe_queue_lo_pc__9_, fe_queue_lo_pc__8_, fe_queue_lo_pc__7_, fe_queue_lo_pc__6_, fe_queue_lo_pc__5_, fe_queue_lo_pc__4_, fe_queue_lo_pc__3_, fe_queue_lo_pc__2_, fe_queue_lo_pc__1_, fe_queue_lo_pc__0_, fe_queue_lo_instr__79_, fe_queue_lo_instr__78_, fe_queue_lo_instr__77_, fe_queue_lo_instr__76_, fe_queue_lo_instr__75_, fe_queue_lo_instr__74_, fe_queue_lo_instr__73_, fe_queue_lo_instr__72_, fe_queue_lo_instr__71_, fe_queue_lo_instr__70_, fe_queue_lo_instr__69_, fe_queue_lo_instr__68_, fe_queue_lo_instr__67_, fe_queue_lo_instr__66_, fe_queue_lo_instr__65_, fe_queue_lo_instr__64_, fe_queue_lo_instr__63_, fe_queue_lo_instr__62_, fe_queue_lo_instr__61_, fe_queue_lo_instr__60_, fe_queue_lo_instr__59_, fe_queue_lo_instr__58_, fe_queue_lo_instr__57_, fe_queue_lo_instr__56_, fe_queue_lo_instr__55_, fe_queue_lo_instr__54_, fe_queue_lo_instr__53_, fe_queue_lo_instr__52_, fe_queue_lo_instr__51_, fe_queue_lo_instr__50_, fe_queue_lo_instr__49_, fe_queue_lo_instr__48_, fe_queue_lo_instr__47_, fe_queue_lo_instr__46_, fe_queue_lo_instr__45_, fe_queue_lo_instr__44_, fe_queue_lo_instr__43_, fe_queue_lo_instr__42_, fe_queue_lo_instr__41_, fe_queue_lo_instr__40_, fe_queue_lo_instr__39_, fe_queue_lo_instr__38_, fe_queue_lo_instr__37_, fe_queue_lo_instr__36_, fe_queue_lo_instr__35_, fe_queue_lo_instr__34_, fe_queue_lo_instr__33_, fe_queue_lo_instr__32_, fe_queue_lo_instr__31_, fe_queue_lo_instr__30_, fe_queue_lo_instr__29_, fe_queue_lo_instr__28_, fe_queue_lo_instr__27_, fe_queue_lo_instr__26_, fe_queue_lo_instr__25_, fe_queue_lo_instr__24_, fe_queue_lo_instr__23_, fe_queue_lo_instr__22_, fe_queue_lo_instr__21_, fe_queue_lo_instr__20_, fe_queue_lo_instr__19_, fe_queue_lo_instr__18_, fe_queue_lo_instr__17_, fe_queue_lo_instr__16_, fe_queue_lo_instr__15_, fe_queue_lo_instr__14_, fe_queue_lo_instr__13_, fe_queue_lo_instr__12_, fe_queue_lo_instr__11_, fe_queue_lo_instr__10_, fe_queue_lo_instr__9_, fe_queue_lo_instr__8_, fe_queue_lo_instr__7_, fe_queue_lo_instr__6_, fe_queue_lo_instr__5_, fe_queue_lo_instr__4_, fe_queue_lo_instr__3_, fe_queue_lo_instr__2_, fe_queue_lo_instr__1_, fe_queue_lo_instr__0_, issue_pkt_o[48:0], issue_pkt_o[173:171], fe_queue_lo_msg_type__2_, fe_queue_lo_msg_type__1_, fe_queue_lo_msg_type__0_ })
  );


  bp_be_instr_decoder_00
  instr_decoder
  (
    .preissue_pkt_i({ preissue_pkt_r_irs1_v_, preissue_pkt_r_irs2_v_, preissue_pkt_r_frs1_v_, preissue_pkt_r_frs2_v_, preissue_pkt_r_frs3_v_, issue_pkt_o[205:174], preissue_pkt_r_size__1_, preissue_pkt_r_size__0_ }),
    .decode_info_i(decode_info_i),
    .decode_o(issue_pkt_o[168:115]),
    .illegal_instr_o(illegal_instr_lo),
    .ecall_m_o(issue_pkt_o[256]),
    .ecall_s_o(issue_pkt_o[255]),
    .ecall_u_o(issue_pkt_o[254]),
    .ebreak_o(issue_pkt_o[253]),
    .dbreak_o(issue_pkt_o[252]),
    .dret_o(issue_pkt_o[251]),
    .mret_o(issue_pkt_o[250]),
    .sret_o(issue_pkt_o[249]),
    .wfi_o(issue_pkt_o[248]),
    .sfence_vma_o(issue_pkt_o[247]),
    .fencei_o(issue_pkt_o[246]),
    .csrw_o(issue_pkt_o[245]),
    .imm_o(issue_pkt_o[112:49])
  );

  assign N601 = fe_queue_lo_msg_type__1_ | fe_queue_lo_msg_type__2_;
  assign N602 = fe_queue_lo_msg_type__0_ | N601;
  assign issue_pkt_o[261] = ~N602;
  assign N604 = ~fe_queue_lo_msg_type__1_;
  assign N605 = N604 | fe_queue_lo_msg_type__2_;
  assign N606 = fe_queue_lo_msg_type__0_ | N605;
  assign issue_pkt_o[260] = ~N606;
  assign N608 = ~fe_queue_lo_msg_type__0_;
  assign N609 = fe_queue_lo_msg_type__1_ | fe_queue_lo_msg_type__2_;
  assign N610 = N608 | N609;
  assign issue_pkt_o[259] = ~N610;
  assign N612 = N604 | fe_queue_lo_msg_type__2_;
  assign N613 = N608 | N612;
  assign issue_pkt_o[258] = ~N613;
  assign N615 = ~fe_queue_lo_msg_type__2_;
  assign N616 = fe_queue_lo_msg_type__1_ | N615;
  assign N617 = fe_queue_lo_msg_type__0_ | N616;
  assign N618 = ~N617;
  assign N619 = fe_queue_lo_msg_type__1_ | N615;
  assign N620 = fe_queue_lo_msg_type__0_ | N619;
  assign N621 = ~N620;
  assign N622 = ~preissue_size_0__0_;
  assign N623 = N622 | preissue_size_0__1_;
  assign N624 = ~N623;
  assign N625 = ~preissue_size_1__0_;
  assign N626 = N625 | preissue_size_1__1_;
  assign N627 = ~N626;
  assign N628 = ~preissue_size_2__0_;
  assign N629 = N628 | preissue_size_2__1_;
  assign N630 = ~N629;
  assign N631 = ~preissue_size_3__0_;
  assign N632 = N631 | preissue_size_3__1_;
  assign N633 = ~N632;
  assign N634 = ~preissue_size_4__0_;
  assign N635 = N634 | preissue_size_4__1_;
  assign N636 = ~N635;
  assign { N78, N77, N76, N75 } = cptr_r[2:0] + cmt_size_i;
  assign { N74, N73, N72, N71 } = rptr_r[2:0] + read_size_i;
  assign issue_pkt_o[244:206] = { fe_queue_lo_pc__38_, fe_queue_lo_pc__37_, fe_queue_lo_pc__36_, fe_queue_lo_pc__35_, fe_queue_lo_pc__34_, fe_queue_lo_pc__33_, fe_queue_lo_pc__32_, fe_queue_lo_pc__31_, fe_queue_lo_pc__30_, fe_queue_lo_pc__29_, fe_queue_lo_pc__28_, fe_queue_lo_pc__27_, fe_queue_lo_pc__26_, fe_queue_lo_pc__25_, fe_queue_lo_pc__24_, fe_queue_lo_pc__23_, fe_queue_lo_pc__22_, fe_queue_lo_pc__21_, fe_queue_lo_pc__20_, fe_queue_lo_pc__19_, fe_queue_lo_pc__18_, fe_queue_lo_pc__17_, fe_queue_lo_pc__16_, fe_queue_lo_pc__15_, fe_queue_lo_pc__14_, fe_queue_lo_pc__13_, fe_queue_lo_pc__12_, fe_queue_lo_pc__11_, fe_queue_lo_pc__10_, fe_queue_lo_pc__9_, fe_queue_lo_pc__8_, fe_queue_lo_pc__7_, fe_queue_lo_pc__6_, fe_queue_lo_pc__5_, fe_queue_lo_pc__4_, fe_queue_lo_pc__3_, fe_queue_lo_pc__2_, fe_queue_lo_pc__1_, fe_queue_lo_pc__0_ } + { rptr_r[2:0], 1'b0 };
  assign { N152, N151, N150, N149, N148, N147, N146 } = 1'b0 - cptr_r;
  assign { N145, N144, N143, N142, N141, N140, N139 } = 1'b0 - wptr_r;
  assign { N120, N119, N118, N117, N116, N115, N114 } = 1'b0 - rptr_r;
  assign { N107, N106, N105, N104 } = { 1'b1, 1'b0, 1'b0, 1'b0 } - cptr_r[2:0];
  assign { N96, N95, N94, N93 } = { 1'b1, 1'b0, 1'b0, 1'b0 } - rptr_r[2:0];
  assign { N128, N127, N126, N125, N124, N123, N122 } = cptr_r - rptr_r;
  assign { N135, N134, N133, N132, N131, N130, N129 } = { N128, N127, N126, N125, N124, N123, N122 } + deq;
  assign { N85, N84, N83, N82 } = { 1'b1, 1'b0, 1'b0, 1'b0 } - wptr_r[2:0];
  assign N159 = N0 & N1 & N2;
  assign N0 = ~preissue_entry_sel[2];
  assign N1 = ~preissue_entry_sel[0];
  assign N2 = ~preissue_entry_sel[1];
  assign N160 = preissue_entry_sel[0] & N3;
  assign N3 = ~preissue_entry_sel[1];
  assign N161 = N4 & preissue_entry_sel[1];
  assign N4 = ~preissue_entry_sel[0];
  assign N162 = preissue_entry_sel[0] & preissue_entry_sel[1];
  assign N163 = N5 & N6 & N7;
  assign N5 = ~preissue_entry_sel[2];
  assign N6 = ~preissue_entry_sel[0];
  assign N7 = ~preissue_entry_sel[1];
  assign N164 = preissue_entry_sel[0] & N8;
  assign N8 = ~preissue_entry_sel[1];
  assign N165 = N9 & preissue_entry_sel[1];
  assign N9 = ~preissue_entry_sel[0];
  assign N166 = preissue_entry_sel[0] & preissue_entry_sel[1];
  assign N167 = N10 & N11 & N12;
  assign N10 = ~preissue_entry_sel[2];
  assign N11 = ~preissue_entry_sel[0];
  assign N12 = ~preissue_entry_sel[1];
  assign N168 = preissue_entry_sel[0] & N13;
  assign N13 = ~preissue_entry_sel[1];
  assign N169 = N14 & preissue_entry_sel[1];
  assign N14 = ~preissue_entry_sel[0];
  assign N170 = preissue_entry_sel[0] & preissue_entry_sel[1];
  assign { N89, N88, N87, N86 } = (N15)? { N85, N84, N83, N82 } : 
                                  (N16)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = 1'b1;
  assign N16 = N81;
  assign enq = (N17)? { N89, N88, N87, N86 } : 
               (N18)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N17 = ack;
  assign N18 = N79;
  assign { N100, N99, N98, N97 } = (N19)? { N96, N95, N94, N93 } : 
                                   (N20)? read_size_i : 1'b0;
  assign N19 = read_catchup;
  assign N20 = N92;
  assign read = (N21)? { N100, N99, N98, N97 } : 
                (N22)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N21 = read_i;
  assign N22 = N90;
  assign { N111, N110, N109, N108 } = (N23)? { N107, N106, N105, N104 } : 
                                      (N24)? cmt_size_i : 1'b0;
  assign N23 = deq_catchup;
  assign N24 = N103;
  assign deq = (N25)? { N111, N110, N109, N108 } : 
               (N26)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N25 = cmt_i;
  assign N26 = N101;
  assign rptr_jmp = (N27)? { N120, N119, N118, N117, N116, N115, N114 } : 
                    (N137)? { N135, N134, N133, N132, N131, N130, N129 } : 
                    (N113)? { 1'b0, 1'b0, 1'b0, read } : 1'b0;
  assign N27 = clr_i;
  assign wptr_jmp = (N27)? { N145, N144, N143, N142, N141, N140, N139 } : 
                    (N28)? { 1'b0, 1'b0, 1'b0, enq } : 1'b0;
  assign N28 = N138;
  assign cptr_jmp = (N27)? { N152, N151, N150, N149, N148, N147, N146 } : 
                    (N28)? { 1'b0, 1'b0, 1'b0, deq } : 1'b0;
  assign preissue_entry_sel = (N29)? wptr_r[2:0] : 
                              (N30)? rptr_n[2:0] : 1'b0;
  assign N29 = bypass_preissue;
  assign N30 = N153;
  assign { queue_instr_raw_4__15_, queue_instr_raw_4__14_, queue_instr_raw_4__13_, queue_instr_raw_4__12_, queue_instr_raw_4__11_, queue_instr_raw_4__10_, queue_instr_raw_4__9_, queue_instr_raw_4__8_, queue_instr_raw_4__7_, queue_instr_raw_4__6_, queue_instr_raw_4__5_, queue_instr_raw_4__4_, queue_instr_raw_4__3_, queue_instr_raw_4__2_, queue_instr_raw_4__1_, queue_instr_raw_4__0_, queue_instr_raw_3__15_, queue_instr_raw_3__14_, queue_instr_raw_3__13_, queue_instr_raw_3__12_, queue_instr_raw_3__11_, queue_instr_raw_3__10_, queue_instr_raw_3__9_, queue_instr_raw_3__8_, queue_instr_raw_3__7_, queue_instr_raw_3__6_, queue_instr_raw_3__5_, queue_instr_raw_3__4_, queue_instr_raw_3__3_, queue_instr_raw_3__2_, queue_instr_raw_3__1_, queue_instr_raw_3__0_, queue_instr_raw_2__15_, queue_instr_raw_2__14_, queue_instr_raw_2__13_, queue_instr_raw_2__12_, queue_instr_raw_2__11_, queue_instr_raw_2__10_, queue_instr_raw_2__9_, queue_instr_raw_2__8_, queue_instr_raw_2__7_, queue_instr_raw_2__6_, queue_instr_raw_2__5_, queue_instr_raw_2__4_, queue_instr_raw_2__3_, queue_instr_raw_2__2_, queue_instr_raw_2__1_, queue_instr_raw_2__0_, queue_instr_raw_1__15_, queue_instr_raw_1__14_, queue_instr_raw_1__13_, queue_instr_raw_1__12_, queue_instr_raw_1__11_, queue_instr_raw_1__10_, queue_instr_raw_1__9_, queue_instr_raw_1__8_, queue_instr_raw_1__7_, queue_instr_raw_1__6_, queue_instr_raw_1__5_, queue_instr_raw_1__4_, queue_instr_raw_1__3_, queue_instr_raw_1__2_, queue_instr_raw_1__1_, queue_instr_raw_1__0_, queue_instr_raw_0__15_, queue_instr_raw_0__14_, queue_instr_raw_0__13_, queue_instr_raw_0__12_, queue_instr_raw_0__11_, queue_instr_raw_0__10_, queue_instr_raw_0__9_, queue_instr_raw_0__8_, queue_instr_raw_0__7_, queue_instr_raw_0__6_, queue_instr_raw_0__5_, queue_instr_raw_0__4_, queue_instr_raw_0__3_, queue_instr_raw_0__2_, queue_instr_raw_0__1_, queue_instr_raw_0__0_ } = (N29)? fe_queue_i[134:55] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (N30)? queue_instr_n : 1'b0;
  assign preissue_size_0__1_ = ~preissue_size_0__0_;
  assign preissue_instr[31:0] = (N31)? \e_0_.instr  : 
                                (N32)? { queue_instr_raw_1__15_, queue_instr_raw_1__14_, queue_instr_raw_1__13_, queue_instr_raw_1__12_, queue_instr_raw_1__11_, queue_instr_raw_1__10_, queue_instr_raw_1__9_, queue_instr_raw_1__8_, queue_instr_raw_1__7_, queue_instr_raw_1__6_, queue_instr_raw_1__5_, queue_instr_raw_1__4_, queue_instr_raw_1__3_, queue_instr_raw_1__2_, queue_instr_raw_1__1_, queue_instr_raw_1__0_, queue_instr_raw_0__15_, queue_instr_raw_0__14_, queue_instr_raw_0__13_, queue_instr_raw_0__12_, queue_instr_raw_0__11_, queue_instr_raw_0__10_, queue_instr_raw_0__9_, queue_instr_raw_0__8_, queue_instr_raw_0__7_, queue_instr_raw_0__6_, queue_instr_raw_0__5_, queue_instr_raw_0__4_, queue_instr_raw_0__3_, queue_instr_raw_0__2_, queue_instr_raw_0__1_, queue_instr_raw_0__0_ } : 1'b0;
  assign N31 = N624;
  assign N32 = N623;
  assign preissue_size_1__1_ = ~preissue_size_1__0_;
  assign preissue_instr[63:32] = (N33)? \e_1_.instr  : 
                                 (N34)? { queue_instr_raw_2__15_, queue_instr_raw_2__14_, queue_instr_raw_2__13_, queue_instr_raw_2__12_, queue_instr_raw_2__11_, queue_instr_raw_2__10_, queue_instr_raw_2__9_, queue_instr_raw_2__8_, queue_instr_raw_2__7_, queue_instr_raw_2__6_, queue_instr_raw_2__5_, queue_instr_raw_2__4_, queue_instr_raw_2__3_, queue_instr_raw_2__2_, queue_instr_raw_2__1_, queue_instr_raw_2__0_, queue_instr_raw_1__15_, queue_instr_raw_1__14_, queue_instr_raw_1__13_, queue_instr_raw_1__12_, queue_instr_raw_1__11_, queue_instr_raw_1__10_, queue_instr_raw_1__9_, queue_instr_raw_1__8_, queue_instr_raw_1__7_, queue_instr_raw_1__6_, queue_instr_raw_1__5_, queue_instr_raw_1__4_, queue_instr_raw_1__3_, queue_instr_raw_1__2_, queue_instr_raw_1__1_, queue_instr_raw_1__0_ } : 1'b0;
  assign N33 = N627;
  assign N34 = N626;
  assign preissue_size_2__1_ = ~preissue_size_2__0_;
  assign preissue_instr[95:64] = (N35)? \e_2_.instr  : 
                                 (N36)? { queue_instr_raw_3__15_, queue_instr_raw_3__14_, queue_instr_raw_3__13_, queue_instr_raw_3__12_, queue_instr_raw_3__11_, queue_instr_raw_3__10_, queue_instr_raw_3__9_, queue_instr_raw_3__8_, queue_instr_raw_3__7_, queue_instr_raw_3__6_, queue_instr_raw_3__5_, queue_instr_raw_3__4_, queue_instr_raw_3__3_, queue_instr_raw_3__2_, queue_instr_raw_3__1_, queue_instr_raw_3__0_, queue_instr_raw_2__15_, queue_instr_raw_2__14_, queue_instr_raw_2__13_, queue_instr_raw_2__12_, queue_instr_raw_2__11_, queue_instr_raw_2__10_, queue_instr_raw_2__9_, queue_instr_raw_2__8_, queue_instr_raw_2__7_, queue_instr_raw_2__6_, queue_instr_raw_2__5_, queue_instr_raw_2__4_, queue_instr_raw_2__3_, queue_instr_raw_2__2_, queue_instr_raw_2__1_, queue_instr_raw_2__0_ } : 1'b0;
  assign N35 = N630;
  assign N36 = N629;
  assign preissue_size_3__1_ = ~preissue_size_3__0_;
  assign preissue_instr[127:96] = (N37)? \e_3_.instr  : 
                                  (N38)? { queue_instr_raw_4__15_, queue_instr_raw_4__14_, queue_instr_raw_4__13_, queue_instr_raw_4__12_, queue_instr_raw_4__11_, queue_instr_raw_4__10_, queue_instr_raw_4__9_, queue_instr_raw_4__8_, queue_instr_raw_4__7_, queue_instr_raw_4__6_, queue_instr_raw_4__5_, queue_instr_raw_4__4_, queue_instr_raw_4__3_, queue_instr_raw_4__2_, queue_instr_raw_4__1_, queue_instr_raw_4__0_, queue_instr_raw_3__15_, queue_instr_raw_3__14_, queue_instr_raw_3__13_, queue_instr_raw_3__12_, queue_instr_raw_3__11_, queue_instr_raw_3__10_, queue_instr_raw_3__9_, queue_instr_raw_3__8_, queue_instr_raw_3__7_, queue_instr_raw_3__6_, queue_instr_raw_3__5_, queue_instr_raw_3__4_, queue_instr_raw_3__3_, queue_instr_raw_3__2_, queue_instr_raw_3__1_, queue_instr_raw_3__0_ } : 1'b0;
  assign N37 = N633;
  assign N38 = N632;
  assign preissue_size_4__1_ = ~preissue_size_4__0_;
  assign preissue_instr[159:128] = (N39)? \e_4_.instr  : 
                                   (N40)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, queue_instr_raw_4__15_, queue_instr_raw_4__14_, queue_instr_raw_4__13_, queue_instr_raw_4__12_, queue_instr_raw_4__11_, queue_instr_raw_4__10_, queue_instr_raw_4__9_, queue_instr_raw_4__8_, queue_instr_raw_4__7_, queue_instr_raw_4__6_, queue_instr_raw_4__5_, queue_instr_raw_4__4_, queue_instr_raw_4__3_, queue_instr_raw_4__2_, queue_instr_raw_4__1_, queue_instr_raw_4__0_ } : 1'b0;
  assign N39 = N636;
  assign N40 = N635;
  assign { N308, N307 } = (N41)? { preissue_v, preissue_v } : 
                          (N306)? { 1'b0, 1'b0 } : 1'b0;
  assign N41 = N305;
  assign { N311, N310 } = (N42)? { N308, N307 } : 
                          (N309)? { 1'b0, 1'b0 } : 1'b0;
  assign N42 = N287;
  assign N590 = (N43)? preissue_v : 
                (N589)? 1'b0 : 1'b0;
  assign N43 = N587;
  assign N591 = (N44)? preissue_v : 
                (N45)? 1'b0 : 
                (N43)? preissue_v : 1'b0;
  assign N44 = N477;
  assign N45 = N565;
  assign N594 = (N45)? preissue_v : 
                (N593)? 1'b0 : 1'b0;
  assign { N597, N596, N595 } = (N46)? { N594, N591, N590 } : 
                                (N332)? { 1'b0, preissue_v, preissue_v } : 1'b0;
  assign N46 = N331;
  assign preissue_pkt_o[34] = (N47)? preissue_v : 
                              (N599)? 1'b0 : 1'b0;
  assign N47 = N234;
  assign preissue_pkt_o[38:35] = (N48)? { preissue_v, 1'b0, 1'b0, 1'b0 } : 
                                 (N49)? { preissue_v, preissue_v, 1'b0, 1'b0 } : 
                                 (N50)? { N311, N310, 1'b0, 1'b0 } : 
                                 (N51)? { preissue_v, 1'b0, 1'b0, 1'b0 } : 
                                 (N52)? { preissue_v, 1'b0, 1'b0, preissue_v } : 
                                 (N53)? { N597, 1'b0, N596, N595 } : 
                                 (N47)? { 1'b0, 1'b0, preissue_v, preissue_v } : 
                                 (N54)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N48 = N204;
  assign N49 = N216;
  assign N50 = N219;
  assign N51 = N221;
  assign N52 = N223;
  assign N53 = N227;
  assign N54 = N245;
  assign issue_pkt_o[170:169] = (N55)? { preissue_pkt_r_size__1_, preissue_pkt_r_size__0_ } : 
                                (N600)? { 1'b1, 1'b1 } : 1'b0;
  assign N55 = issue_pkt_o[262];
  assign preissue_pkt_o[0] = (N56)? preissue_size_0__0_ : 
                             (N57)? preissue_size_1__0_ : 
                             (N58)? preissue_size_2__0_ : 
                             (N59)? preissue_size_3__0_ : 
                             (N60)? preissue_size_4__0_ : 1'b0;
  assign N56 = N159;
  assign N57 = N160;
  assign N58 = N161;
  assign N59 = N162;
  assign N60 = preissue_entry_sel[2];
  assign preissue_pkt_o[1] = (N56)? preissue_size_0__1_ : 
                             (N57)? preissue_size_1__1_ : 
                             (N58)? preissue_size_2__1_ : 
                             (N59)? preissue_size_3__1_ : 
                             (N60)? preissue_size_4__1_ : 1'b0;
  assign preissue_pkt_o[2] = (N61)? preissue_instr[0] : 
                             (N62)? preissue_instr[32] : 
                             (N63)? preissue_instr[64] : 
                             (N64)? preissue_instr[96] : 
                             (N60)? preissue_instr[128] : 1'b0;
  assign N61 = N163;
  assign N62 = N164;
  assign N63 = N165;
  assign N64 = N166;
  assign N177 = (N65)? preissue_instr[0] : 
                (N66)? preissue_instr[32] : 
                (N67)? preissue_instr[64] : 
                (N68)? preissue_instr[96] : 
                (N60)? preissue_instr[128] : 1'b0;
  assign N65 = N167;
  assign N66 = N168;
  assign N67 = N169;
  assign N68 = N170;
  assign preissue_pkt_o[3] = (N61)? preissue_instr[1] : 
                             (N62)? preissue_instr[33] : 
                             (N63)? preissue_instr[65] : 
                             (N64)? preissue_instr[97] : 
                             (N60)? preissue_instr[129] : 1'b0;
  assign N176 = (N65)? preissue_instr[1] : 
                (N66)? preissue_instr[33] : 
                (N67)? preissue_instr[65] : 
                (N68)? preissue_instr[97] : 
                (N60)? preissue_instr[129] : 1'b0;
  assign preissue_pkt_o[4] = (N61)? preissue_instr[2] : 
                             (N62)? preissue_instr[34] : 
                             (N63)? preissue_instr[66] : 
                             (N64)? preissue_instr[98] : 
                             (N60)? preissue_instr[130] : 1'b0;
  assign N175 = (N65)? preissue_instr[2] : 
                (N66)? preissue_instr[34] : 
                (N67)? preissue_instr[66] : 
                (N68)? preissue_instr[98] : 
                (N60)? preissue_instr[130] : 1'b0;
  assign preissue_pkt_o[5] = (N61)? preissue_instr[3] : 
                             (N62)? preissue_instr[35] : 
                             (N63)? preissue_instr[67] : 
                             (N64)? preissue_instr[99] : 
                             (N60)? preissue_instr[131] : 1'b0;
  assign N174 = (N65)? preissue_instr[3] : 
                (N66)? preissue_instr[35] : 
                (N67)? preissue_instr[67] : 
                (N68)? preissue_instr[99] : 
                (N60)? preissue_instr[131] : 1'b0;
  assign preissue_pkt_o[6] = (N61)? preissue_instr[4] : 
                             (N62)? preissue_instr[36] : 
                             (N63)? preissue_instr[68] : 
                             (N64)? preissue_instr[100] : 
                             (N60)? preissue_instr[132] : 1'b0;
  assign N173 = (N65)? preissue_instr[4] : 
                (N66)? preissue_instr[36] : 
                (N67)? preissue_instr[68] : 
                (N68)? preissue_instr[100] : 
                (N60)? preissue_instr[132] : 1'b0;
  assign preissue_pkt_o[7] = (N61)? preissue_instr[5] : 
                             (N62)? preissue_instr[37] : 
                             (N63)? preissue_instr[69] : 
                             (N64)? preissue_instr[101] : 
                             (N60)? preissue_instr[133] : 1'b0;
  assign N172 = (N65)? preissue_instr[5] : 
                (N66)? preissue_instr[37] : 
                (N67)? preissue_instr[69] : 
                (N68)? preissue_instr[101] : 
                (N60)? preissue_instr[133] : 1'b0;
  assign preissue_pkt_o[8] = (N61)? preissue_instr[6] : 
                             (N62)? preissue_instr[38] : 
                             (N63)? preissue_instr[70] : 
                             (N64)? preissue_instr[102] : 
                             (N60)? preissue_instr[134] : 1'b0;
  assign N171 = (N65)? preissue_instr[6] : 
                (N66)? preissue_instr[38] : 
                (N67)? preissue_instr[70] : 
                (N68)? preissue_instr[102] : 
                (N60)? preissue_instr[134] : 1'b0;
  assign preissue_pkt_o[9] = (N61)? preissue_instr[7] : 
                             (N62)? preissue_instr[39] : 
                             (N63)? preissue_instr[71] : 
                             (N64)? preissue_instr[103] : 
                             (N60)? preissue_instr[135] : 1'b0;
  assign preissue_pkt_o[10] = (N61)? preissue_instr[8] : 
                              (N62)? preissue_instr[40] : 
                              (N63)? preissue_instr[72] : 
                              (N64)? preissue_instr[104] : 
                              (N60)? preissue_instr[136] : 1'b0;
  assign preissue_pkt_o[11] = (N61)? preissue_instr[9] : 
                              (N62)? preissue_instr[41] : 
                              (N63)? preissue_instr[73] : 
                              (N64)? preissue_instr[105] : 
                              (N60)? preissue_instr[137] : 1'b0;
  assign preissue_pkt_o[12] = (N61)? preissue_instr[10] : 
                              (N62)? preissue_instr[42] : 
                              (N63)? preissue_instr[74] : 
                              (N64)? preissue_instr[106] : 
                              (N60)? preissue_instr[138] : 1'b0;
  assign preissue_pkt_o[13] = (N61)? preissue_instr[11] : 
                              (N62)? preissue_instr[43] : 
                              (N63)? preissue_instr[75] : 
                              (N64)? preissue_instr[107] : 
                              (N60)? preissue_instr[139] : 1'b0;
  assign preissue_pkt_o[14] = (N61)? preissue_instr[12] : 
                              (N62)? preissue_instr[44] : 
                              (N63)? preissue_instr[76] : 
                              (N64)? preissue_instr[108] : 
                              (N60)? preissue_instr[140] : 1'b0;
  assign preissue_pkt_o[15] = (N61)? preissue_instr[13] : 
                              (N62)? preissue_instr[45] : 
                              (N63)? preissue_instr[77] : 
                              (N64)? preissue_instr[109] : 
                              (N60)? preissue_instr[141] : 1'b0;
  assign preissue_pkt_o[16] = (N61)? preissue_instr[14] : 
                              (N62)? preissue_instr[46] : 
                              (N63)? preissue_instr[78] : 
                              (N64)? preissue_instr[110] : 
                              (N60)? preissue_instr[142] : 1'b0;
  assign preissue_pkt_o[17] = (N61)? preissue_instr[15] : 
                              (N62)? preissue_instr[47] : 
                              (N63)? preissue_instr[79] : 
                              (N64)? preissue_instr[111] : 
                              (N60)? preissue_instr[143] : 1'b0;
  assign preissue_pkt_o[18] = (N61)? preissue_instr[16] : 
                              (N62)? preissue_instr[48] : 
                              (N63)? preissue_instr[80] : 
                              (N64)? preissue_instr[112] : 
                              (N60)? preissue_instr[144] : 1'b0;
  assign preissue_pkt_o[19] = (N61)? preissue_instr[17] : 
                              (N62)? preissue_instr[49] : 
                              (N63)? preissue_instr[81] : 
                              (N64)? preissue_instr[113] : 
                              (N60)? preissue_instr[145] : 1'b0;
  assign preissue_pkt_o[20] = (N61)? preissue_instr[18] : 
                              (N62)? preissue_instr[50] : 
                              (N63)? preissue_instr[82] : 
                              (N64)? preissue_instr[114] : 
                              (N60)? preissue_instr[146] : 1'b0;
  assign preissue_pkt_o[21] = (N61)? preissue_instr[19] : 
                              (N62)? preissue_instr[51] : 
                              (N63)? preissue_instr[83] : 
                              (N64)? preissue_instr[115] : 
                              (N60)? preissue_instr[147] : 1'b0;
  assign preissue_pkt_o[22] = (N61)? preissue_instr[20] : 
                              (N62)? preissue_instr[52] : 
                              (N63)? preissue_instr[84] : 
                              (N64)? preissue_instr[116] : 
                              (N60)? preissue_instr[148] : 1'b0;
  assign preissue_pkt_o[23] = (N61)? preissue_instr[21] : 
                              (N62)? preissue_instr[53] : 
                              (N63)? preissue_instr[85] : 
                              (N64)? preissue_instr[117] : 
                              (N60)? preissue_instr[149] : 1'b0;
  assign preissue_pkt_o[24] = (N61)? preissue_instr[22] : 
                              (N62)? preissue_instr[54] : 
                              (N63)? preissue_instr[86] : 
                              (N64)? preissue_instr[118] : 
                              (N60)? preissue_instr[150] : 1'b0;
  assign preissue_pkt_o[25] = (N61)? preissue_instr[23] : 
                              (N62)? preissue_instr[55] : 
                              (N63)? preissue_instr[87] : 
                              (N64)? preissue_instr[119] : 
                              (N60)? preissue_instr[151] : 1'b0;
  assign preissue_pkt_o[26] = (N61)? preissue_instr[24] : 
                              (N62)? preissue_instr[56] : 
                              (N63)? preissue_instr[88] : 
                              (N64)? preissue_instr[120] : 
                              (N60)? preissue_instr[152] : 1'b0;
  assign preissue_pkt_o[27] = (N61)? preissue_instr[25] : 
                              (N62)? preissue_instr[57] : 
                              (N63)? preissue_instr[89] : 
                              (N64)? preissue_instr[121] : 
                              (N60)? preissue_instr[153] : 1'b0;
  assign preissue_pkt_o[28] = (N61)? preissue_instr[26] : 
                              (N62)? preissue_instr[58] : 
                              (N63)? preissue_instr[90] : 
                              (N64)? preissue_instr[122] : 
                              (N60)? preissue_instr[154] : 1'b0;
  assign preissue_pkt_o[29] = (N61)? preissue_instr[27] : 
                              (N62)? preissue_instr[59] : 
                              (N63)? preissue_instr[91] : 
                              (N64)? preissue_instr[123] : 
                              (N60)? preissue_instr[155] : 1'b0;
  assign preissue_pkt_o[30] = (N61)? preissue_instr[28] : 
                              (N62)? preissue_instr[60] : 
                              (N63)? preissue_instr[92] : 
                              (N64)? preissue_instr[124] : 
                              (N60)? preissue_instr[156] : 1'b0;
  assign preissue_pkt_o[31] = (N61)? preissue_instr[29] : 
                              (N62)? preissue_instr[61] : 
                              (N63)? preissue_instr[93] : 
                              (N64)? preissue_instr[125] : 
                              (N60)? preissue_instr[157] : 1'b0;
  assign preissue_pkt_o[32] = (N61)? preissue_instr[30] : 
                              (N62)? preissue_instr[62] : 
                              (N63)? preissue_instr[94] : 
                              (N64)? preissue_instr[126] : 
                              (N60)? preissue_instr[158] : 1'b0;
  assign preissue_pkt_o[33] = (N61)? preissue_instr[31] : 
                              (N62)? preissue_instr[63] : 
                              (N63)? preissue_instr[95] : 
                              (N64)? preissue_instr[127] : 
                              (N60)? preissue_instr[159] : 1'b0;
  assign ack = fe_queue_ready_and_o & fe_queue_v_i;
  assign full = N69 & N70;
  assign N79 = ~ack;
  assign N80 = ack;
  assign N81 = ~1'b1;
  assign N90 = ~read_i;
  assign N91 = read_i;
  assign N92 = ~read_catchup;
  assign N101 = ~cmt_i;
  assign N102 = cmt_i;
  assign N103 = ~deq_catchup;
  assign N112 = roll_i | clr_i;
  assign N113 = ~N112;
  assign N121 = N137;
  assign N136 = ~clr_i;
  assign N137 = roll_i & N136;
  assign N138 = ~clr_i;
  assign preissue_v = N642 | N646;
  assign N642 = N641 | roll_i;
  assign N641 = N639 & N640;
  assign N639 = N638 | read[0];
  assign N638 = N637 | read[1];
  assign N637 = read[3] | read[2];
  assign N640 = ~empty_n;
  assign N646 = N645 & empty;
  assign N645 = N644 | enq[0];
  assign N644 = N643 | enq[1];
  assign N643 = enq[3] | enq[2];
  assign _2_net_ = ~bypass_preissue;
  assign _0_net_ = N648 | enq[0];
  assign N648 = N647 | enq[1];
  assign N647 = enq[3] | enq[2];
  assign N153 = ~bypass_preissue;
  assign N154 = ~N649;
  assign N649 = queue_instr_raw_0__1_ & queue_instr_raw_0__0_;
  assign preissue_size_0__0_ = N154;
  assign N155 = ~N650;
  assign N650 = queue_instr_raw_1__1_ & queue_instr_raw_1__0_;
  assign preissue_size_1__0_ = N155;
  assign N156 = ~N651;
  assign N651 = queue_instr_raw_2__1_ & queue_instr_raw_2__0_;
  assign preissue_size_2__0_ = N156;
  assign N157 = ~N652;
  assign N652 = queue_instr_raw_3__1_ & queue_instr_raw_3__0_;
  assign preissue_size_3__0_ = N157;
  assign N158 = ~N653;
  assign N653 = queue_instr_raw_4__1_ & queue_instr_raw_4__0_;
  assign preissue_size_4__0_ = N158;
  assign N178 = ~N171;
  assign N179 = ~N172;
  assign N180 = ~N175;
  assign N181 = ~N176;
  assign N182 = ~N177;
  assign N194 = ~N173;
  assign N198 = ~N174;
  assign N204 = N660 | N661;
  assign N660 = N658 | N659;
  assign N658 = N656 | N657;
  assign N656 = N654 | N655;
  assign N654 = ~N188;
  assign N655 = ~N193;
  assign N657 = ~N197;
  assign N659 = ~N201;
  assign N661 = ~N203;
  assign N216 = N668 | N669;
  assign N668 = N666 | N667;
  assign N666 = N664 | N665;
  assign N664 = N662 | N663;
  assign N662 = ~N205;
  assign N663 = ~N208;
  assign N665 = ~N210;
  assign N667 = ~N212;
  assign N669 = ~N215;
  assign N219 = ~N218;
  assign N221 = ~N220;
  assign N223 = ~N222;
  assign N227 = ~N226;
  assign N234 = N674 | N675;
  assign N674 = N672 | N673;
  assign N672 = N670 | N671;
  assign N670 = ~N229;
  assign N671 = ~N230;
  assign N673 = ~N232;
  assign N675 = ~N233;
  assign N245 = N181 | N680;
  assign N680 = N182 | N679;
  assign N679 = N236 | N678;
  assign N678 = N239 | N677;
  assign N677 = N241 | N676;
  assign N676 = N242 | N244;
  assign N246 = ~preissue_pkt_o[33];
  assign N247 = ~preissue_pkt_o[32];
  assign N248 = ~preissue_pkt_o[31];
  assign N249 = ~preissue_pkt_o[30];
  assign N250 = ~preissue_pkt_o[29];
  assign N251 = ~preissue_pkt_o[28];
  assign N252 = ~preissue_pkt_o[27];
  assign N253 = ~preissue_pkt_o[26];
  assign N254 = ~preissue_pkt_o[25];
  assign N255 = ~preissue_pkt_o[16];
  assign N256 = ~preissue_pkt_o[14];
  assign N257 = ~preissue_pkt_o[13];
  assign N258 = ~preissue_pkt_o[12];
  assign N259 = ~preissue_pkt_o[11];
  assign N260 = ~preissue_pkt_o[10];
  assign N261 = ~preissue_pkt_o[9];
  assign N262 = ~preissue_pkt_o[8];
  assign N263 = ~preissue_pkt_o[7];
  assign N264 = ~preissue_pkt_o[6];
  assign N288 = ~preissue_pkt_o[23];
  assign N289 = ~preissue_pkt_o[22];
  assign N292 = ~preissue_pkt_o[24];
  assign N293 = ~preissue_pkt_o[23];
  assign N296 = ~preissue_pkt_o[24];
  assign N297 = ~preissue_pkt_o[23];
  assign N298 = ~preissue_pkt_o[22];
  assign N301 = ~preissue_pkt_o[24];
  assign N302 = ~preissue_pkt_o[22];
  assign N305 = N682 | N304;
  assign N682 = N681 | N300;
  assign N681 = N291 | N295;
  assign N306 = ~N305;
  assign N309 = ~N287;
  assign N312 = ~preissue_pkt_o[29];
  assign N313 = ~preissue_pkt_o[28];
  assign N314 = ~preissue_pkt_o[26];
  assign N315 = ~preissue_pkt_o[25];
  assign N316 = ~preissue_pkt_o[24];
  assign N317 = ~preissue_pkt_o[7];
  assign N318 = ~preissue_pkt_o[5];
  assign N319 = ~preissue_pkt_o[4];
  assign N332 = ~N331;
  assign N333 = ~preissue_pkt_o[31];
  assign N334 = ~preissue_pkt_o[30];
  assign N335 = ~preissue_pkt_o[27];
  assign N336 = ~preissue_pkt_o[23];
  assign N337 = ~preissue_pkt_o[22];
  assign N343 = ~preissue_pkt_o[31];
  assign N344 = ~preissue_pkt_o[30];
  assign N345 = ~preissue_pkt_o[27];
  assign N346 = ~preissue_pkt_o[23];
  assign N352 = ~preissue_pkt_o[31];
  assign N353 = ~preissue_pkt_o[30];
  assign N354 = ~preissue_pkt_o[27];
  assign N355 = ~preissue_pkt_o[22];
  assign N361 = ~preissue_pkt_o[31];
  assign N362 = ~preissue_pkt_o[30];
  assign N363 = ~preissue_pkt_o[27];
  assign N369 = ~preissue_pkt_o[31];
  assign N370 = ~preissue_pkt_o[30];
  assign N371 = ~preissue_pkt_o[23];
  assign N372 = ~preissue_pkt_o[22];
  assign N378 = ~preissue_pkt_o[31];
  assign N379 = ~preissue_pkt_o[30];
  assign N380 = ~preissue_pkt_o[23];
  assign N386 = ~preissue_pkt_o[31];
  assign N387 = ~preissue_pkt_o[30];
  assign N388 = ~preissue_pkt_o[22];
  assign N394 = ~preissue_pkt_o[31];
  assign N395 = ~preissue_pkt_o[30];
  assign N401 = ~preissue_pkt_o[33];
  assign N402 = ~preissue_pkt_o[31];
  assign N403 = ~preissue_pkt_o[30];
  assign N404 = ~preissue_pkt_o[27];
  assign N405 = ~preissue_pkt_o[23];
  assign N411 = ~preissue_pkt_o[33];
  assign N412 = ~preissue_pkt_o[31];
  assign N413 = ~preissue_pkt_o[30];
  assign N414 = ~preissue_pkt_o[23];
  assign N415 = ~preissue_pkt_o[22];
  assign N421 = ~preissue_pkt_o[30];
  assign N422 = ~preissue_pkt_o[27];
  assign N423 = ~preissue_pkt_o[23];
  assign N424 = ~preissue_pkt_o[22];
  assign N425 = ~preissue_pkt_o[16];
  assign N426 = ~preissue_pkt_o[15];
  assign N427 = ~preissue_pkt_o[14];
  assign N436 = ~preissue_pkt_o[30];
  assign N437 = ~preissue_pkt_o[23];
  assign N438 = ~preissue_pkt_o[22];
  assign N439 = ~preissue_pkt_o[16];
  assign N440 = ~preissue_pkt_o[15];
  assign N441 = ~preissue_pkt_o[14];
  assign N450 = ~preissue_pkt_o[30];
  assign N451 = ~preissue_pkt_o[27];
  assign N452 = ~preissue_pkt_o[23];
  assign N453 = ~preissue_pkt_o[22];
  assign N454 = ~preissue_pkt_o[16];
  assign N455 = ~preissue_pkt_o[15];
  assign N464 = ~preissue_pkt_o[30];
  assign N465 = ~preissue_pkt_o[23];
  assign N466 = ~preissue_pkt_o[22];
  assign N467 = ~preissue_pkt_o[16];
  assign N468 = ~preissue_pkt_o[15];
  assign N477 = N694 | N476;
  assign N694 = N693 | N463;
  assign N693 = N692 | N449;
  assign N692 = N691 | N435;
  assign N691 = N690 | N420;
  assign N690 = N689 | N410;
  assign N689 = N688 | N400;
  assign N688 = N687 | N393;
  assign N687 = N686 | N385;
  assign N686 = N685 | N377;
  assign N685 = N684 | N368;
  assign N684 = N683 | N360;
  assign N683 = N342 | N351;
  assign N478 = ~preissue_pkt_o[31];
  assign N479 = ~preissue_pkt_o[27];
  assign N480 = ~preissue_pkt_o[23];
  assign N481 = ~preissue_pkt_o[22];
  assign N487 = ~preissue_pkt_o[31];
  assign N488 = ~preissue_pkt_o[27];
  assign N489 = ~preissue_pkt_o[23];
  assign N495 = ~preissue_pkt_o[31];
  assign N496 = ~preissue_pkt_o[27];
  assign N497 = ~preissue_pkt_o[22];
  assign N503 = ~preissue_pkt_o[31];
  assign N504 = ~preissue_pkt_o[27];
  assign N510 = ~preissue_pkt_o[31];
  assign N511 = ~preissue_pkt_o[23];
  assign N512 = ~preissue_pkt_o[22];
  assign N518 = ~preissue_pkt_o[31];
  assign N519 = ~preissue_pkt_o[23];
  assign N525 = ~preissue_pkt_o[31];
  assign N526 = ~preissue_pkt_o[22];
  assign N532 = ~preissue_pkt_o[31];
  assign N538 = ~preissue_pkt_o[27];
  assign N539 = ~preissue_pkt_o[23];
  assign N540 = ~preissue_pkt_o[22];
  assign N541 = ~preissue_pkt_o[16];
  assign N542 = ~preissue_pkt_o[15];
  assign N543 = ~preissue_pkt_o[14];
  assign N552 = ~preissue_pkt_o[23];
  assign N553 = ~preissue_pkt_o[22];
  assign N554 = ~preissue_pkt_o[16];
  assign N555 = ~preissue_pkt_o[15];
  assign N556 = ~preissue_pkt_o[14];
  assign N565 = N702 | N564;
  assign N702 = N701 | N551;
  assign N701 = N700 | N537;
  assign N700 = N699 | N531;
  assign N699 = N698 | N524;
  assign N698 = N697 | N517;
  assign N697 = N696 | N509;
  assign N696 = N695 | N502;
  assign N695 = N486 | N494;
  assign N566 = ~preissue_pkt_o[33];
  assign N569 = ~preissue_pkt_o[33];
  assign N573 = ~preissue_pkt_o[33];
  assign N575 = ~preissue_pkt_o[33];
  assign N577 = ~preissue_pkt_o[33];
  assign N578 = ~preissue_pkt_o[27];
  assign N579 = ~preissue_pkt_o[22];
  assign N587 = N568 | N710;
  assign N710 = N571 | N709;
  assign N709 = N572 | N708;
  assign N708 = N574 | N707;
  assign N707 = N576 | N706;
  assign N706 = N581 | N705;
  assign N705 = N583 | N704;
  assign N704 = N584 | N703;
  assign N703 = N585 | N586;
  assign N588 = ~N587;
  assign N589 = N588;
  assign N592 = ~N565;
  assign N593 = N592;
  assign N598 = ~N234;
  assign N599 = N598;
  assign _6_net_ = ~bypass_issue;
  assign _4_net_ = N712 | enq[0];
  assign N712 = N711 | enq[1];
  assign N711 = enq[3] | enq[2];
  assign fe_queue_ready_and_o = ~full;
  assign N600 = ~issue_pkt_o[262];
  assign issue_pkt_o[263] = en_i & N713;
  assign N713 = ~empty;
  assign issue_pkt_o[262] = N621 & N714;
  assign N714 = ~illegal_instr_lo;
  assign issue_pkt_o[257] = N618 & illegal_instr_lo;

endmodule



module bsg_mem_2r1w_sync_width_p66_els_p32
(
  clk_i,
  reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r0_v_i,
  r0_addr_i,
  r0_data_o,
  r1_v_i,
  r1_addr_i,
  r1_data_o
);

  input [4:0] w_addr_i;
  input [65:0] w_data_i;
  input [4:0] r0_addr_i;
  output [65:0] r0_data_o;
  input [4:0] r1_addr_i;
  output [65:0] r1_data_o;
  input clk_i;
  input reset_i;
  input w_v_i;
  input r0_v_i;
  input r1_v_i;
  wire [65:0] r0_data_o,r1_data_o;

  bsg_mem_2r1w_sync_synth
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r0_v_i(r0_v_i),
    .r0_addr_i(r0_addr_i),
    .r0_data_o(r0_data_o),
    .r1_v_i(r1_v_i),
    .r1_addr_i(r1_addr_i),
    .r1_data_o(r1_data_o)
  );


endmodule



module bsg_dff_width_p66
(
  clk_i,
  data_i,
  data_o
);

  input [65:0] data_i;
  output [65:0] data_o;
  input clk_i;
  wire [65:0] data_o;
  reg data_o_65_sv2v_reg,data_o_64_sv2v_reg,data_o_63_sv2v_reg,data_o_62_sv2v_reg,
  data_o_61_sv2v_reg,data_o_60_sv2v_reg,data_o_59_sv2v_reg,data_o_58_sv2v_reg,
  data_o_57_sv2v_reg,data_o_56_sv2v_reg,data_o_55_sv2v_reg,data_o_54_sv2v_reg,
  data_o_53_sv2v_reg,data_o_52_sv2v_reg,data_o_51_sv2v_reg,data_o_50_sv2v_reg,
  data_o_49_sv2v_reg,data_o_48_sv2v_reg,data_o_47_sv2v_reg,data_o_46_sv2v_reg,data_o_45_sv2v_reg,
  data_o_44_sv2v_reg,data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,
  data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,
  data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,
  data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,
  data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,
  data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,
  data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,
  data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_width_p3
(
  clk_i,
  data_i,
  data_o
);

  input [2:0] data_i;
  output [2:0] data_o;
  input clk_i;
  wire [2:0] data_o;
  reg data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_width_p5
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [4:0] data_i;
  output [4:0] data_o;
  input clk_i;
  input en_i;
  wire [4:0] data_o;
  reg data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_width_p66
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [65:0] data_i;
  output [65:0] data_o;
  input clk_i;
  input en_i;
  wire [65:0] data_o;
  reg data_o_65_sv2v_reg,data_o_64_sv2v_reg,data_o_63_sv2v_reg,data_o_62_sv2v_reg,
  data_o_61_sv2v_reg,data_o_60_sv2v_reg,data_o_59_sv2v_reg,data_o_58_sv2v_reg,
  data_o_57_sv2v_reg,data_o_56_sv2v_reg,data_o_55_sv2v_reg,data_o_54_sv2v_reg,
  data_o_53_sv2v_reg,data_o_52_sv2v_reg,data_o_51_sv2v_reg,data_o_50_sv2v_reg,
  data_o_49_sv2v_reg,data_o_48_sv2v_reg,data_o_47_sv2v_reg,data_o_46_sv2v_reg,data_o_45_sv2v_reg,
  data_o_44_sv2v_reg,data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,
  data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,
  data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,
  data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,
  data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,
  data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,
  data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,
  data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bp_be_regfile_00_66_2_1
(
  clk_i,
  reset_i,
  rs_r_v_i,
  rs_addr_i,
  rs_data_o,
  rd_w_v_i,
  rd_addr_i,
  rd_data_i
);

  input [1:0] rs_r_v_i;
  input [9:0] rs_addr_i;
  output [131:0] rs_data_o;
  input [4:0] rd_addr_i;
  input [65:0] rd_data_i;
  input clk_i;
  input reset_i;
  input rd_w_v_i;
  wire [131:0] rs_data_o,rs_data_lo;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,\bypass_0_.zero_rs ,N10,\bypass_0_.fwd_rs ,
  \bypass_0_.zero_rs_r ,\bypass_0_.fwd_rs_r ,\bypass_0_.rs_r_v_r ,N11,N12,N13,N14,N15,
  \bypass_0_.replace_rs ,N16,_2_net_,N17,\bypass_1_.zero_rs ,N18,\bypass_1_.fwd_rs ,
  \bypass_1_.zero_rs_r ,\bypass_1_.fwd_rs_r ,\bypass_1_.rs_r_v_r ,N19,N20,N21,N22,
  N23,\bypass_1_.replace_rs ,N24,_5_net_,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,
  N35,N36,N37,N38,N39;
  wire [1:0] rs_v_li;
  wire [65:0] rd_data_r,\bypass_0_.fwd_data_lo ,\bypass_0_.rs_data_n ,\bypass_0_.rs_data_r ,
  \bypass_1_.fwd_data_lo ,\bypass_1_.rs_data_n ,\bypass_1_.rs_data_r ;
  wire [4:0] \bypass_0_.rs_addr_r ,\bypass_1_.rs_addr_r ;

  bsg_mem_2r1w_sync_width_p66_els_p32
  \tworonew.rf 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(rd_w_v_i),
    .w_addr_i(rd_addr_i),
    .w_data_i(rd_data_i),
    .r0_v_i(rs_v_li[0]),
    .r0_addr_i(rs_addr_i[4:0]),
    .r0_data_o(rs_data_lo[65:0]),
    .r1_v_i(rs_v_li[1]),
    .r1_addr_i(rs_addr_i[9:5]),
    .r1_data_o(rs_data_lo[131:66])
  );


  bsg_dff_width_p66
  rd_reg
  (
    .clk_i(clk_i),
    .data_i(rd_data_i),
    .data_o(rd_data_r)
  );

  assign N10 = rd_addr_i == rs_addr_i[4:0];

  bsg_dff_width_p3
  \bypass_0_.rs_r_v_reg 
  (
    .clk_i(clk_i),
    .data_i({ \bypass_0_.zero_rs , \bypass_0_.fwd_rs , rs_r_v_i[0:0] }),
    .data_o({ \bypass_0_.zero_rs_r , \bypass_0_.fwd_rs_r , \bypass_0_.rs_r_v_r  })
  );


  bsg_dff_en_width_p5
  \bypass_0_.rs_addr_reg 
  (
    .clk_i(clk_i),
    .data_i(rs_addr_i[4:0]),
    .en_i(rs_r_v_i[0]),
    .data_o(\bypass_0_.rs_addr_r )
  );

  assign N15 = \bypass_0_.rs_addr_r  == rd_addr_i;

  bsg_dff_en_width_p66
  \bypass_0_.rs_data_reg 
  (
    .clk_i(clk_i),
    .data_i(\bypass_0_.rs_data_n ),
    .en_i(_2_net_),
    .data_o(\bypass_0_.rs_data_r )
  );

  assign N18 = rd_addr_i == rs_addr_i[9:5];

  bsg_dff_width_p3
  \bypass_1_.rs_r_v_reg 
  (
    .clk_i(clk_i),
    .data_i({ \bypass_1_.zero_rs , \bypass_1_.fwd_rs , rs_r_v_i[1:1] }),
    .data_o({ \bypass_1_.zero_rs_r , \bypass_1_.fwd_rs_r , \bypass_1_.rs_r_v_r  })
  );


  bsg_dff_en_width_p5
  \bypass_1_.rs_addr_reg 
  (
    .clk_i(clk_i),
    .data_i(rs_addr_i[9:5]),
    .en_i(rs_r_v_i[1]),
    .data_o(\bypass_1_.rs_addr_r )
  );

  assign N23 = \bypass_1_.rs_addr_r  == rd_addr_i;

  bsg_dff_en_width_p66
  \bypass_1_.rs_data_reg 
  (
    .clk_i(clk_i),
    .data_i(\bypass_1_.rs_data_n ),
    .en_i(_5_net_),
    .data_o(\bypass_1_.rs_data_r )
  );

  assign N26 = rs_addr_i[3] | rs_addr_i[4];
  assign N27 = rs_addr_i[2] | N26;
  assign N28 = rs_addr_i[1] | N27;
  assign N29 = rs_addr_i[0] | N28;
  assign N30 = ~N29;
  assign N31 = rs_addr_i[8] | rs_addr_i[9];
  assign N32 = rs_addr_i[7] | N31;
  assign N33 = rs_addr_i[6] | N32;
  assign N34 = rs_addr_i[5] | N33;
  assign N35 = ~N34;
  assign \bypass_0_.fwd_data_lo  = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N14)? rd_data_r : 
                                   (N12)? rs_data_lo[65:0] : 1'b0;
  assign N0 = \bypass_0_.zero_rs_r ;
  assign \bypass_0_.rs_data_n  = (N1)? rd_data_i : 
                                 (N2)? \bypass_0_.fwd_data_lo  : 1'b0;
  assign N1 = \bypass_0_.replace_rs ;
  assign N2 = N16;
  assign rs_data_o[65:0] = (N3)? \bypass_0_.fwd_data_lo  : 
                           (N4)? \bypass_0_.rs_data_r  : 1'b0;
  assign N3 = \bypass_0_.rs_r_v_r ;
  assign N4 = N17;
  assign \bypass_1_.fwd_data_lo  = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N22)? rd_data_r : 
                                   (N20)? rs_data_lo[131:66] : 1'b0;
  assign N5 = \bypass_1_.zero_rs_r ;
  assign \bypass_1_.rs_data_n  = (N6)? rd_data_i : 
                                 (N7)? \bypass_1_.fwd_data_lo  : 1'b0;
  assign N6 = \bypass_1_.replace_rs ;
  assign N7 = N24;
  assign rs_data_o[131:66] = (N8)? \bypass_1_.fwd_data_lo  : 
                             (N9)? \bypass_1_.rs_data_r  : 1'b0;
  assign N8 = \bypass_1_.rs_r_v_r ;
  assign N9 = N25;
  assign \bypass_0_.zero_rs  = rs_r_v_i[0] & N30;
  assign \bypass_0_.fwd_rs  = N36 & N10;
  assign N36 = rd_w_v_i & rs_r_v_i[0];
  assign N11 = \bypass_0_.fwd_rs_r  | \bypass_0_.zero_rs_r ;
  assign N12 = ~N11;
  assign N13 = ~\bypass_0_.zero_rs_r ;
  assign N14 = \bypass_0_.fwd_rs_r  & N13;
  assign \bypass_0_.replace_rs  = rd_w_v_i & N15;
  assign N16 = ~\bypass_0_.replace_rs ;
  assign _2_net_ = \bypass_0_.rs_r_v_r  | \bypass_0_.replace_rs ;
  assign rs_v_li[0] = rs_r_v_i[0] & N37;
  assign N37 = ~\bypass_0_.fwd_rs ;
  assign N17 = ~\bypass_0_.rs_r_v_r ;
  assign \bypass_1_.zero_rs  = rs_r_v_i[1] & N35;
  assign \bypass_1_.fwd_rs  = N38 & N18;
  assign N38 = rd_w_v_i & rs_r_v_i[1];
  assign N19 = \bypass_1_.fwd_rs_r  | \bypass_1_.zero_rs_r ;
  assign N20 = ~N19;
  assign N21 = ~\bypass_1_.zero_rs_r ;
  assign N22 = \bypass_1_.fwd_rs_r  & N21;
  assign \bypass_1_.replace_rs  = rd_w_v_i & N23;
  assign N24 = ~\bypass_1_.replace_rs ;
  assign _5_net_ = \bypass_1_.rs_r_v_r  | \bypass_1_.replace_rs ;
  assign rs_v_li[1] = rs_r_v_i[1] & N39;
  assign N39 = ~\bypass_1_.fwd_rs ;
  assign N25 = ~\bypass_1_.rs_r_v_r ;

endmodule



module bp_be_int_regfile_00
(
  clk_i,
  reset_i,
  rs_r_v_i,
  rs_addr_i,
  rs_data_o,
  rd_w_v_i,
  rd_addr_i,
  rd_data_i
);

  input [1:0] rs_r_v_i;
  input [9:0] rs_addr_i;
  output [131:0] rs_data_o;
  input [4:0] rd_addr_i;
  input [65:0] rd_data_i;
  input clk_i;
  input reset_i;
  input rd_w_v_i;
  wire [131:0] rs_data_o;

  bp_be_regfile_00_66_2_1
  regfile
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .rs_r_v_i(rs_r_v_i),
    .rs_addr_i(rs_addr_i),
    .rs_data_o(rs_data_o),
    .rd_w_v_i(rd_w_v_i),
    .rd_addr_i(rd_addr_i),
    .rd_data_i(rd_data_i)
  );


endmodule



module bsg_mem_3r1w_sync_width_p66_els_p32
(
  clk_i,
  reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r0_v_i,
  r0_addr_i,
  r0_data_o,
  r1_v_i,
  r1_addr_i,
  r1_data_o,
  r2_v_i,
  r2_addr_i,
  r2_data_o
);

  input [4:0] w_addr_i;
  input [65:0] w_data_i;
  input [4:0] r0_addr_i;
  output [65:0] r0_data_o;
  input [4:0] r1_addr_i;
  output [65:0] r1_data_o;
  input [4:0] r2_addr_i;
  output [65:0] r2_data_o;
  input clk_i;
  input reset_i;
  input w_v_i;
  input r0_v_i;
  input r1_v_i;
  input r2_v_i;
  wire [65:0] r0_data_o,r1_data_o,r2_data_o;

  bsg_mem_3r1w_sync_synth
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r0_v_i(r0_v_i),
    .r0_addr_i(r0_addr_i),
    .r0_data_o(r0_data_o),
    .r1_v_i(r1_v_i),
    .r1_addr_i(r1_addr_i),
    .r1_data_o(r1_data_o),
    .r2_v_i(r2_v_i),
    .r2_addr_i(r2_addr_i),
    .r2_data_o(r2_data_o)
  );


endmodule



module bp_be_regfile_00_66_3_0
(
  clk_i,
  reset_i,
  rs_r_v_i,
  rs_addr_i,
  rs_data_o,
  rd_w_v_i,
  rd_addr_i,
  rd_data_i
);

  input [2:0] rs_r_v_i;
  input [14:0] rs_addr_i;
  output [197:0] rs_data_o;
  input [4:0] rd_addr_i;
  input [65:0] rd_data_i;
  input clk_i;
  input reset_i;
  input rd_w_v_i;
  wire [197:0] rs_data_o,rs_data_lo;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,\bypass_0_.fwd_rs ,
  \bypass_0_.zero_rs_r ,\bypass_0_.fwd_rs_r ,\bypass_0_.rs_r_v_r ,N16,N17,N18,N19,N20,
  \bypass_0_.replace_rs ,N21,_2_net_,N22,N23,\bypass_1_.fwd_rs ,
  \bypass_1_.zero_rs_r ,\bypass_1_.fwd_rs_r ,\bypass_1_.rs_r_v_r ,N24,N25,N26,N27,N28,
  \bypass_1_.replace_rs ,N29,_5_net_,N30,N31,\bypass_2_.fwd_rs ,\bypass_2_.zero_rs_r ,
  \bypass_2_.fwd_rs_r ,\bypass_2_.rs_r_v_r ,N32,N33,N34,N35,N36,\bypass_2_.replace_rs ,N37,
  _8_net_,N38,N39,N40,N41,N42,N43,N44;
  wire [2:0] rs_v_li;
  wire [65:0] rd_data_r,\bypass_0_.fwd_data_lo ,\bypass_0_.rs_data_n ,\bypass_0_.rs_data_r ,
  \bypass_1_.fwd_data_lo ,\bypass_1_.rs_data_n ,\bypass_1_.rs_data_r ,
  \bypass_2_.fwd_data_lo ,\bypass_2_.rs_data_n ,\bypass_2_.rs_data_r ;
  wire [4:0] \bypass_0_.rs_addr_r ,\bypass_1_.rs_addr_r ,\bypass_2_.rs_addr_r ;

  bsg_mem_3r1w_sync_width_p66_els_p32
  \threeronew.rf 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(rd_w_v_i),
    .w_addr_i(rd_addr_i),
    .w_data_i(rd_data_i),
    .r0_v_i(rs_v_li[0]),
    .r0_addr_i(rs_addr_i[4:0]),
    .r0_data_o(rs_data_lo[65:0]),
    .r1_v_i(rs_v_li[1]),
    .r1_addr_i(rs_addr_i[9:5]),
    .r1_data_o(rs_data_lo[131:66]),
    .r2_v_i(rs_v_li[2]),
    .r2_addr_i(rs_addr_i[14:10]),
    .r2_data_o(rs_data_lo[197:132])
  );


  bsg_dff_width_p66
  rd_reg
  (
    .clk_i(clk_i),
    .data_i(rd_data_i),
    .data_o(rd_data_r)
  );

  assign N15 = rd_addr_i == rs_addr_i[4:0];

  bsg_dff_width_p3
  \bypass_0_.rs_r_v_reg 
  (
    .clk_i(clk_i),
    .data_i({ 1'b0, \bypass_0_.fwd_rs , rs_r_v_i[0:0] }),
    .data_o({ \bypass_0_.zero_rs_r , \bypass_0_.fwd_rs_r , \bypass_0_.rs_r_v_r  })
  );


  bsg_dff_en_width_p5
  \bypass_0_.rs_addr_reg 
  (
    .clk_i(clk_i),
    .data_i(rs_addr_i[4:0]),
    .en_i(rs_r_v_i[0]),
    .data_o(\bypass_0_.rs_addr_r )
  );

  assign N20 = \bypass_0_.rs_addr_r  == rd_addr_i;

  bsg_dff_en_width_p66
  \bypass_0_.rs_data_reg 
  (
    .clk_i(clk_i),
    .data_i(\bypass_0_.rs_data_n ),
    .en_i(_2_net_),
    .data_o(\bypass_0_.rs_data_r )
  );

  assign N23 = rd_addr_i == rs_addr_i[9:5];

  bsg_dff_width_p3
  \bypass_1_.rs_r_v_reg 
  (
    .clk_i(clk_i),
    .data_i({ 1'b0, \bypass_1_.fwd_rs , rs_r_v_i[1:1] }),
    .data_o({ \bypass_1_.zero_rs_r , \bypass_1_.fwd_rs_r , \bypass_1_.rs_r_v_r  })
  );


  bsg_dff_en_width_p5
  \bypass_1_.rs_addr_reg 
  (
    .clk_i(clk_i),
    .data_i(rs_addr_i[9:5]),
    .en_i(rs_r_v_i[1]),
    .data_o(\bypass_1_.rs_addr_r )
  );

  assign N28 = \bypass_1_.rs_addr_r  == rd_addr_i;

  bsg_dff_en_width_p66
  \bypass_1_.rs_data_reg 
  (
    .clk_i(clk_i),
    .data_i(\bypass_1_.rs_data_n ),
    .en_i(_5_net_),
    .data_o(\bypass_1_.rs_data_r )
  );

  assign N31 = rd_addr_i == rs_addr_i[14:10];

  bsg_dff_width_p3
  \bypass_2_.rs_r_v_reg 
  (
    .clk_i(clk_i),
    .data_i({ 1'b0, \bypass_2_.fwd_rs , rs_r_v_i[2:2] }),
    .data_o({ \bypass_2_.zero_rs_r , \bypass_2_.fwd_rs_r , \bypass_2_.rs_r_v_r  })
  );


  bsg_dff_en_width_p5
  \bypass_2_.rs_addr_reg 
  (
    .clk_i(clk_i),
    .data_i(rs_addr_i[14:10]),
    .en_i(rs_r_v_i[2]),
    .data_o(\bypass_2_.rs_addr_r )
  );

  assign N36 = \bypass_2_.rs_addr_r  == rd_addr_i;

  bsg_dff_en_width_p66
  \bypass_2_.rs_data_reg 
  (
    .clk_i(clk_i),
    .data_i(\bypass_2_.rs_data_n ),
    .en_i(_8_net_),
    .data_o(\bypass_2_.rs_data_r )
  );

  assign \bypass_0_.fwd_data_lo  = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N19)? rd_data_r : 
                                   (N17)? rs_data_lo[65:0] : 1'b0;
  assign N0 = \bypass_0_.zero_rs_r ;
  assign \bypass_0_.rs_data_n  = (N1)? rd_data_i : 
                                 (N2)? \bypass_0_.fwd_data_lo  : 1'b0;
  assign N1 = \bypass_0_.replace_rs ;
  assign N2 = N21;
  assign rs_data_o[65:0] = (N3)? \bypass_0_.fwd_data_lo  : 
                           (N4)? \bypass_0_.rs_data_r  : 1'b0;
  assign N3 = \bypass_0_.rs_r_v_r ;
  assign N4 = N22;
  assign \bypass_1_.fwd_data_lo  = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N27)? rd_data_r : 
                                   (N25)? rs_data_lo[131:66] : 1'b0;
  assign N5 = \bypass_1_.zero_rs_r ;
  assign \bypass_1_.rs_data_n  = (N6)? rd_data_i : 
                                 (N7)? \bypass_1_.fwd_data_lo  : 1'b0;
  assign N6 = \bypass_1_.replace_rs ;
  assign N7 = N29;
  assign rs_data_o[131:66] = (N8)? \bypass_1_.fwd_data_lo  : 
                             (N9)? \bypass_1_.rs_data_r  : 1'b0;
  assign N8 = \bypass_1_.rs_r_v_r ;
  assign N9 = N30;
  assign \bypass_2_.fwd_data_lo  = (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N35)? rd_data_r : 
                                   (N33)? rs_data_lo[197:132] : 1'b0;
  assign N10 = \bypass_2_.zero_rs_r ;
  assign \bypass_2_.rs_data_n  = (N11)? rd_data_i : 
                                 (N12)? \bypass_2_.fwd_data_lo  : 1'b0;
  assign N11 = \bypass_2_.replace_rs ;
  assign N12 = N37;
  assign rs_data_o[197:132] = (N13)? \bypass_2_.fwd_data_lo  : 
                              (N14)? \bypass_2_.rs_data_r  : 1'b0;
  assign N13 = \bypass_2_.rs_r_v_r ;
  assign N14 = N38;
  assign \bypass_0_.fwd_rs  = N39 & N15;
  assign N39 = rd_w_v_i & rs_r_v_i[0];
  assign N16 = \bypass_0_.fwd_rs_r  | \bypass_0_.zero_rs_r ;
  assign N17 = ~N16;
  assign N18 = ~\bypass_0_.zero_rs_r ;
  assign N19 = \bypass_0_.fwd_rs_r  & N18;
  assign \bypass_0_.replace_rs  = rd_w_v_i & N20;
  assign N21 = ~\bypass_0_.replace_rs ;
  assign _2_net_ = \bypass_0_.rs_r_v_r  | \bypass_0_.replace_rs ;
  assign rs_v_li[0] = rs_r_v_i[0] & N40;
  assign N40 = ~\bypass_0_.fwd_rs ;
  assign N22 = ~\bypass_0_.rs_r_v_r ;
  assign \bypass_1_.fwd_rs  = N41 & N23;
  assign N41 = rd_w_v_i & rs_r_v_i[1];
  assign N24 = \bypass_1_.fwd_rs_r  | \bypass_1_.zero_rs_r ;
  assign N25 = ~N24;
  assign N26 = ~\bypass_1_.zero_rs_r ;
  assign N27 = \bypass_1_.fwd_rs_r  & N26;
  assign \bypass_1_.replace_rs  = rd_w_v_i & N28;
  assign N29 = ~\bypass_1_.replace_rs ;
  assign _5_net_ = \bypass_1_.rs_r_v_r  | \bypass_1_.replace_rs ;
  assign rs_v_li[1] = rs_r_v_i[1] & N42;
  assign N42 = ~\bypass_1_.fwd_rs ;
  assign N30 = ~\bypass_1_.rs_r_v_r ;
  assign \bypass_2_.fwd_rs  = N43 & N31;
  assign N43 = rd_w_v_i & rs_r_v_i[2];
  assign N32 = \bypass_2_.fwd_rs_r  | \bypass_2_.zero_rs_r ;
  assign N33 = ~N32;
  assign N34 = ~\bypass_2_.zero_rs_r ;
  assign N35 = \bypass_2_.fwd_rs_r  & N34;
  assign \bypass_2_.replace_rs  = rd_w_v_i & N36;
  assign N37 = ~\bypass_2_.replace_rs ;
  assign _8_net_ = \bypass_2_.rs_r_v_r  | \bypass_2_.replace_rs ;
  assign rs_v_li[2] = rs_r_v_i[2] & N44;
  assign N44 = ~\bypass_2_.fwd_rs ;
  assign N38 = ~\bypass_2_.rs_r_v_r ;

endmodule



module bp_be_fp_regfile_00
(
  clk_i,
  reset_i,
  rs_r_v_i,
  rs_addr_i,
  rs_data_o,
  rd_w_v_i,
  rd_addr_i,
  rd_data_i
);

  input [2:0] rs_r_v_i;
  input [14:0] rs_addr_i;
  output [197:0] rs_data_o;
  input [4:0] rd_addr_i;
  input [65:0] rd_data_i;
  input clk_i;
  input reset_i;
  input rd_w_v_i;
  wire [197:0] rs_data_o;

  bp_be_regfile_00_66_3_0
  regfile
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .rs_r_v_i(rs_r_v_i),
    .rs_addr_i(rs_addr_i),
    .rs_data_o(rs_data_o),
    .rd_w_v_i(rd_w_v_i),
    .rd_addr_i(rd_addr_i),
    .rd_data_i(rd_data_i)
  );


endmodule



module bp_be_scheduler_00
(
  clk_i,
  reset_i,
  issue_pkt_o,
  expected_npc_i,
  clear_iss_i,
  suppress_iss_i,
  resume_i,
  decode_info_i,
  hazard_v_i,
  irq_pending_i,
  ispec_v_i,
  poison_isd_i,
  ordered_v_i,
  trans_info_i,
  fe_queue_i,
  fe_queue_v_i,
  fe_queue_ready_and_o,
  dispatch_pkt_o,
  commit_pkt_i,
  iwb_pkt_i,
  fwb_pkt_i,
  late_wb_pkt_i,
  late_wb_v_i,
  late_wb_force_i,
  late_wb_yumi_o
);

  output [263:0] issue_pkt_o;
  input [38:0] expected_npc_i;
  input [12:0] decode_info_i;
  input [32:0] trans_info_i;
  input [173:0] fe_queue_i;
  output [365:0] dispatch_pkt_o;
  input [213:0] commit_pkt_i;
  input [78:0] iwb_pkt_i;
  input [78:0] fwb_pkt_i;
  input [78:0] late_wb_pkt_i;
  input clk_i;
  input reset_i;
  input clear_iss_i;
  input suppress_iss_i;
  input resume_i;
  input hazard_v_i;
  input irq_pending_i;
  input ispec_v_i;
  input poison_isd_i;
  input ordered_v_i;
  input fe_queue_v_i;
  input late_wb_v_i;
  input late_wb_force_i;
  output fe_queue_ready_and_o;
  output late_wb_yumi_o;
  wire [263:0] issue_pkt_o;
  wire [365:0] dispatch_pkt_o;
  wire fe_queue_ready_and_o,late_wb_yumi_o,N0,N1,dispatch_pkt_o_361_,
  dispatch_pkt_o_360_,dispatch_pkt_o_359_,dispatch_pkt_o_358_,dispatch_pkt_o_357_,
  dispatch_pkt_o_356_,dispatch_pkt_o_355_,dispatch_pkt_o_354_,dispatch_pkt_o_353_,
  dispatch_pkt_o_352_,dispatch_pkt_o_351_,dispatch_pkt_o_350_,dispatch_pkt_o_349_,
  dispatch_pkt_o_348_,dispatch_pkt_o_347_,dispatch_pkt_o_346_,dispatch_pkt_o_345_,
  dispatch_pkt_o_344_,dispatch_pkt_o_343_,dispatch_pkt_o_342_,dispatch_pkt_o_341_,
  dispatch_pkt_o_340_,dispatch_pkt_o_339_,dispatch_pkt_o_338_,dispatch_pkt_o_337_,
  dispatch_pkt_o_336_,dispatch_pkt_o_335_,dispatch_pkt_o_334_,dispatch_pkt_o_333_,
  dispatch_pkt_o_332_,dispatch_pkt_o_331_,dispatch_pkt_o_330_,dispatch_pkt_o_329_,
  dispatch_pkt_o_328_,dispatch_pkt_o_327_,dispatch_pkt_o_326_,dispatch_pkt_o_325_,
  dispatch_pkt_o_324_,dispatch_pkt_o_323_,ptw_v_li,ptw_busy_lo,ptw_v_lo,ptw_itlb_fill_lo,
  ptw_dtlb_fill_lo,ptw_instr_page_fault_lo,ptw_load_page_fault_lo,ptw_store_page_fault_lo,
  resume_v,interrupt_v,be_exc_not_instr_li,fe_exc_not_instr_li,fe_instr_not_exc_li,
  fe_queue_en_li,fe_queue_read_li,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,
  walk_decode_li_pipe_mem_final_v_,be_exc_decode_li_pipe_mem_final_v_,
  be_exc_decode_li_irf_w_v_,be_exc_decode_li_frf_w_v_,be_exc_decode_li_dcache_mmu_v_,
  be_exc_decode_li_fu_op__t__5_,be_exc_decode_li_fu_op__t__4_,be_exc_decode_li_fu_op__t__3_,N14,N15,
  N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,
  N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,
  N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73;
  wire [2:0] ptw_count_lo,be_exc_count_li;
  wire [63:0] ptw_addr_lo,ptw_pte_lo,be_exc_vaddr_li;
  wire [38:0] preissue_pkt,fe_exc_vaddr_li;
  wire [65:0] irf_rs2,irf_rs1,frf_rs3,frf_rs2,frf_rs1,be_exc_data_li;
  wire [4:0] be_exc_imm_li;
  wire [31:0] be_exc_instr_li;
  assign dispatch_pkt_o[8] = 1'b0;
  assign dispatch_pkt_o[9] = 1'b0;
  assign dispatch_pkt_o[10] = 1'b0;
  assign dispatch_pkt_o[14] = 1'b0;
  assign dispatch_pkt_o[15] = 1'b0;
  assign dispatch_pkt_o[16] = 1'b0;
  assign dispatch_pkt_o[20] = 1'b0;
  assign dispatch_pkt_o[24] = 1'b0;
  assign dispatch_pkt_o[25] = 1'b0;
  assign dispatch_pkt_o[26] = 1'b0;
  assign dispatch_pkt_o[27] = 1'b0;
  assign dispatch_pkt_o_361_ = expected_npc_i[38];
  assign dispatch_pkt_o[361] = dispatch_pkt_o_361_;
  assign dispatch_pkt_o_360_ = expected_npc_i[37];
  assign dispatch_pkt_o[360] = dispatch_pkt_o_360_;
  assign dispatch_pkt_o_359_ = expected_npc_i[36];
  assign dispatch_pkt_o[359] = dispatch_pkt_o_359_;
  assign dispatch_pkt_o_358_ = expected_npc_i[35];
  assign dispatch_pkt_o[358] = dispatch_pkt_o_358_;
  assign dispatch_pkt_o_357_ = expected_npc_i[34];
  assign dispatch_pkt_o[357] = dispatch_pkt_o_357_;
  assign dispatch_pkt_o_356_ = expected_npc_i[33];
  assign dispatch_pkt_o[356] = dispatch_pkt_o_356_;
  assign dispatch_pkt_o_355_ = expected_npc_i[32];
  assign dispatch_pkt_o[355] = dispatch_pkt_o_355_;
  assign dispatch_pkt_o_354_ = expected_npc_i[31];
  assign dispatch_pkt_o[354] = dispatch_pkt_o_354_;
  assign dispatch_pkt_o_353_ = expected_npc_i[30];
  assign dispatch_pkt_o[353] = dispatch_pkt_o_353_;
  assign dispatch_pkt_o_352_ = expected_npc_i[29];
  assign dispatch_pkt_o[352] = dispatch_pkt_o_352_;
  assign dispatch_pkt_o_351_ = expected_npc_i[28];
  assign dispatch_pkt_o[351] = dispatch_pkt_o_351_;
  assign dispatch_pkt_o_350_ = expected_npc_i[27];
  assign dispatch_pkt_o[350] = dispatch_pkt_o_350_;
  assign dispatch_pkt_o_349_ = expected_npc_i[26];
  assign dispatch_pkt_o[349] = dispatch_pkt_o_349_;
  assign dispatch_pkt_o_348_ = expected_npc_i[25];
  assign dispatch_pkt_o[348] = dispatch_pkt_o_348_;
  assign dispatch_pkt_o_347_ = expected_npc_i[24];
  assign dispatch_pkt_o[347] = dispatch_pkt_o_347_;
  assign dispatch_pkt_o_346_ = expected_npc_i[23];
  assign dispatch_pkt_o[346] = dispatch_pkt_o_346_;
  assign dispatch_pkt_o_345_ = expected_npc_i[22];
  assign dispatch_pkt_o[345] = dispatch_pkt_o_345_;
  assign dispatch_pkt_o_344_ = expected_npc_i[21];
  assign dispatch_pkt_o[344] = dispatch_pkt_o_344_;
  assign dispatch_pkt_o_343_ = expected_npc_i[20];
  assign dispatch_pkt_o[343] = dispatch_pkt_o_343_;
  assign dispatch_pkt_o_342_ = expected_npc_i[19];
  assign dispatch_pkt_o[342] = dispatch_pkt_o_342_;
  assign dispatch_pkt_o_341_ = expected_npc_i[18];
  assign dispatch_pkt_o[341] = dispatch_pkt_o_341_;
  assign dispatch_pkt_o_340_ = expected_npc_i[17];
  assign dispatch_pkt_o[340] = dispatch_pkt_o_340_;
  assign dispatch_pkt_o_339_ = expected_npc_i[16];
  assign dispatch_pkt_o[339] = dispatch_pkt_o_339_;
  assign dispatch_pkt_o_338_ = expected_npc_i[15];
  assign dispatch_pkt_o[338] = dispatch_pkt_o_338_;
  assign dispatch_pkt_o_337_ = expected_npc_i[14];
  assign dispatch_pkt_o[337] = dispatch_pkt_o_337_;
  assign dispatch_pkt_o_336_ = expected_npc_i[13];
  assign dispatch_pkt_o[336] = dispatch_pkt_o_336_;
  assign dispatch_pkt_o_335_ = expected_npc_i[12];
  assign dispatch_pkt_o[335] = dispatch_pkt_o_335_;
  assign dispatch_pkt_o_334_ = expected_npc_i[11];
  assign dispatch_pkt_o[334] = dispatch_pkt_o_334_;
  assign dispatch_pkt_o_333_ = expected_npc_i[10];
  assign dispatch_pkt_o[333] = dispatch_pkt_o_333_;
  assign dispatch_pkt_o_332_ = expected_npc_i[9];
  assign dispatch_pkt_o[332] = dispatch_pkt_o_332_;
  assign dispatch_pkt_o_331_ = expected_npc_i[8];
  assign dispatch_pkt_o[331] = dispatch_pkt_o_331_;
  assign dispatch_pkt_o_330_ = expected_npc_i[7];
  assign dispatch_pkt_o[330] = dispatch_pkt_o_330_;
  assign dispatch_pkt_o_329_ = expected_npc_i[6];
  assign dispatch_pkt_o[329] = dispatch_pkt_o_329_;
  assign dispatch_pkt_o_328_ = expected_npc_i[5];
  assign dispatch_pkt_o[328] = dispatch_pkt_o_328_;
  assign dispatch_pkt_o_327_ = expected_npc_i[4];
  assign dispatch_pkt_o[327] = dispatch_pkt_o_327_;
  assign dispatch_pkt_o_326_ = expected_npc_i[3];
  assign dispatch_pkt_o[326] = dispatch_pkt_o_326_;
  assign dispatch_pkt_o_325_ = expected_npc_i[2];
  assign dispatch_pkt_o[325] = dispatch_pkt_o_325_;
  assign dispatch_pkt_o_324_ = expected_npc_i[1];
  assign dispatch_pkt_o[324] = dispatch_pkt_o_324_;
  assign dispatch_pkt_o_323_ = expected_npc_i[0];
  assign dispatch_pkt_o[323] = dispatch_pkt_o_323_;

  bp_be_ptw_00_64_3_8_9
  ptw
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .busy_o(ptw_busy_lo),
    .commit_pkt_i(commit_pkt_i),
    .trans_info_i(trans_info_i),
    .ordered_i(ordered_v_i),
    .v_o(ptw_v_lo),
    .walk_o(walk_decode_li_pipe_mem_final_v_),
    .itlb_fill_o(ptw_itlb_fill_lo),
    .dtlb_fill_o(ptw_dtlb_fill_lo),
    .instr_page_fault_o(ptw_instr_page_fault_lo),
    .load_page_fault_o(ptw_load_page_fault_lo),
    .store_page_fault_o(ptw_store_page_fault_lo),
    .count_o(ptw_count_lo),
    .addr_o(ptw_addr_lo),
    .pte_o(ptw_pte_lo),
    .v_i(ptw_v_li),
    .data_i(late_wb_pkt_i[68:5])
  );


  bp_be_issue_queue_00
  issue_queue
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(fe_queue_en_li),
    .clr_i(clear_iss_i),
    .roll_i(commit_pkt_i[213]),
    .read_i(fe_queue_read_li),
    .read_cnt_i({ 1'b0, issue_pkt_o[173:171] }),
    .read_size_i({ 1'b0, 1'b0, issue_pkt_o[170:169] }),
    .cmt_i(commit_pkt_i[211]),
    .cmt_cnt_i({ 1'b0, commit_pkt_i[210:208] }),
    .cmt_size_i({ 1'b0, 1'b0, commit_pkt_i[207:206] }),
    .fe_queue_i(fe_queue_i),
    .fe_queue_v_i(fe_queue_v_i),
    .fe_queue_ready_and_o(fe_queue_ready_and_o),
    .decode_info_i(decode_info_i),
    .preissue_pkt_o(preissue_pkt),
    .issue_pkt_o(issue_pkt_o)
  );


  bp_be_int_regfile_00
  int_regfile
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .rs_r_v_i({ preissue_pkt[37:37], preissue_pkt[38:38] }),
    .rs_addr_i(preissue_pkt[26:17]),
    .rs_data_o({ irf_rs2, irf_rs1 }),
    .rd_w_v_i(iwb_pkt_i[78]),
    .rd_addr_i(iwb_pkt_i[75:71]),
    .rd_data_i(iwb_pkt_i[70:5])
  );


  bp_be_fp_regfile_00
  fp_regfile
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .rs_r_v_i({ preissue_pkt[34:34], preissue_pkt[35:35], preissue_pkt[36:36] }),
    .rs_addr_i({ preissue_pkt[33:29], preissue_pkt[26:17] }),
    .rs_data_o({ frf_rs3, frf_rs2, frf_rs1 }),
    .rd_w_v_i(fwb_pkt_i[77]),
    .rd_addr_i(fwb_pkt_i[75:71]),
    .rd_data_i(fwb_pkt_i[70:5])
  );

  assign fe_exc_vaddr_li = issue_pkt_o[244:206] + { issue_pkt_o[173:171], 1'b0 };
  assign be_exc_vaddr_li = (N0)? ptw_addr_lo : 
                           (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = ptw_v_lo;
  assign be_exc_data_li = (N0)? { 1'b0, 1'b0, ptw_pte_lo } : 
                          (N8)? late_wb_pkt_i[70:5] : 
                          (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign be_exc_imm_li = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N11)? late_wb_pkt_i[4:0] : 
                         (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { be_exc_decode_li_pipe_mem_final_v_, be_exc_decode_li_irf_w_v_, be_exc_decode_li_frf_w_v_, be_exc_decode_li_dcache_mmu_v_, be_exc_decode_li_fu_op__t__5_, be_exc_decode_li_fu_op__t__4_, be_exc_decode_li_fu_op__t__3_ } = (N0)? { walk_decode_li_pipe_mem_final_v_, 1'b0, 1'b0, walk_decode_li_pipe_mem_final_v_, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                                                     (N14)? { 1'b0, late_wb_pkt_i[78:77], 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                     (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign be_exc_instr_li = (N0)? issue_pkt_o[205:174] : 
                           (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, late_wb_pkt_i[75:71], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign be_exc_count_li = (N0)? ptw_count_lo : 
                           (N20)? { 1'b0, 1'b0, 1'b0 } : 
                           (N19)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign dispatch_pkt_o[322:291] = (N1)? be_exc_instr_li : 
                                   (N40)? issue_pkt_o[205:174] : 
                                   (N22)? issue_pkt_o[205:174] : 1'b0;
  assign N1 = be_exc_not_instr_li;
  assign dispatch_pkt_o[287:286] = (N1)? { 1'b0, 1'b0 } : 
                                   (N41)? issue_pkt_o[170:169] : 
                                   (N24)? issue_pkt_o[170:169] : 1'b0;
  assign dispatch_pkt_o[290:288] = (N1)? be_exc_count_li : 
                                   (N42)? issue_pkt_o[173:171] : 
                                   (N26)? issue_pkt_o[173:171] : 1'b0;
  assign dispatch_pkt_o[231:166] = (N1)? { 1'b0, 1'b0, be_exc_vaddr_li } : 
                                   (N43)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fe_exc_vaddr_li } : 
                                   (N46)? frf_rs1 : 
                                   (N29)? irf_rs1 : 1'b0;
  assign dispatch_pkt_o[165:100] = (N1)? be_exc_data_li : 
                                   (N47)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N49)? frf_rs2 : 
                                   (N32)? irf_rs2 : 1'b0;
  assign dispatch_pkt_o[99:34] = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, be_exc_imm_li } : 
                                 (N50)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N52)? frf_rs3 : 
                                 (N35)? issue_pkt_o[114:49] : 1'b0;
  assign dispatch_pkt_o[285:232] = (N1)? { 1'b0, 1'b0, 1'b0, be_exc_decode_li_pipe_mem_final_v_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, be_exc_decode_li_irf_w_v_, be_exc_decode_li_frf_w_v_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, be_exc_decode_li_dcache_mmu_v_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, be_exc_decode_li_fu_op__t__5_, be_exc_decode_li_fu_op__t__4_, be_exc_decode_li_fu_op__t__3_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N53)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N37)? issue_pkt_o[168:115] : 1'b0;
  assign ptw_v_li = late_wb_yumi_o & late_wb_pkt_i[76];
  assign late_wb_yumi_o = late_wb_v_i & N55;
  assign N55 = late_wb_force_i | N54;
  assign N54 = ~issue_pkt_o[263];
  assign resume_v = N58 & resume_i;
  assign N58 = N56 & N57;
  assign N56 = ~late_wb_yumi_o;
  assign N57 = ~ptw_busy_lo;
  assign interrupt_v = N61 & irq_pending_i;
  assign N61 = N59 & N60;
  assign N59 = N56 & N57;
  assign N60 = ~resume_i;
  assign be_exc_not_instr_li = N63 | interrupt_v;
  assign N63 = N62 | resume_v;
  assign N62 = ptw_v_lo | late_wb_yumi_o;
  assign fe_exc_not_instr_li = N65 & N66;
  assign N65 = N64 & issue_pkt_o[263];
  assign N64 = ~be_exc_not_instr_li;
  assign N66 = ~issue_pkt_o[262];
  assign fe_instr_not_exc_li = N67 & issue_pkt_o[262];
  assign N67 = N64 & issue_pkt_o[263];
  assign fe_queue_en_li = N69 & N70;
  assign N69 = N68 & N57;
  assign N68 = ~suppress_iss_i;
  assign N70 = ~hazard_v_i;
  assign fe_queue_read_li = fe_instr_not_exc_li | fe_exc_not_instr_li;
  assign N2 = late_wb_yumi_o | ptw_v_lo;
  assign N3 = ~N2;
  assign N4 = ~ptw_v_lo;
  assign N5 = late_wb_yumi_o & N4;
  assign N6 = late_wb_yumi_o | ptw_v_lo;
  assign N7 = ~N6;
  assign N8 = late_wb_yumi_o & N4;
  assign N9 = late_wb_yumi_o | ptw_v_lo;
  assign N10 = ~N9;
  assign N11 = late_wb_yumi_o & N4;
  assign N12 = late_wb_yumi_o | ptw_v_lo;
  assign N13 = ~N12;
  assign N14 = late_wb_yumi_o & N4;
  assign N15 = late_wb_yumi_o | ptw_v_lo;
  assign N16 = ~N15;
  assign N17 = late_wb_yumi_o & N4;
  assign N18 = late_wb_yumi_o | ptw_v_lo;
  assign N19 = ~N18;
  assign N20 = late_wb_yumi_o & N4;
  assign dispatch_pkt_o[365] = N72 | be_exc_not_instr_li;
  assign N72 = fe_queue_read_li & N71;
  assign N71 = ~poison_isd_i;
  assign dispatch_pkt_o[364] = fe_queue_read_li & N71;
  assign dispatch_pkt_o[363] = fe_instr_not_exc_li & ispec_v_i;
  assign dispatch_pkt_o[362] = ptw_v_lo | late_wb_yumi_o;
  assign N21 = fe_exc_not_instr_li | be_exc_not_instr_li;
  assign N22 = ~N21;
  assign N23 = fe_exc_not_instr_li | be_exc_not_instr_li;
  assign N24 = ~N23;
  assign N25 = fe_exc_not_instr_li | be_exc_not_instr_li;
  assign N26 = ~N25;
  assign N27 = fe_exc_not_instr_li | be_exc_not_instr_li;
  assign N28 = issue_pkt_o[158] | N27;
  assign N29 = ~N28;
  assign N30 = fe_exc_not_instr_li | be_exc_not_instr_li;
  assign N31 = issue_pkt_o[157] | N30;
  assign N32 = ~N31;
  assign N33 = fe_exc_not_instr_li | be_exc_not_instr_li;
  assign N34 = issue_pkt_o[156] | N33;
  assign N35 = ~N34;
  assign N36 = fe_exc_not_instr_li | be_exc_not_instr_li;
  assign N37 = ~N36;
  assign N38 = be_exc_not_instr_li & ptw_instr_page_fault_lo;
  assign dispatch_pkt_o[32] = be_exc_not_instr_li & ptw_load_page_fault_lo;
  assign dispatch_pkt_o[33] = be_exc_not_instr_li & ptw_store_page_fault_lo;
  assign dispatch_pkt_o[13] = be_exc_not_instr_li & ptw_itlb_fill_lo;
  assign dispatch_pkt_o[12] = be_exc_not_instr_li & ptw_dtlb_fill_lo;
  assign dispatch_pkt_o[19] = be_exc_not_instr_li & resume_v;
  assign dispatch_pkt_o[11] = be_exc_not_instr_li & interrupt_v;
  assign dispatch_pkt_o[21] = fe_exc_not_instr_li & issue_pkt_o[260];
  assign dispatch_pkt_o[31] = N38 | N73;
  assign N73 = fe_exc_not_instr_li & issue_pkt_o[259];
  assign dispatch_pkt_o[18] = fe_exc_not_instr_li & issue_pkt_o[261];
  assign dispatch_pkt_o[17] = fe_exc_not_instr_li & issue_pkt_o[258];
  assign dispatch_pkt_o[22] = fe_exc_not_instr_li & issue_pkt_o[257];
  assign dispatch_pkt_o[30] = fe_instr_not_exc_li & issue_pkt_o[256];
  assign dispatch_pkt_o[29] = fe_instr_not_exc_li & issue_pkt_o[255];
  assign dispatch_pkt_o[28] = fe_instr_not_exc_li & issue_pkt_o[254];
  assign dispatch_pkt_o[23] = fe_instr_not_exc_li & issue_pkt_o[253];
  assign dispatch_pkt_o[5] = fe_instr_not_exc_li & issue_pkt_o[252];
  assign dispatch_pkt_o[4] = fe_instr_not_exc_li & issue_pkt_o[251];
  assign dispatch_pkt_o[3] = fe_instr_not_exc_li & issue_pkt_o[250];
  assign dispatch_pkt_o[2] = fe_instr_not_exc_li & issue_pkt_o[249];
  assign dispatch_pkt_o[1] = fe_instr_not_exc_li & issue_pkt_o[248];
  assign dispatch_pkt_o[6] = fe_instr_not_exc_li & issue_pkt_o[247];
  assign dispatch_pkt_o[7] = fe_instr_not_exc_li & issue_pkt_o[246];
  assign dispatch_pkt_o[0] = fe_instr_not_exc_li & issue_pkt_o[245];
  assign N39 = ~be_exc_not_instr_li;
  assign N40 = fe_exc_not_instr_li & N39;
  assign N41 = fe_exc_not_instr_li & N39;
  assign N42 = fe_exc_not_instr_li & N39;
  assign N43 = fe_exc_not_instr_li & N39;
  assign N44 = ~fe_exc_not_instr_li;
  assign N45 = N39 & N44;
  assign N46 = issue_pkt_o[158] & N45;
  assign N47 = fe_exc_not_instr_li & N39;
  assign N48 = N39 & N44;
  assign N49 = issue_pkt_o[157] & N48;
  assign N50 = fe_exc_not_instr_li & N39;
  assign N51 = N39 & N44;
  assign N52 = issue_pkt_o[156] & N51;
  assign N53 = fe_exc_not_instr_li & N39;

endmodule



module bsg_scan_width_p6_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [5:0] i;
  output [5:0] o;
  wire [5:0] o;
  wire t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,
  t_1__1_,t_1__0_;
  assign t_1__5_ = i[0] | 1'b0;
  assign t_1__4_ = i[1] | i[0];
  assign t_1__3_ = i[2] | i[1];
  assign t_1__2_ = i[3] | i[2];
  assign t_1__1_ = i[4] | i[3];
  assign t_1__0_ = i[5] | i[4];
  assign t_2__5_ = t_1__5_ | 1'b0;
  assign t_2__4_ = t_1__4_ | 1'b0;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign o[0] = t_2__5_ | 1'b0;
  assign o[1] = t_2__4_ | 1'b0;
  assign o[2] = t_2__3_ | 1'b0;
  assign o[3] = t_2__2_ | 1'b0;
  assign o[4] = t_2__1_ | t_2__5_;
  assign o[5] = t_2__0_ | t_2__4_;

endmodule



module bsg_priority_encode_one_hot_out_width_p6_lo_to_hi_p1
(
  i,
  o,
  v_o
);

  input [5:0] i;
  output [5:0] o;
  output v_o;
  wire [5:0] o;
  wire v_o,N0,N1,N2,N3,N4;
  wire [4:1] scan_lo;

  bsg_scan_width_p6_or_p1_lo_to_hi_p1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, scan_lo, o[0:0] })
  );

  assign o[5] = v_o & N0;
  assign N0 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N1;
  assign N1 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N2;
  assign N2 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N3;
  assign N3 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N4;
  assign N4 = ~o[0];

endmodule



module bsg_mux_one_hot_width_p66_els_p6
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [395:0] data_i;
  input [5:0] sel_one_hot_i;
  output [65:0] data_o;
  wire [65:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263;
  wire [395:0] data_masked;
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[1];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[1];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[1];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[1];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[1];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[1];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[1];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[2];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[2];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[2];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[2];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[2];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[2];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[2];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[2];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[2];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[2];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[2];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[2];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[2];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[2];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[2];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[2];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[2];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[2];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[2];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[2];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[2];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[2];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[2];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[2];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[2];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[2];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[2];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[2];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[2];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[2];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[2];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[2];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[2];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[2];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[2];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[2];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[2];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[2];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[2];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[2];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[2];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[2];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[2];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[2];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[2];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[2];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[2];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[2];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[2];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[2];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[2];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[2];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[2];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[2];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[2];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[2];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[2];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[2];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[2];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[2];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[2];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[2];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[2];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[2];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[2];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[2];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[3];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[3];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[3];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[3];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[3];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[3];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[3];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[3];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[3];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[3];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[3];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[3];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[3];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[3];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[3];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[3];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[3];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[3];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[3];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[3];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[3];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[3];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[3];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[3];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[3];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[3];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[3];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[3];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[3];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[3];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[3];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[3];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[3];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[3];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[3];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[3];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[3];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[3];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[3];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[3];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[3];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[3];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[3];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[3];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[3];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[3];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[3];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[3];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[3];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[3];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[3];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[3];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[3];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[3];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[3];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[3];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[3];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[3];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[3];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[3];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[3];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[3];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[3];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[3];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[3];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[3];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[4];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[4];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[4];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[4];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[4];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[4];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[4];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[4];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[4];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[4];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[4];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[4];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[4];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[4];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[4];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[4];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[4];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[4];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[4];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[4];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[4];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[4];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[4];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[4];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[4];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[4];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[4];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[4];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[4];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[4];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[4];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[4];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[4];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[4];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[4];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[4];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[4];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[4];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[4];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[4];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[4];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[4];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[4];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[4];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[4];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[4];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[4];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[4];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[4];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[4];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[4];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[4];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[4];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[4];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[4];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[4];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[4];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[4];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[4];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[4];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[4];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[4];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[4];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[4];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[4];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[4];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[5];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[5];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[5];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[5];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[5];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[5];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[5];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[5];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[5];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[5];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[5];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[5];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[5];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[5];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[5];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[5];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[5];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[5];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[5];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[5];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[5];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[5];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[5];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[5];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[5];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[5];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[5];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[5];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[5];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[5];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[5];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[5];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[5];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[5];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[5];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[5];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[5];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[5];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[5];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[5];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[5];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[5];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[5];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[5];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[5];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[5];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[5];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[5];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[5];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[5];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[5];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[5];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[5];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[5];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[5];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[5];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[5];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[5];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[5];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[5];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[5];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[5];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[5];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[5];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[5];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[5];
  assign data_o[0] = N3 | data_masked[0];
  assign N3 = N2 | data_masked[66];
  assign N2 = N1 | data_masked[132];
  assign N1 = N0 | data_masked[198];
  assign N0 = data_masked[330] | data_masked[264];
  assign data_o[1] = N7 | data_masked[1];
  assign N7 = N6 | data_masked[67];
  assign N6 = N5 | data_masked[133];
  assign N5 = N4 | data_masked[199];
  assign N4 = data_masked[331] | data_masked[265];
  assign data_o[2] = N11 | data_masked[2];
  assign N11 = N10 | data_masked[68];
  assign N10 = N9 | data_masked[134];
  assign N9 = N8 | data_masked[200];
  assign N8 = data_masked[332] | data_masked[266];
  assign data_o[3] = N15 | data_masked[3];
  assign N15 = N14 | data_masked[69];
  assign N14 = N13 | data_masked[135];
  assign N13 = N12 | data_masked[201];
  assign N12 = data_masked[333] | data_masked[267];
  assign data_o[4] = N19 | data_masked[4];
  assign N19 = N18 | data_masked[70];
  assign N18 = N17 | data_masked[136];
  assign N17 = N16 | data_masked[202];
  assign N16 = data_masked[334] | data_masked[268];
  assign data_o[5] = N23 | data_masked[5];
  assign N23 = N22 | data_masked[71];
  assign N22 = N21 | data_masked[137];
  assign N21 = N20 | data_masked[203];
  assign N20 = data_masked[335] | data_masked[269];
  assign data_o[6] = N27 | data_masked[6];
  assign N27 = N26 | data_masked[72];
  assign N26 = N25 | data_masked[138];
  assign N25 = N24 | data_masked[204];
  assign N24 = data_masked[336] | data_masked[270];
  assign data_o[7] = N31 | data_masked[7];
  assign N31 = N30 | data_masked[73];
  assign N30 = N29 | data_masked[139];
  assign N29 = N28 | data_masked[205];
  assign N28 = data_masked[337] | data_masked[271];
  assign data_o[8] = N35 | data_masked[8];
  assign N35 = N34 | data_masked[74];
  assign N34 = N33 | data_masked[140];
  assign N33 = N32 | data_masked[206];
  assign N32 = data_masked[338] | data_masked[272];
  assign data_o[9] = N39 | data_masked[9];
  assign N39 = N38 | data_masked[75];
  assign N38 = N37 | data_masked[141];
  assign N37 = N36 | data_masked[207];
  assign N36 = data_masked[339] | data_masked[273];
  assign data_o[10] = N43 | data_masked[10];
  assign N43 = N42 | data_masked[76];
  assign N42 = N41 | data_masked[142];
  assign N41 = N40 | data_masked[208];
  assign N40 = data_masked[340] | data_masked[274];
  assign data_o[11] = N47 | data_masked[11];
  assign N47 = N46 | data_masked[77];
  assign N46 = N45 | data_masked[143];
  assign N45 = N44 | data_masked[209];
  assign N44 = data_masked[341] | data_masked[275];
  assign data_o[12] = N51 | data_masked[12];
  assign N51 = N50 | data_masked[78];
  assign N50 = N49 | data_masked[144];
  assign N49 = N48 | data_masked[210];
  assign N48 = data_masked[342] | data_masked[276];
  assign data_o[13] = N55 | data_masked[13];
  assign N55 = N54 | data_masked[79];
  assign N54 = N53 | data_masked[145];
  assign N53 = N52 | data_masked[211];
  assign N52 = data_masked[343] | data_masked[277];
  assign data_o[14] = N59 | data_masked[14];
  assign N59 = N58 | data_masked[80];
  assign N58 = N57 | data_masked[146];
  assign N57 = N56 | data_masked[212];
  assign N56 = data_masked[344] | data_masked[278];
  assign data_o[15] = N63 | data_masked[15];
  assign N63 = N62 | data_masked[81];
  assign N62 = N61 | data_masked[147];
  assign N61 = N60 | data_masked[213];
  assign N60 = data_masked[345] | data_masked[279];
  assign data_o[16] = N67 | data_masked[16];
  assign N67 = N66 | data_masked[82];
  assign N66 = N65 | data_masked[148];
  assign N65 = N64 | data_masked[214];
  assign N64 = data_masked[346] | data_masked[280];
  assign data_o[17] = N71 | data_masked[17];
  assign N71 = N70 | data_masked[83];
  assign N70 = N69 | data_masked[149];
  assign N69 = N68 | data_masked[215];
  assign N68 = data_masked[347] | data_masked[281];
  assign data_o[18] = N75 | data_masked[18];
  assign N75 = N74 | data_masked[84];
  assign N74 = N73 | data_masked[150];
  assign N73 = N72 | data_masked[216];
  assign N72 = data_masked[348] | data_masked[282];
  assign data_o[19] = N79 | data_masked[19];
  assign N79 = N78 | data_masked[85];
  assign N78 = N77 | data_masked[151];
  assign N77 = N76 | data_masked[217];
  assign N76 = data_masked[349] | data_masked[283];
  assign data_o[20] = N83 | data_masked[20];
  assign N83 = N82 | data_masked[86];
  assign N82 = N81 | data_masked[152];
  assign N81 = N80 | data_masked[218];
  assign N80 = data_masked[350] | data_masked[284];
  assign data_o[21] = N87 | data_masked[21];
  assign N87 = N86 | data_masked[87];
  assign N86 = N85 | data_masked[153];
  assign N85 = N84 | data_masked[219];
  assign N84 = data_masked[351] | data_masked[285];
  assign data_o[22] = N91 | data_masked[22];
  assign N91 = N90 | data_masked[88];
  assign N90 = N89 | data_masked[154];
  assign N89 = N88 | data_masked[220];
  assign N88 = data_masked[352] | data_masked[286];
  assign data_o[23] = N95 | data_masked[23];
  assign N95 = N94 | data_masked[89];
  assign N94 = N93 | data_masked[155];
  assign N93 = N92 | data_masked[221];
  assign N92 = data_masked[353] | data_masked[287];
  assign data_o[24] = N99 | data_masked[24];
  assign N99 = N98 | data_masked[90];
  assign N98 = N97 | data_masked[156];
  assign N97 = N96 | data_masked[222];
  assign N96 = data_masked[354] | data_masked[288];
  assign data_o[25] = N103 | data_masked[25];
  assign N103 = N102 | data_masked[91];
  assign N102 = N101 | data_masked[157];
  assign N101 = N100 | data_masked[223];
  assign N100 = data_masked[355] | data_masked[289];
  assign data_o[26] = N107 | data_masked[26];
  assign N107 = N106 | data_masked[92];
  assign N106 = N105 | data_masked[158];
  assign N105 = N104 | data_masked[224];
  assign N104 = data_masked[356] | data_masked[290];
  assign data_o[27] = N111 | data_masked[27];
  assign N111 = N110 | data_masked[93];
  assign N110 = N109 | data_masked[159];
  assign N109 = N108 | data_masked[225];
  assign N108 = data_masked[357] | data_masked[291];
  assign data_o[28] = N115 | data_masked[28];
  assign N115 = N114 | data_masked[94];
  assign N114 = N113 | data_masked[160];
  assign N113 = N112 | data_masked[226];
  assign N112 = data_masked[358] | data_masked[292];
  assign data_o[29] = N119 | data_masked[29];
  assign N119 = N118 | data_masked[95];
  assign N118 = N117 | data_masked[161];
  assign N117 = N116 | data_masked[227];
  assign N116 = data_masked[359] | data_masked[293];
  assign data_o[30] = N123 | data_masked[30];
  assign N123 = N122 | data_masked[96];
  assign N122 = N121 | data_masked[162];
  assign N121 = N120 | data_masked[228];
  assign N120 = data_masked[360] | data_masked[294];
  assign data_o[31] = N127 | data_masked[31];
  assign N127 = N126 | data_masked[97];
  assign N126 = N125 | data_masked[163];
  assign N125 = N124 | data_masked[229];
  assign N124 = data_masked[361] | data_masked[295];
  assign data_o[32] = N131 | data_masked[32];
  assign N131 = N130 | data_masked[98];
  assign N130 = N129 | data_masked[164];
  assign N129 = N128 | data_masked[230];
  assign N128 = data_masked[362] | data_masked[296];
  assign data_o[33] = N135 | data_masked[33];
  assign N135 = N134 | data_masked[99];
  assign N134 = N133 | data_masked[165];
  assign N133 = N132 | data_masked[231];
  assign N132 = data_masked[363] | data_masked[297];
  assign data_o[34] = N139 | data_masked[34];
  assign N139 = N138 | data_masked[100];
  assign N138 = N137 | data_masked[166];
  assign N137 = N136 | data_masked[232];
  assign N136 = data_masked[364] | data_masked[298];
  assign data_o[35] = N143 | data_masked[35];
  assign N143 = N142 | data_masked[101];
  assign N142 = N141 | data_masked[167];
  assign N141 = N140 | data_masked[233];
  assign N140 = data_masked[365] | data_masked[299];
  assign data_o[36] = N147 | data_masked[36];
  assign N147 = N146 | data_masked[102];
  assign N146 = N145 | data_masked[168];
  assign N145 = N144 | data_masked[234];
  assign N144 = data_masked[366] | data_masked[300];
  assign data_o[37] = N151 | data_masked[37];
  assign N151 = N150 | data_masked[103];
  assign N150 = N149 | data_masked[169];
  assign N149 = N148 | data_masked[235];
  assign N148 = data_masked[367] | data_masked[301];
  assign data_o[38] = N155 | data_masked[38];
  assign N155 = N154 | data_masked[104];
  assign N154 = N153 | data_masked[170];
  assign N153 = N152 | data_masked[236];
  assign N152 = data_masked[368] | data_masked[302];
  assign data_o[39] = N159 | data_masked[39];
  assign N159 = N158 | data_masked[105];
  assign N158 = N157 | data_masked[171];
  assign N157 = N156 | data_masked[237];
  assign N156 = data_masked[369] | data_masked[303];
  assign data_o[40] = N163 | data_masked[40];
  assign N163 = N162 | data_masked[106];
  assign N162 = N161 | data_masked[172];
  assign N161 = N160 | data_masked[238];
  assign N160 = data_masked[370] | data_masked[304];
  assign data_o[41] = N167 | data_masked[41];
  assign N167 = N166 | data_masked[107];
  assign N166 = N165 | data_masked[173];
  assign N165 = N164 | data_masked[239];
  assign N164 = data_masked[371] | data_masked[305];
  assign data_o[42] = N171 | data_masked[42];
  assign N171 = N170 | data_masked[108];
  assign N170 = N169 | data_masked[174];
  assign N169 = N168 | data_masked[240];
  assign N168 = data_masked[372] | data_masked[306];
  assign data_o[43] = N175 | data_masked[43];
  assign N175 = N174 | data_masked[109];
  assign N174 = N173 | data_masked[175];
  assign N173 = N172 | data_masked[241];
  assign N172 = data_masked[373] | data_masked[307];
  assign data_o[44] = N179 | data_masked[44];
  assign N179 = N178 | data_masked[110];
  assign N178 = N177 | data_masked[176];
  assign N177 = N176 | data_masked[242];
  assign N176 = data_masked[374] | data_masked[308];
  assign data_o[45] = N183 | data_masked[45];
  assign N183 = N182 | data_masked[111];
  assign N182 = N181 | data_masked[177];
  assign N181 = N180 | data_masked[243];
  assign N180 = data_masked[375] | data_masked[309];
  assign data_o[46] = N187 | data_masked[46];
  assign N187 = N186 | data_masked[112];
  assign N186 = N185 | data_masked[178];
  assign N185 = N184 | data_masked[244];
  assign N184 = data_masked[376] | data_masked[310];
  assign data_o[47] = N191 | data_masked[47];
  assign N191 = N190 | data_masked[113];
  assign N190 = N189 | data_masked[179];
  assign N189 = N188 | data_masked[245];
  assign N188 = data_masked[377] | data_masked[311];
  assign data_o[48] = N195 | data_masked[48];
  assign N195 = N194 | data_masked[114];
  assign N194 = N193 | data_masked[180];
  assign N193 = N192 | data_masked[246];
  assign N192 = data_masked[378] | data_masked[312];
  assign data_o[49] = N199 | data_masked[49];
  assign N199 = N198 | data_masked[115];
  assign N198 = N197 | data_masked[181];
  assign N197 = N196 | data_masked[247];
  assign N196 = data_masked[379] | data_masked[313];
  assign data_o[50] = N203 | data_masked[50];
  assign N203 = N202 | data_masked[116];
  assign N202 = N201 | data_masked[182];
  assign N201 = N200 | data_masked[248];
  assign N200 = data_masked[380] | data_masked[314];
  assign data_o[51] = N207 | data_masked[51];
  assign N207 = N206 | data_masked[117];
  assign N206 = N205 | data_masked[183];
  assign N205 = N204 | data_masked[249];
  assign N204 = data_masked[381] | data_masked[315];
  assign data_o[52] = N211 | data_masked[52];
  assign N211 = N210 | data_masked[118];
  assign N210 = N209 | data_masked[184];
  assign N209 = N208 | data_masked[250];
  assign N208 = data_masked[382] | data_masked[316];
  assign data_o[53] = N215 | data_masked[53];
  assign N215 = N214 | data_masked[119];
  assign N214 = N213 | data_masked[185];
  assign N213 = N212 | data_masked[251];
  assign N212 = data_masked[383] | data_masked[317];
  assign data_o[54] = N219 | data_masked[54];
  assign N219 = N218 | data_masked[120];
  assign N218 = N217 | data_masked[186];
  assign N217 = N216 | data_masked[252];
  assign N216 = data_masked[384] | data_masked[318];
  assign data_o[55] = N223 | data_masked[55];
  assign N223 = N222 | data_masked[121];
  assign N222 = N221 | data_masked[187];
  assign N221 = N220 | data_masked[253];
  assign N220 = data_masked[385] | data_masked[319];
  assign data_o[56] = N227 | data_masked[56];
  assign N227 = N226 | data_masked[122];
  assign N226 = N225 | data_masked[188];
  assign N225 = N224 | data_masked[254];
  assign N224 = data_masked[386] | data_masked[320];
  assign data_o[57] = N231 | data_masked[57];
  assign N231 = N230 | data_masked[123];
  assign N230 = N229 | data_masked[189];
  assign N229 = N228 | data_masked[255];
  assign N228 = data_masked[387] | data_masked[321];
  assign data_o[58] = N235 | data_masked[58];
  assign N235 = N234 | data_masked[124];
  assign N234 = N233 | data_masked[190];
  assign N233 = N232 | data_masked[256];
  assign N232 = data_masked[388] | data_masked[322];
  assign data_o[59] = N239 | data_masked[59];
  assign N239 = N238 | data_masked[125];
  assign N238 = N237 | data_masked[191];
  assign N237 = N236 | data_masked[257];
  assign N236 = data_masked[389] | data_masked[323];
  assign data_o[60] = N243 | data_masked[60];
  assign N243 = N242 | data_masked[126];
  assign N242 = N241 | data_masked[192];
  assign N241 = N240 | data_masked[258];
  assign N240 = data_masked[390] | data_masked[324];
  assign data_o[61] = N247 | data_masked[61];
  assign N247 = N246 | data_masked[127];
  assign N246 = N245 | data_masked[193];
  assign N245 = N244 | data_masked[259];
  assign N244 = data_masked[391] | data_masked[325];
  assign data_o[62] = N251 | data_masked[62];
  assign N251 = N250 | data_masked[128];
  assign N250 = N249 | data_masked[194];
  assign N249 = N248 | data_masked[260];
  assign N248 = data_masked[392] | data_masked[326];
  assign data_o[63] = N255 | data_masked[63];
  assign N255 = N254 | data_masked[129];
  assign N254 = N253 | data_masked[195];
  assign N253 = N252 | data_masked[261];
  assign N252 = data_masked[393] | data_masked[327];
  assign data_o[64] = N259 | data_masked[64];
  assign N259 = N258 | data_masked[130];
  assign N258 = N257 | data_masked[196];
  assign N257 = N256 | data_masked[262];
  assign N256 = data_masked[394] | data_masked[328];
  assign data_o[65] = N263 | data_masked[65];
  assign N263 = N262 | data_masked[131];
  assign N262 = N261 | data_masked[197];
  assign N261 = N260 | data_masked[263];
  assign N260 = data_masked[395] | data_masked[329];

endmodule



module bsg_dff_0000016e
(
  clk_i,
  data_i,
  data_o
);

  input [365:0] data_i;
  output [365:0] data_o;
  input clk_i;
  wire [365:0] data_o;
  reg data_o_365_sv2v_reg,data_o_364_sv2v_reg,data_o_363_sv2v_reg,data_o_362_sv2v_reg,
  data_o_361_sv2v_reg,data_o_360_sv2v_reg,data_o_359_sv2v_reg,data_o_358_sv2v_reg,
  data_o_357_sv2v_reg,data_o_356_sv2v_reg,data_o_355_sv2v_reg,data_o_354_sv2v_reg,
  data_o_353_sv2v_reg,data_o_352_sv2v_reg,data_o_351_sv2v_reg,data_o_350_sv2v_reg,
  data_o_349_sv2v_reg,data_o_348_sv2v_reg,data_o_347_sv2v_reg,data_o_346_sv2v_reg,
  data_o_345_sv2v_reg,data_o_344_sv2v_reg,data_o_343_sv2v_reg,data_o_342_sv2v_reg,
  data_o_341_sv2v_reg,data_o_340_sv2v_reg,data_o_339_sv2v_reg,data_o_338_sv2v_reg,
  data_o_337_sv2v_reg,data_o_336_sv2v_reg,data_o_335_sv2v_reg,data_o_334_sv2v_reg,
  data_o_333_sv2v_reg,data_o_332_sv2v_reg,data_o_331_sv2v_reg,data_o_330_sv2v_reg,
  data_o_329_sv2v_reg,data_o_328_sv2v_reg,data_o_327_sv2v_reg,data_o_326_sv2v_reg,
  data_o_325_sv2v_reg,data_o_324_sv2v_reg,data_o_323_sv2v_reg,data_o_322_sv2v_reg,
  data_o_321_sv2v_reg,data_o_320_sv2v_reg,data_o_319_sv2v_reg,data_o_318_sv2v_reg,
  data_o_317_sv2v_reg,data_o_316_sv2v_reg,data_o_315_sv2v_reg,data_o_314_sv2v_reg,
  data_o_313_sv2v_reg,data_o_312_sv2v_reg,data_o_311_sv2v_reg,data_o_310_sv2v_reg,
  data_o_309_sv2v_reg,data_o_308_sv2v_reg,data_o_307_sv2v_reg,data_o_306_sv2v_reg,
  data_o_305_sv2v_reg,data_o_304_sv2v_reg,data_o_303_sv2v_reg,data_o_302_sv2v_reg,
  data_o_301_sv2v_reg,data_o_300_sv2v_reg,data_o_299_sv2v_reg,data_o_298_sv2v_reg,
  data_o_297_sv2v_reg,data_o_296_sv2v_reg,data_o_295_sv2v_reg,data_o_294_sv2v_reg,
  data_o_293_sv2v_reg,data_o_292_sv2v_reg,data_o_291_sv2v_reg,data_o_290_sv2v_reg,
  data_o_289_sv2v_reg,data_o_288_sv2v_reg,data_o_287_sv2v_reg,data_o_286_sv2v_reg,
  data_o_285_sv2v_reg,data_o_284_sv2v_reg,data_o_283_sv2v_reg,data_o_282_sv2v_reg,
  data_o_281_sv2v_reg,data_o_280_sv2v_reg,data_o_279_sv2v_reg,data_o_278_sv2v_reg,
  data_o_277_sv2v_reg,data_o_276_sv2v_reg,data_o_275_sv2v_reg,data_o_274_sv2v_reg,
  data_o_273_sv2v_reg,data_o_272_sv2v_reg,data_o_271_sv2v_reg,data_o_270_sv2v_reg,
  data_o_269_sv2v_reg,data_o_268_sv2v_reg,data_o_267_sv2v_reg,data_o_266_sv2v_reg,
  data_o_265_sv2v_reg,data_o_264_sv2v_reg,data_o_263_sv2v_reg,data_o_262_sv2v_reg,
  data_o_261_sv2v_reg,data_o_260_sv2v_reg,data_o_259_sv2v_reg,data_o_258_sv2v_reg,
  data_o_257_sv2v_reg,data_o_256_sv2v_reg,data_o_255_sv2v_reg,data_o_254_sv2v_reg,
  data_o_253_sv2v_reg,data_o_252_sv2v_reg,data_o_251_sv2v_reg,data_o_250_sv2v_reg,
  data_o_249_sv2v_reg,data_o_248_sv2v_reg,data_o_247_sv2v_reg,data_o_246_sv2v_reg,
  data_o_245_sv2v_reg,data_o_244_sv2v_reg,data_o_243_sv2v_reg,data_o_242_sv2v_reg,
  data_o_241_sv2v_reg,data_o_240_sv2v_reg,data_o_239_sv2v_reg,data_o_238_sv2v_reg,
  data_o_237_sv2v_reg,data_o_236_sv2v_reg,data_o_235_sv2v_reg,data_o_234_sv2v_reg,
  data_o_233_sv2v_reg,data_o_232_sv2v_reg,data_o_231_sv2v_reg,data_o_230_sv2v_reg,
  data_o_229_sv2v_reg,data_o_228_sv2v_reg,data_o_227_sv2v_reg,data_o_226_sv2v_reg,
  data_o_225_sv2v_reg,data_o_224_sv2v_reg,data_o_223_sv2v_reg,data_o_222_sv2v_reg,
  data_o_221_sv2v_reg,data_o_220_sv2v_reg,data_o_219_sv2v_reg,data_o_218_sv2v_reg,
  data_o_217_sv2v_reg,data_o_216_sv2v_reg,data_o_215_sv2v_reg,data_o_214_sv2v_reg,
  data_o_213_sv2v_reg,data_o_212_sv2v_reg,data_o_211_sv2v_reg,data_o_210_sv2v_reg,
  data_o_209_sv2v_reg,data_o_208_sv2v_reg,data_o_207_sv2v_reg,data_o_206_sv2v_reg,
  data_o_205_sv2v_reg,data_o_204_sv2v_reg,data_o_203_sv2v_reg,data_o_202_sv2v_reg,
  data_o_201_sv2v_reg,data_o_200_sv2v_reg,data_o_199_sv2v_reg,data_o_198_sv2v_reg,
  data_o_197_sv2v_reg,data_o_196_sv2v_reg,data_o_195_sv2v_reg,data_o_194_sv2v_reg,
  data_o_193_sv2v_reg,data_o_192_sv2v_reg,data_o_191_sv2v_reg,data_o_190_sv2v_reg,
  data_o_189_sv2v_reg,data_o_188_sv2v_reg,data_o_187_sv2v_reg,data_o_186_sv2v_reg,
  data_o_185_sv2v_reg,data_o_184_sv2v_reg,data_o_183_sv2v_reg,data_o_182_sv2v_reg,
  data_o_181_sv2v_reg,data_o_180_sv2v_reg,data_o_179_sv2v_reg,data_o_178_sv2v_reg,
  data_o_177_sv2v_reg,data_o_176_sv2v_reg,data_o_175_sv2v_reg,data_o_174_sv2v_reg,
  data_o_173_sv2v_reg,data_o_172_sv2v_reg,data_o_171_sv2v_reg,data_o_170_sv2v_reg,
  data_o_169_sv2v_reg,data_o_168_sv2v_reg,data_o_167_sv2v_reg,data_o_166_sv2v_reg,
  data_o_165_sv2v_reg,data_o_164_sv2v_reg,data_o_163_sv2v_reg,data_o_162_sv2v_reg,
  data_o_161_sv2v_reg,data_o_160_sv2v_reg,data_o_159_sv2v_reg,data_o_158_sv2v_reg,
  data_o_157_sv2v_reg,data_o_156_sv2v_reg,data_o_155_sv2v_reg,data_o_154_sv2v_reg,
  data_o_153_sv2v_reg,data_o_152_sv2v_reg,data_o_151_sv2v_reg,data_o_150_sv2v_reg,
  data_o_149_sv2v_reg,data_o_148_sv2v_reg,data_o_147_sv2v_reg,data_o_146_sv2v_reg,
  data_o_145_sv2v_reg,data_o_144_sv2v_reg,data_o_143_sv2v_reg,data_o_142_sv2v_reg,
  data_o_141_sv2v_reg,data_o_140_sv2v_reg,data_o_139_sv2v_reg,data_o_138_sv2v_reg,
  data_o_137_sv2v_reg,data_o_136_sv2v_reg,data_o_135_sv2v_reg,data_o_134_sv2v_reg,
  data_o_133_sv2v_reg,data_o_132_sv2v_reg,data_o_131_sv2v_reg,data_o_130_sv2v_reg,
  data_o_129_sv2v_reg,data_o_128_sv2v_reg,data_o_127_sv2v_reg,data_o_126_sv2v_reg,
  data_o_125_sv2v_reg,data_o_124_sv2v_reg,data_o_123_sv2v_reg,data_o_122_sv2v_reg,
  data_o_121_sv2v_reg,data_o_120_sv2v_reg,data_o_119_sv2v_reg,data_o_118_sv2v_reg,
  data_o_117_sv2v_reg,data_o_116_sv2v_reg,data_o_115_sv2v_reg,data_o_114_sv2v_reg,
  data_o_113_sv2v_reg,data_o_112_sv2v_reg,data_o_111_sv2v_reg,data_o_110_sv2v_reg,
  data_o_109_sv2v_reg,data_o_108_sv2v_reg,data_o_107_sv2v_reg,data_o_106_sv2v_reg,
  data_o_105_sv2v_reg,data_o_104_sv2v_reg,data_o_103_sv2v_reg,data_o_102_sv2v_reg,
  data_o_101_sv2v_reg,data_o_100_sv2v_reg,data_o_99_sv2v_reg,data_o_98_sv2v_reg,
  data_o_97_sv2v_reg,data_o_96_sv2v_reg,data_o_95_sv2v_reg,data_o_94_sv2v_reg,
  data_o_93_sv2v_reg,data_o_92_sv2v_reg,data_o_91_sv2v_reg,data_o_90_sv2v_reg,
  data_o_89_sv2v_reg,data_o_88_sv2v_reg,data_o_87_sv2v_reg,data_o_86_sv2v_reg,
  data_o_85_sv2v_reg,data_o_84_sv2v_reg,data_o_83_sv2v_reg,data_o_82_sv2v_reg,
  data_o_81_sv2v_reg,data_o_80_sv2v_reg,data_o_79_sv2v_reg,data_o_78_sv2v_reg,data_o_77_sv2v_reg,
  data_o_76_sv2v_reg,data_o_75_sv2v_reg,data_o_74_sv2v_reg,data_o_73_sv2v_reg,
  data_o_72_sv2v_reg,data_o_71_sv2v_reg,data_o_70_sv2v_reg,data_o_69_sv2v_reg,
  data_o_68_sv2v_reg,data_o_67_sv2v_reg,data_o_66_sv2v_reg,data_o_65_sv2v_reg,
  data_o_64_sv2v_reg,data_o_63_sv2v_reg,data_o_62_sv2v_reg,data_o_61_sv2v_reg,data_o_60_sv2v_reg,
  data_o_59_sv2v_reg,data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,
  data_o_55_sv2v_reg,data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,
  data_o_51_sv2v_reg,data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,
  data_o_47_sv2v_reg,data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,
  data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,
  data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,
  data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,
  data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,
  data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,
  data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,
  data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[365] = data_o_365_sv2v_reg;
  assign data_o[364] = data_o_364_sv2v_reg;
  assign data_o[363] = data_o_363_sv2v_reg;
  assign data_o[362] = data_o_362_sv2v_reg;
  assign data_o[361] = data_o_361_sv2v_reg;
  assign data_o[360] = data_o_360_sv2v_reg;
  assign data_o[359] = data_o_359_sv2v_reg;
  assign data_o[358] = data_o_358_sv2v_reg;
  assign data_o[357] = data_o_357_sv2v_reg;
  assign data_o[356] = data_o_356_sv2v_reg;
  assign data_o[355] = data_o_355_sv2v_reg;
  assign data_o[354] = data_o_354_sv2v_reg;
  assign data_o[353] = data_o_353_sv2v_reg;
  assign data_o[352] = data_o_352_sv2v_reg;
  assign data_o[351] = data_o_351_sv2v_reg;
  assign data_o[350] = data_o_350_sv2v_reg;
  assign data_o[349] = data_o_349_sv2v_reg;
  assign data_o[348] = data_o_348_sv2v_reg;
  assign data_o[347] = data_o_347_sv2v_reg;
  assign data_o[346] = data_o_346_sv2v_reg;
  assign data_o[345] = data_o_345_sv2v_reg;
  assign data_o[344] = data_o_344_sv2v_reg;
  assign data_o[343] = data_o_343_sv2v_reg;
  assign data_o[342] = data_o_342_sv2v_reg;
  assign data_o[341] = data_o_341_sv2v_reg;
  assign data_o[340] = data_o_340_sv2v_reg;
  assign data_o[339] = data_o_339_sv2v_reg;
  assign data_o[338] = data_o_338_sv2v_reg;
  assign data_o[337] = data_o_337_sv2v_reg;
  assign data_o[336] = data_o_336_sv2v_reg;
  assign data_o[335] = data_o_335_sv2v_reg;
  assign data_o[334] = data_o_334_sv2v_reg;
  assign data_o[333] = data_o_333_sv2v_reg;
  assign data_o[332] = data_o_332_sv2v_reg;
  assign data_o[331] = data_o_331_sv2v_reg;
  assign data_o[330] = data_o_330_sv2v_reg;
  assign data_o[329] = data_o_329_sv2v_reg;
  assign data_o[328] = data_o_328_sv2v_reg;
  assign data_o[327] = data_o_327_sv2v_reg;
  assign data_o[326] = data_o_326_sv2v_reg;
  assign data_o[325] = data_o_325_sv2v_reg;
  assign data_o[324] = data_o_324_sv2v_reg;
  assign data_o[323] = data_o_323_sv2v_reg;
  assign data_o[322] = data_o_322_sv2v_reg;
  assign data_o[321] = data_o_321_sv2v_reg;
  assign data_o[320] = data_o_320_sv2v_reg;
  assign data_o[319] = data_o_319_sv2v_reg;
  assign data_o[318] = data_o_318_sv2v_reg;
  assign data_o[317] = data_o_317_sv2v_reg;
  assign data_o[316] = data_o_316_sv2v_reg;
  assign data_o[315] = data_o_315_sv2v_reg;
  assign data_o[314] = data_o_314_sv2v_reg;
  assign data_o[313] = data_o_313_sv2v_reg;
  assign data_o[312] = data_o_312_sv2v_reg;
  assign data_o[311] = data_o_311_sv2v_reg;
  assign data_o[310] = data_o_310_sv2v_reg;
  assign data_o[309] = data_o_309_sv2v_reg;
  assign data_o[308] = data_o_308_sv2v_reg;
  assign data_o[307] = data_o_307_sv2v_reg;
  assign data_o[306] = data_o_306_sv2v_reg;
  assign data_o[305] = data_o_305_sv2v_reg;
  assign data_o[304] = data_o_304_sv2v_reg;
  assign data_o[303] = data_o_303_sv2v_reg;
  assign data_o[302] = data_o_302_sv2v_reg;
  assign data_o[301] = data_o_301_sv2v_reg;
  assign data_o[300] = data_o_300_sv2v_reg;
  assign data_o[299] = data_o_299_sv2v_reg;
  assign data_o[298] = data_o_298_sv2v_reg;
  assign data_o[297] = data_o_297_sv2v_reg;
  assign data_o[296] = data_o_296_sv2v_reg;
  assign data_o[295] = data_o_295_sv2v_reg;
  assign data_o[294] = data_o_294_sv2v_reg;
  assign data_o[293] = data_o_293_sv2v_reg;
  assign data_o[292] = data_o_292_sv2v_reg;
  assign data_o[291] = data_o_291_sv2v_reg;
  assign data_o[290] = data_o_290_sv2v_reg;
  assign data_o[289] = data_o_289_sv2v_reg;
  assign data_o[288] = data_o_288_sv2v_reg;
  assign data_o[287] = data_o_287_sv2v_reg;
  assign data_o[286] = data_o_286_sv2v_reg;
  assign data_o[285] = data_o_285_sv2v_reg;
  assign data_o[284] = data_o_284_sv2v_reg;
  assign data_o[283] = data_o_283_sv2v_reg;
  assign data_o[282] = data_o_282_sv2v_reg;
  assign data_o[281] = data_o_281_sv2v_reg;
  assign data_o[280] = data_o_280_sv2v_reg;
  assign data_o[279] = data_o_279_sv2v_reg;
  assign data_o[278] = data_o_278_sv2v_reg;
  assign data_o[277] = data_o_277_sv2v_reg;
  assign data_o[276] = data_o_276_sv2v_reg;
  assign data_o[275] = data_o_275_sv2v_reg;
  assign data_o[274] = data_o_274_sv2v_reg;
  assign data_o[273] = data_o_273_sv2v_reg;
  assign data_o[272] = data_o_272_sv2v_reg;
  assign data_o[271] = data_o_271_sv2v_reg;
  assign data_o[270] = data_o_270_sv2v_reg;
  assign data_o[269] = data_o_269_sv2v_reg;
  assign data_o[268] = data_o_268_sv2v_reg;
  assign data_o[267] = data_o_267_sv2v_reg;
  assign data_o[266] = data_o_266_sv2v_reg;
  assign data_o[265] = data_o_265_sv2v_reg;
  assign data_o[264] = data_o_264_sv2v_reg;
  assign data_o[263] = data_o_263_sv2v_reg;
  assign data_o[262] = data_o_262_sv2v_reg;
  assign data_o[261] = data_o_261_sv2v_reg;
  assign data_o[260] = data_o_260_sv2v_reg;
  assign data_o[259] = data_o_259_sv2v_reg;
  assign data_o[258] = data_o_258_sv2v_reg;
  assign data_o[257] = data_o_257_sv2v_reg;
  assign data_o[256] = data_o_256_sv2v_reg;
  assign data_o[255] = data_o_255_sv2v_reg;
  assign data_o[254] = data_o_254_sv2v_reg;
  assign data_o[253] = data_o_253_sv2v_reg;
  assign data_o[252] = data_o_252_sv2v_reg;
  assign data_o[251] = data_o_251_sv2v_reg;
  assign data_o[250] = data_o_250_sv2v_reg;
  assign data_o[249] = data_o_249_sv2v_reg;
  assign data_o[248] = data_o_248_sv2v_reg;
  assign data_o[247] = data_o_247_sv2v_reg;
  assign data_o[246] = data_o_246_sv2v_reg;
  assign data_o[245] = data_o_245_sv2v_reg;
  assign data_o[244] = data_o_244_sv2v_reg;
  assign data_o[243] = data_o_243_sv2v_reg;
  assign data_o[242] = data_o_242_sv2v_reg;
  assign data_o[241] = data_o_241_sv2v_reg;
  assign data_o[240] = data_o_240_sv2v_reg;
  assign data_o[239] = data_o_239_sv2v_reg;
  assign data_o[238] = data_o_238_sv2v_reg;
  assign data_o[237] = data_o_237_sv2v_reg;
  assign data_o[236] = data_o_236_sv2v_reg;
  assign data_o[235] = data_o_235_sv2v_reg;
  assign data_o[234] = data_o_234_sv2v_reg;
  assign data_o[233] = data_o_233_sv2v_reg;
  assign data_o[232] = data_o_232_sv2v_reg;
  assign data_o[231] = data_o_231_sv2v_reg;
  assign data_o[230] = data_o_230_sv2v_reg;
  assign data_o[229] = data_o_229_sv2v_reg;
  assign data_o[228] = data_o_228_sv2v_reg;
  assign data_o[227] = data_o_227_sv2v_reg;
  assign data_o[226] = data_o_226_sv2v_reg;
  assign data_o[225] = data_o_225_sv2v_reg;
  assign data_o[224] = data_o_224_sv2v_reg;
  assign data_o[223] = data_o_223_sv2v_reg;
  assign data_o[222] = data_o_222_sv2v_reg;
  assign data_o[221] = data_o_221_sv2v_reg;
  assign data_o[220] = data_o_220_sv2v_reg;
  assign data_o[219] = data_o_219_sv2v_reg;
  assign data_o[218] = data_o_218_sv2v_reg;
  assign data_o[217] = data_o_217_sv2v_reg;
  assign data_o[216] = data_o_216_sv2v_reg;
  assign data_o[215] = data_o_215_sv2v_reg;
  assign data_o[214] = data_o_214_sv2v_reg;
  assign data_o[213] = data_o_213_sv2v_reg;
  assign data_o[212] = data_o_212_sv2v_reg;
  assign data_o[211] = data_o_211_sv2v_reg;
  assign data_o[210] = data_o_210_sv2v_reg;
  assign data_o[209] = data_o_209_sv2v_reg;
  assign data_o[208] = data_o_208_sv2v_reg;
  assign data_o[207] = data_o_207_sv2v_reg;
  assign data_o[206] = data_o_206_sv2v_reg;
  assign data_o[205] = data_o_205_sv2v_reg;
  assign data_o[204] = data_o_204_sv2v_reg;
  assign data_o[203] = data_o_203_sv2v_reg;
  assign data_o[202] = data_o_202_sv2v_reg;
  assign data_o[201] = data_o_201_sv2v_reg;
  assign data_o[200] = data_o_200_sv2v_reg;
  assign data_o[199] = data_o_199_sv2v_reg;
  assign data_o[198] = data_o_198_sv2v_reg;
  assign data_o[197] = data_o_197_sv2v_reg;
  assign data_o[196] = data_o_196_sv2v_reg;
  assign data_o[195] = data_o_195_sv2v_reg;
  assign data_o[194] = data_o_194_sv2v_reg;
  assign data_o[193] = data_o_193_sv2v_reg;
  assign data_o[192] = data_o_192_sv2v_reg;
  assign data_o[191] = data_o_191_sv2v_reg;
  assign data_o[190] = data_o_190_sv2v_reg;
  assign data_o[189] = data_o_189_sv2v_reg;
  assign data_o[188] = data_o_188_sv2v_reg;
  assign data_o[187] = data_o_187_sv2v_reg;
  assign data_o[186] = data_o_186_sv2v_reg;
  assign data_o[185] = data_o_185_sv2v_reg;
  assign data_o[184] = data_o_184_sv2v_reg;
  assign data_o[183] = data_o_183_sv2v_reg;
  assign data_o[182] = data_o_182_sv2v_reg;
  assign data_o[181] = data_o_181_sv2v_reg;
  assign data_o[180] = data_o_180_sv2v_reg;
  assign data_o[179] = data_o_179_sv2v_reg;
  assign data_o[178] = data_o_178_sv2v_reg;
  assign data_o[177] = data_o_177_sv2v_reg;
  assign data_o[176] = data_o_176_sv2v_reg;
  assign data_o[175] = data_o_175_sv2v_reg;
  assign data_o[174] = data_o_174_sv2v_reg;
  assign data_o[173] = data_o_173_sv2v_reg;
  assign data_o[172] = data_o_172_sv2v_reg;
  assign data_o[171] = data_o_171_sv2v_reg;
  assign data_o[170] = data_o_170_sv2v_reg;
  assign data_o[169] = data_o_169_sv2v_reg;
  assign data_o[168] = data_o_168_sv2v_reg;
  assign data_o[167] = data_o_167_sv2v_reg;
  assign data_o[166] = data_o_166_sv2v_reg;
  assign data_o[165] = data_o_165_sv2v_reg;
  assign data_o[164] = data_o_164_sv2v_reg;
  assign data_o[163] = data_o_163_sv2v_reg;
  assign data_o[162] = data_o_162_sv2v_reg;
  assign data_o[161] = data_o_161_sv2v_reg;
  assign data_o[160] = data_o_160_sv2v_reg;
  assign data_o[159] = data_o_159_sv2v_reg;
  assign data_o[158] = data_o_158_sv2v_reg;
  assign data_o[157] = data_o_157_sv2v_reg;
  assign data_o[156] = data_o_156_sv2v_reg;
  assign data_o[155] = data_o_155_sv2v_reg;
  assign data_o[154] = data_o_154_sv2v_reg;
  assign data_o[153] = data_o_153_sv2v_reg;
  assign data_o[152] = data_o_152_sv2v_reg;
  assign data_o[151] = data_o_151_sv2v_reg;
  assign data_o[150] = data_o_150_sv2v_reg;
  assign data_o[149] = data_o_149_sv2v_reg;
  assign data_o[148] = data_o_148_sv2v_reg;
  assign data_o[147] = data_o_147_sv2v_reg;
  assign data_o[146] = data_o_146_sv2v_reg;
  assign data_o[145] = data_o_145_sv2v_reg;
  assign data_o[144] = data_o_144_sv2v_reg;
  assign data_o[143] = data_o_143_sv2v_reg;
  assign data_o[142] = data_o_142_sv2v_reg;
  assign data_o[141] = data_o_141_sv2v_reg;
  assign data_o[140] = data_o_140_sv2v_reg;
  assign data_o[139] = data_o_139_sv2v_reg;
  assign data_o[138] = data_o_138_sv2v_reg;
  assign data_o[137] = data_o_137_sv2v_reg;
  assign data_o[136] = data_o_136_sv2v_reg;
  assign data_o[135] = data_o_135_sv2v_reg;
  assign data_o[134] = data_o_134_sv2v_reg;
  assign data_o[133] = data_o_133_sv2v_reg;
  assign data_o[132] = data_o_132_sv2v_reg;
  assign data_o[131] = data_o_131_sv2v_reg;
  assign data_o[130] = data_o_130_sv2v_reg;
  assign data_o[129] = data_o_129_sv2v_reg;
  assign data_o[128] = data_o_128_sv2v_reg;
  assign data_o[127] = data_o_127_sv2v_reg;
  assign data_o[126] = data_o_126_sv2v_reg;
  assign data_o[125] = data_o_125_sv2v_reg;
  assign data_o[124] = data_o_124_sv2v_reg;
  assign data_o[123] = data_o_123_sv2v_reg;
  assign data_o[122] = data_o_122_sv2v_reg;
  assign data_o[121] = data_o_121_sv2v_reg;
  assign data_o[120] = data_o_120_sv2v_reg;
  assign data_o[119] = data_o_119_sv2v_reg;
  assign data_o[118] = data_o_118_sv2v_reg;
  assign data_o[117] = data_o_117_sv2v_reg;
  assign data_o[116] = data_o_116_sv2v_reg;
  assign data_o[115] = data_o_115_sv2v_reg;
  assign data_o[114] = data_o_114_sv2v_reg;
  assign data_o[113] = data_o_113_sv2v_reg;
  assign data_o[112] = data_o_112_sv2v_reg;
  assign data_o[111] = data_o_111_sv2v_reg;
  assign data_o[110] = data_o_110_sv2v_reg;
  assign data_o[109] = data_o_109_sv2v_reg;
  assign data_o[108] = data_o_108_sv2v_reg;
  assign data_o[107] = data_o_107_sv2v_reg;
  assign data_o[106] = data_o_106_sv2v_reg;
  assign data_o[105] = data_o_105_sv2v_reg;
  assign data_o[104] = data_o_104_sv2v_reg;
  assign data_o[103] = data_o_103_sv2v_reg;
  assign data_o[102] = data_o_102_sv2v_reg;
  assign data_o[101] = data_o_101_sv2v_reg;
  assign data_o[100] = data_o_100_sv2v_reg;
  assign data_o[99] = data_o_99_sv2v_reg;
  assign data_o[98] = data_o_98_sv2v_reg;
  assign data_o[97] = data_o_97_sv2v_reg;
  assign data_o[96] = data_o_96_sv2v_reg;
  assign data_o[95] = data_o_95_sv2v_reg;
  assign data_o[94] = data_o_94_sv2v_reg;
  assign data_o[93] = data_o_93_sv2v_reg;
  assign data_o[92] = data_o_92_sv2v_reg;
  assign data_o[91] = data_o_91_sv2v_reg;
  assign data_o[90] = data_o_90_sv2v_reg;
  assign data_o[89] = data_o_89_sv2v_reg;
  assign data_o[88] = data_o_88_sv2v_reg;
  assign data_o[87] = data_o_87_sv2v_reg;
  assign data_o[86] = data_o_86_sv2v_reg;
  assign data_o[85] = data_o_85_sv2v_reg;
  assign data_o[84] = data_o_84_sv2v_reg;
  assign data_o[83] = data_o_83_sv2v_reg;
  assign data_o[82] = data_o_82_sv2v_reg;
  assign data_o[81] = data_o_81_sv2v_reg;
  assign data_o[80] = data_o_80_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_365_sv2v_reg <= data_i[365];
      data_o_364_sv2v_reg <= data_i[364];
      data_o_363_sv2v_reg <= data_i[363];
      data_o_362_sv2v_reg <= data_i[362];
      data_o_361_sv2v_reg <= data_i[361];
      data_o_360_sv2v_reg <= data_i[360];
      data_o_359_sv2v_reg <= data_i[359];
      data_o_358_sv2v_reg <= data_i[358];
      data_o_357_sv2v_reg <= data_i[357];
      data_o_356_sv2v_reg <= data_i[356];
      data_o_355_sv2v_reg <= data_i[355];
      data_o_354_sv2v_reg <= data_i[354];
      data_o_353_sv2v_reg <= data_i[353];
      data_o_352_sv2v_reg <= data_i[352];
      data_o_351_sv2v_reg <= data_i[351];
      data_o_350_sv2v_reg <= data_i[350];
      data_o_349_sv2v_reg <= data_i[349];
      data_o_348_sv2v_reg <= data_i[348];
      data_o_347_sv2v_reg <= data_i[347];
      data_o_346_sv2v_reg <= data_i[346];
      data_o_345_sv2v_reg <= data_i[345];
      data_o_344_sv2v_reg <= data_i[344];
      data_o_343_sv2v_reg <= data_i[343];
      data_o_342_sv2v_reg <= data_i[342];
      data_o_341_sv2v_reg <= data_i[341];
      data_o_340_sv2v_reg <= data_i[340];
      data_o_339_sv2v_reg <= data_i[339];
      data_o_338_sv2v_reg <= data_i[338];
      data_o_337_sv2v_reg <= data_i[337];
      data_o_336_sv2v_reg <= data_i[336];
      data_o_335_sv2v_reg <= data_i[335];
      data_o_334_sv2v_reg <= data_i[334];
      data_o_333_sv2v_reg <= data_i[333];
      data_o_332_sv2v_reg <= data_i[332];
      data_o_331_sv2v_reg <= data_i[331];
      data_o_330_sv2v_reg <= data_i[330];
      data_o_329_sv2v_reg <= data_i[329];
      data_o_328_sv2v_reg <= data_i[328];
      data_o_327_sv2v_reg <= data_i[327];
      data_o_326_sv2v_reg <= data_i[326];
      data_o_325_sv2v_reg <= data_i[325];
      data_o_324_sv2v_reg <= data_i[324];
      data_o_323_sv2v_reg <= data_i[323];
      data_o_322_sv2v_reg <= data_i[322];
      data_o_321_sv2v_reg <= data_i[321];
      data_o_320_sv2v_reg <= data_i[320];
      data_o_319_sv2v_reg <= data_i[319];
      data_o_318_sv2v_reg <= data_i[318];
      data_o_317_sv2v_reg <= data_i[317];
      data_o_316_sv2v_reg <= data_i[316];
      data_o_315_sv2v_reg <= data_i[315];
      data_o_314_sv2v_reg <= data_i[314];
      data_o_313_sv2v_reg <= data_i[313];
      data_o_312_sv2v_reg <= data_i[312];
      data_o_311_sv2v_reg <= data_i[311];
      data_o_310_sv2v_reg <= data_i[310];
      data_o_309_sv2v_reg <= data_i[309];
      data_o_308_sv2v_reg <= data_i[308];
      data_o_307_sv2v_reg <= data_i[307];
      data_o_306_sv2v_reg <= data_i[306];
      data_o_305_sv2v_reg <= data_i[305];
      data_o_304_sv2v_reg <= data_i[304];
      data_o_303_sv2v_reg <= data_i[303];
      data_o_302_sv2v_reg <= data_i[302];
      data_o_301_sv2v_reg <= data_i[301];
      data_o_300_sv2v_reg <= data_i[300];
      data_o_299_sv2v_reg <= data_i[299];
      data_o_298_sv2v_reg <= data_i[298];
      data_o_297_sv2v_reg <= data_i[297];
      data_o_296_sv2v_reg <= data_i[296];
      data_o_295_sv2v_reg <= data_i[295];
      data_o_294_sv2v_reg <= data_i[294];
      data_o_293_sv2v_reg <= data_i[293];
      data_o_292_sv2v_reg <= data_i[292];
      data_o_291_sv2v_reg <= data_i[291];
      data_o_290_sv2v_reg <= data_i[290];
      data_o_289_sv2v_reg <= data_i[289];
      data_o_288_sv2v_reg <= data_i[288];
      data_o_287_sv2v_reg <= data_i[287];
      data_o_286_sv2v_reg <= data_i[286];
      data_o_285_sv2v_reg <= data_i[285];
      data_o_284_sv2v_reg <= data_i[284];
      data_o_283_sv2v_reg <= data_i[283];
      data_o_282_sv2v_reg <= data_i[282];
      data_o_281_sv2v_reg <= data_i[281];
      data_o_280_sv2v_reg <= data_i[280];
      data_o_279_sv2v_reg <= data_i[279];
      data_o_278_sv2v_reg <= data_i[278];
      data_o_277_sv2v_reg <= data_i[277];
      data_o_276_sv2v_reg <= data_i[276];
      data_o_275_sv2v_reg <= data_i[275];
      data_o_274_sv2v_reg <= data_i[274];
      data_o_273_sv2v_reg <= data_i[273];
      data_o_272_sv2v_reg <= data_i[272];
      data_o_271_sv2v_reg <= data_i[271];
      data_o_270_sv2v_reg <= data_i[270];
      data_o_269_sv2v_reg <= data_i[269];
      data_o_268_sv2v_reg <= data_i[268];
      data_o_267_sv2v_reg <= data_i[267];
      data_o_266_sv2v_reg <= data_i[266];
      data_o_265_sv2v_reg <= data_i[265];
      data_o_264_sv2v_reg <= data_i[264];
      data_o_263_sv2v_reg <= data_i[263];
      data_o_262_sv2v_reg <= data_i[262];
      data_o_261_sv2v_reg <= data_i[261];
      data_o_260_sv2v_reg <= data_i[260];
      data_o_259_sv2v_reg <= data_i[259];
      data_o_258_sv2v_reg <= data_i[258];
      data_o_257_sv2v_reg <= data_i[257];
      data_o_256_sv2v_reg <= data_i[256];
      data_o_255_sv2v_reg <= data_i[255];
      data_o_254_sv2v_reg <= data_i[254];
      data_o_253_sv2v_reg <= data_i[253];
      data_o_252_sv2v_reg <= data_i[252];
      data_o_251_sv2v_reg <= data_i[251];
      data_o_250_sv2v_reg <= data_i[250];
      data_o_249_sv2v_reg <= data_i[249];
      data_o_248_sv2v_reg <= data_i[248];
      data_o_247_sv2v_reg <= data_i[247];
      data_o_246_sv2v_reg <= data_i[246];
      data_o_245_sv2v_reg <= data_i[245];
      data_o_244_sv2v_reg <= data_i[244];
      data_o_243_sv2v_reg <= data_i[243];
      data_o_242_sv2v_reg <= data_i[242];
      data_o_241_sv2v_reg <= data_i[241];
      data_o_240_sv2v_reg <= data_i[240];
      data_o_239_sv2v_reg <= data_i[239];
      data_o_238_sv2v_reg <= data_i[238];
      data_o_237_sv2v_reg <= data_i[237];
      data_o_236_sv2v_reg <= data_i[236];
      data_o_235_sv2v_reg <= data_i[235];
      data_o_234_sv2v_reg <= data_i[234];
      data_o_233_sv2v_reg <= data_i[233];
      data_o_232_sv2v_reg <= data_i[232];
      data_o_231_sv2v_reg <= data_i[231];
      data_o_230_sv2v_reg <= data_i[230];
      data_o_229_sv2v_reg <= data_i[229];
      data_o_228_sv2v_reg <= data_i[228];
      data_o_227_sv2v_reg <= data_i[227];
      data_o_226_sv2v_reg <= data_i[226];
      data_o_225_sv2v_reg <= data_i[225];
      data_o_224_sv2v_reg <= data_i[224];
      data_o_223_sv2v_reg <= data_i[223];
      data_o_222_sv2v_reg <= data_i[222];
      data_o_221_sv2v_reg <= data_i[221];
      data_o_220_sv2v_reg <= data_i[220];
      data_o_219_sv2v_reg <= data_i[219];
      data_o_218_sv2v_reg <= data_i[218];
      data_o_217_sv2v_reg <= data_i[217];
      data_o_216_sv2v_reg <= data_i[216];
      data_o_215_sv2v_reg <= data_i[215];
      data_o_214_sv2v_reg <= data_i[214];
      data_o_213_sv2v_reg <= data_i[213];
      data_o_212_sv2v_reg <= data_i[212];
      data_o_211_sv2v_reg <= data_i[211];
      data_o_210_sv2v_reg <= data_i[210];
      data_o_209_sv2v_reg <= data_i[209];
      data_o_208_sv2v_reg <= data_i[208];
      data_o_207_sv2v_reg <= data_i[207];
      data_o_206_sv2v_reg <= data_i[206];
      data_o_205_sv2v_reg <= data_i[205];
      data_o_204_sv2v_reg <= data_i[204];
      data_o_203_sv2v_reg <= data_i[203];
      data_o_202_sv2v_reg <= data_i[202];
      data_o_201_sv2v_reg <= data_i[201];
      data_o_200_sv2v_reg <= data_i[200];
      data_o_199_sv2v_reg <= data_i[199];
      data_o_198_sv2v_reg <= data_i[198];
      data_o_197_sv2v_reg <= data_i[197];
      data_o_196_sv2v_reg <= data_i[196];
      data_o_195_sv2v_reg <= data_i[195];
      data_o_194_sv2v_reg <= data_i[194];
      data_o_193_sv2v_reg <= data_i[193];
      data_o_192_sv2v_reg <= data_i[192];
      data_o_191_sv2v_reg <= data_i[191];
      data_o_190_sv2v_reg <= data_i[190];
      data_o_189_sv2v_reg <= data_i[189];
      data_o_188_sv2v_reg <= data_i[188];
      data_o_187_sv2v_reg <= data_i[187];
      data_o_186_sv2v_reg <= data_i[186];
      data_o_185_sv2v_reg <= data_i[185];
      data_o_184_sv2v_reg <= data_i[184];
      data_o_183_sv2v_reg <= data_i[183];
      data_o_182_sv2v_reg <= data_i[182];
      data_o_181_sv2v_reg <= data_i[181];
      data_o_180_sv2v_reg <= data_i[180];
      data_o_179_sv2v_reg <= data_i[179];
      data_o_178_sv2v_reg <= data_i[178];
      data_o_177_sv2v_reg <= data_i[177];
      data_o_176_sv2v_reg <= data_i[176];
      data_o_175_sv2v_reg <= data_i[175];
      data_o_174_sv2v_reg <= data_i[174];
      data_o_173_sv2v_reg <= data_i[173];
      data_o_172_sv2v_reg <= data_i[172];
      data_o_171_sv2v_reg <= data_i[171];
      data_o_170_sv2v_reg <= data_i[170];
      data_o_169_sv2v_reg <= data_i[169];
      data_o_168_sv2v_reg <= data_i[168];
      data_o_167_sv2v_reg <= data_i[167];
      data_o_166_sv2v_reg <= data_i[166];
      data_o_165_sv2v_reg <= data_i[165];
      data_o_164_sv2v_reg <= data_i[164];
      data_o_163_sv2v_reg <= data_i[163];
      data_o_162_sv2v_reg <= data_i[162];
      data_o_161_sv2v_reg <= data_i[161];
      data_o_160_sv2v_reg <= data_i[160];
      data_o_159_sv2v_reg <= data_i[159];
      data_o_158_sv2v_reg <= data_i[158];
      data_o_157_sv2v_reg <= data_i[157];
      data_o_156_sv2v_reg <= data_i[156];
      data_o_155_sv2v_reg <= data_i[155];
      data_o_154_sv2v_reg <= data_i[154];
      data_o_153_sv2v_reg <= data_i[153];
      data_o_152_sv2v_reg <= data_i[152];
      data_o_151_sv2v_reg <= data_i[151];
      data_o_150_sv2v_reg <= data_i[150];
      data_o_149_sv2v_reg <= data_i[149];
      data_o_148_sv2v_reg <= data_i[148];
      data_o_147_sv2v_reg <= data_i[147];
      data_o_146_sv2v_reg <= data_i[146];
      data_o_145_sv2v_reg <= data_i[145];
      data_o_144_sv2v_reg <= data_i[144];
      data_o_143_sv2v_reg <= data_i[143];
      data_o_142_sv2v_reg <= data_i[142];
      data_o_141_sv2v_reg <= data_i[141];
      data_o_140_sv2v_reg <= data_i[140];
      data_o_139_sv2v_reg <= data_i[139];
      data_o_138_sv2v_reg <= data_i[138];
      data_o_137_sv2v_reg <= data_i[137];
      data_o_136_sv2v_reg <= data_i[136];
      data_o_135_sv2v_reg <= data_i[135];
      data_o_134_sv2v_reg <= data_i[134];
      data_o_133_sv2v_reg <= data_i[133];
      data_o_132_sv2v_reg <= data_i[132];
      data_o_131_sv2v_reg <= data_i[131];
      data_o_130_sv2v_reg <= data_i[130];
      data_o_129_sv2v_reg <= data_i[129];
      data_o_128_sv2v_reg <= data_i[128];
      data_o_127_sv2v_reg <= data_i[127];
      data_o_126_sv2v_reg <= data_i[126];
      data_o_125_sv2v_reg <= data_i[125];
      data_o_124_sv2v_reg <= data_i[124];
      data_o_123_sv2v_reg <= data_i[123];
      data_o_122_sv2v_reg <= data_i[122];
      data_o_121_sv2v_reg <= data_i[121];
      data_o_120_sv2v_reg <= data_i[120];
      data_o_119_sv2v_reg <= data_i[119];
      data_o_118_sv2v_reg <= data_i[118];
      data_o_117_sv2v_reg <= data_i[117];
      data_o_116_sv2v_reg <= data_i[116];
      data_o_115_sv2v_reg <= data_i[115];
      data_o_114_sv2v_reg <= data_i[114];
      data_o_113_sv2v_reg <= data_i[113];
      data_o_112_sv2v_reg <= data_i[112];
      data_o_111_sv2v_reg <= data_i[111];
      data_o_110_sv2v_reg <= data_i[110];
      data_o_109_sv2v_reg <= data_i[109];
      data_o_108_sv2v_reg <= data_i[108];
      data_o_107_sv2v_reg <= data_i[107];
      data_o_106_sv2v_reg <= data_i[106];
      data_o_105_sv2v_reg <= data_i[105];
      data_o_104_sv2v_reg <= data_i[104];
      data_o_103_sv2v_reg <= data_i[103];
      data_o_102_sv2v_reg <= data_i[102];
      data_o_101_sv2v_reg <= data_i[101];
      data_o_100_sv2v_reg <= data_i[100];
      data_o_99_sv2v_reg <= data_i[99];
      data_o_98_sv2v_reg <= data_i[98];
      data_o_97_sv2v_reg <= data_i[97];
      data_o_96_sv2v_reg <= data_i[96];
      data_o_95_sv2v_reg <= data_i[95];
      data_o_94_sv2v_reg <= data_i[94];
      data_o_93_sv2v_reg <= data_i[93];
      data_o_92_sv2v_reg <= data_i[92];
      data_o_91_sv2v_reg <= data_i[91];
      data_o_90_sv2v_reg <= data_i[90];
      data_o_89_sv2v_reg <= data_i[89];
      data_o_88_sv2v_reg <= data_i[88];
      data_o_87_sv2v_reg <= data_i[87];
      data_o_86_sv2v_reg <= data_i[86];
      data_o_85_sv2v_reg <= data_i[85];
      data_o_84_sv2v_reg <= data_i[84];
      data_o_83_sv2v_reg <= data_i[83];
      data_o_82_sv2v_reg <= data_i[82];
      data_o_81_sv2v_reg <= data_i[81];
      data_o_80_sv2v_reg <= data_i[80];
      data_o_79_sv2v_reg <= data_i[79];
      data_o_78_sv2v_reg <= data_i[78];
      data_o_77_sv2v_reg <= data_i[77];
      data_o_76_sv2v_reg <= data_i[76];
      data_o_75_sv2v_reg <= data_i[75];
      data_o_74_sv2v_reg <= data_i[74];
      data_o_73_sv2v_reg <= data_i[73];
      data_o_72_sv2v_reg <= data_i[72];
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module recFNToRawFN_expWidth8_sigWidth24
(
  in,
  isNaN,
  isInf,
  isZero,
  sign,
  sExp,
  sig
);

  input [32:0] in;
  output [9:0] sExp;
  output [24:0] sig;
  output isNaN;
  output isInf;
  output isZero;
  output sign;
  wire [9:0] sExp;
  wire [24:0] sig;
  wire isNaN,isInf,isZero,sign,in_32_,sExp_8_,sExp_7_,sExp_6_,sExp_5_,sExp_4_,sExp_3_,
  sExp_2_,sExp_1_,sExp_0_,sig_22_,sig_21_,sig_20_,sig_19_,sig_18_,sig_17_,sig_16_,
  sig_15_,sig_14_,sig_13_,sig_12_,sig_11_,sig_10_,sig_9_,sig_8_,sig_7_,sig_6_,
  sig_5_,sig_4_,sig_3_,sig_2_,sig_1_,sig_0_,N0,N1,N2,N4;
  assign sig[24] = 1'b0;
  assign sExp[9] = 1'b0;
  assign in_32_ = in[32];
  assign sign = in_32_;
  assign sExp_8_ = in[31];
  assign sExp[8] = sExp_8_;
  assign sExp_7_ = in[30];
  assign sExp[7] = sExp_7_;
  assign sExp_6_ = in[29];
  assign sExp[6] = sExp_6_;
  assign sExp_5_ = in[28];
  assign sExp[5] = sExp_5_;
  assign sExp_4_ = in[27];
  assign sExp[4] = sExp_4_;
  assign sExp_3_ = in[26];
  assign sExp[3] = sExp_3_;
  assign sExp_2_ = in[25];
  assign sExp[2] = sExp_2_;
  assign sExp_1_ = in[24];
  assign sExp[1] = sExp_1_;
  assign sExp_0_ = in[23];
  assign sExp[0] = sExp_0_;
  assign sig_22_ = in[22];
  assign sig[22] = sig_22_;
  assign sig_21_ = in[21];
  assign sig[21] = sig_21_;
  assign sig_20_ = in[20];
  assign sig[20] = sig_20_;
  assign sig_19_ = in[19];
  assign sig[19] = sig_19_;
  assign sig_18_ = in[18];
  assign sig[18] = sig_18_;
  assign sig_17_ = in[17];
  assign sig[17] = sig_17_;
  assign sig_16_ = in[16];
  assign sig[16] = sig_16_;
  assign sig_15_ = in[15];
  assign sig[15] = sig_15_;
  assign sig_14_ = in[14];
  assign sig[14] = sig_14_;
  assign sig_13_ = in[13];
  assign sig[13] = sig_13_;
  assign sig_12_ = in[12];
  assign sig[12] = sig_12_;
  assign sig_11_ = in[11];
  assign sig[11] = sig_11_;
  assign sig_10_ = in[10];
  assign sig[10] = sig_10_;
  assign sig_9_ = in[9];
  assign sig[9] = sig_9_;
  assign sig_8_ = in[8];
  assign sig[8] = sig_8_;
  assign sig_7_ = in[7];
  assign sig[7] = sig_7_;
  assign sig_6_ = in[6];
  assign sig[6] = sig_6_;
  assign sig_5_ = in[5];
  assign sig[5] = sig_5_;
  assign sig_4_ = in[4];
  assign sig[4] = sig_4_;
  assign sig_3_ = in[3];
  assign sig[3] = sig_3_;
  assign sig_2_ = in[2];
  assign sig[2] = sig_2_;
  assign sig_1_ = in[1];
  assign sig[1] = sig_1_;
  assign sig_0_ = in[0];
  assign sig[0] = sig_0_;
  assign N0 = sExp_7_ & sExp_8_;
  assign N1 = sExp_7_ | sExp_8_;
  assign N2 = sExp_6_ | N1;
  assign isZero = ~N2;
  assign isNaN = N0 & sExp_6_;
  assign isInf = N0 & N4;
  assign N4 = ~sExp_6_;
  assign sig[23] = ~isZero;

endmodule



module recFNToFN_expWidth8_sigWidth24
(
  in,
  out
);

  input [32:0] in;
  output [31:0] out;
  wire [31:0] out;
  wire N0,N1,isNaN,isInf,isZero,N2,isSubnormal,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,
  N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,
  N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,sv2v_dc_1;
  wire [9:0] sExp;
  wire [24:0] sig;
  wire [4:0] denormShiftDist;

  recFNToRawFN_expWidth8_sigWidth24
  recFNToRawFN
  (
    .in(in),
    .isNaN(isNaN),
    .isInf(isInf),
    .isZero(isZero),
    .sign(out[31]),
    .sExp(sExp),
    .sig(sig)
  );

  assign N2 = sExp[5:0] <= 1'b1;
  assign N56 = ~sExp[7];
  assign N57 = sExp[8] | sExp[9];
  assign N58 = N56 | N57;
  assign N59 = sExp[6] | N58;
  assign N60 = ~N59;
  assign N61 = sExp[8] | sExp[9];
  assign N62 = sExp[7] | N61;
  assign N63 = ~N62;
  assign denormShiftDist = 1'b1 - sExp[4:0];
  assign { sv2v_dc_1, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31 } = sig[24:1] >> denormShiftDist;
  assign { N11, N10, N9, N8, N7, N6, N5, N4 } = sExp[7:0] - { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 };
  assign { N19, N18, N17, N16, N15, N14, N13, N12 } = { N11, N10, N9, N8, N7, N6, N5, N4 } + 1'b1;
  assign { N27, N26, N25, N24, N23, N22, N21, N20 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                      (N1)? { N19, N18, N17, N16, N15, N14, N13, N12 } : 1'b0;
  assign N0 = isSubnormal;
  assign N1 = N3;
  assign out[22:0] = (N0)? { N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31 } : 
                     (N55)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                     (N30)? sig[22:0] : 1'b0;
  assign isSubnormal = N64 | N63;
  assign N64 = N60 & N2;
  assign N3 = ~isSubnormal;
  assign N28 = isNaN | isInf;
  assign out[30] = N27 | N28;
  assign out[29] = N26 | N28;
  assign out[28] = N25 | N28;
  assign out[27] = N24 | N28;
  assign out[26] = N23 | N28;
  assign out[25] = N22 | N28;
  assign out[24] = N21 | N28;
  assign out[23] = N20 | N28;
  assign N29 = isInf | isSubnormal;
  assign N30 = ~N29;
  assign N54 = ~isSubnormal;
  assign N55 = isInf & N54;

endmodule



module recFNToRawFN_expWidth11_sigWidth53
(
  in,
  isNaN,
  isInf,
  isZero,
  sign,
  sExp,
  sig
);

  input [64:0] in;
  output [12:0] sExp;
  output [53:0] sig;
  output isNaN;
  output isInf;
  output isZero;
  output sign;
  wire [12:0] sExp;
  wire [53:0] sig;
  wire isNaN,isInf,isZero,sign,in_64_,sExp_11_,sExp_10_,sExp_9_,sExp_8_,sExp_7_,
  sExp_6_,sExp_5_,sExp_4_,sExp_3_,sExp_2_,sExp_1_,sExp_0_,sig_51_,sig_50_,sig_49_,
  sig_48_,sig_47_,sig_46_,sig_45_,sig_44_,sig_43_,sig_42_,sig_41_,sig_40_,sig_39_,
  sig_38_,sig_37_,sig_36_,sig_35_,sig_34_,sig_33_,sig_32_,sig_31_,sig_30_,sig_29_,
  sig_28_,sig_27_,sig_26_,sig_25_,sig_24_,sig_23_,sig_22_,sig_21_,sig_20_,sig_19_,
  sig_18_,sig_17_,sig_16_,sig_15_,sig_14_,sig_13_,sig_12_,sig_11_,sig_10_,sig_9_,sig_8_,
  sig_7_,sig_6_,sig_5_,sig_4_,sig_3_,sig_2_,sig_1_,sig_0_,N0,N1,N2,N4;
  assign sig[53] = 1'b0;
  assign sExp[12] = 1'b0;
  assign in_64_ = in[64];
  assign sign = in_64_;
  assign sExp_11_ = in[63];
  assign sExp[11] = sExp_11_;
  assign sExp_10_ = in[62];
  assign sExp[10] = sExp_10_;
  assign sExp_9_ = in[61];
  assign sExp[9] = sExp_9_;
  assign sExp_8_ = in[60];
  assign sExp[8] = sExp_8_;
  assign sExp_7_ = in[59];
  assign sExp[7] = sExp_7_;
  assign sExp_6_ = in[58];
  assign sExp[6] = sExp_6_;
  assign sExp_5_ = in[57];
  assign sExp[5] = sExp_5_;
  assign sExp_4_ = in[56];
  assign sExp[4] = sExp_4_;
  assign sExp_3_ = in[55];
  assign sExp[3] = sExp_3_;
  assign sExp_2_ = in[54];
  assign sExp[2] = sExp_2_;
  assign sExp_1_ = in[53];
  assign sExp[1] = sExp_1_;
  assign sExp_0_ = in[52];
  assign sExp[0] = sExp_0_;
  assign sig_51_ = in[51];
  assign sig[51] = sig_51_;
  assign sig_50_ = in[50];
  assign sig[50] = sig_50_;
  assign sig_49_ = in[49];
  assign sig[49] = sig_49_;
  assign sig_48_ = in[48];
  assign sig[48] = sig_48_;
  assign sig_47_ = in[47];
  assign sig[47] = sig_47_;
  assign sig_46_ = in[46];
  assign sig[46] = sig_46_;
  assign sig_45_ = in[45];
  assign sig[45] = sig_45_;
  assign sig_44_ = in[44];
  assign sig[44] = sig_44_;
  assign sig_43_ = in[43];
  assign sig[43] = sig_43_;
  assign sig_42_ = in[42];
  assign sig[42] = sig_42_;
  assign sig_41_ = in[41];
  assign sig[41] = sig_41_;
  assign sig_40_ = in[40];
  assign sig[40] = sig_40_;
  assign sig_39_ = in[39];
  assign sig[39] = sig_39_;
  assign sig_38_ = in[38];
  assign sig[38] = sig_38_;
  assign sig_37_ = in[37];
  assign sig[37] = sig_37_;
  assign sig_36_ = in[36];
  assign sig[36] = sig_36_;
  assign sig_35_ = in[35];
  assign sig[35] = sig_35_;
  assign sig_34_ = in[34];
  assign sig[34] = sig_34_;
  assign sig_33_ = in[33];
  assign sig[33] = sig_33_;
  assign sig_32_ = in[32];
  assign sig[32] = sig_32_;
  assign sig_31_ = in[31];
  assign sig[31] = sig_31_;
  assign sig_30_ = in[30];
  assign sig[30] = sig_30_;
  assign sig_29_ = in[29];
  assign sig[29] = sig_29_;
  assign sig_28_ = in[28];
  assign sig[28] = sig_28_;
  assign sig_27_ = in[27];
  assign sig[27] = sig_27_;
  assign sig_26_ = in[26];
  assign sig[26] = sig_26_;
  assign sig_25_ = in[25];
  assign sig[25] = sig_25_;
  assign sig_24_ = in[24];
  assign sig[24] = sig_24_;
  assign sig_23_ = in[23];
  assign sig[23] = sig_23_;
  assign sig_22_ = in[22];
  assign sig[22] = sig_22_;
  assign sig_21_ = in[21];
  assign sig[21] = sig_21_;
  assign sig_20_ = in[20];
  assign sig[20] = sig_20_;
  assign sig_19_ = in[19];
  assign sig[19] = sig_19_;
  assign sig_18_ = in[18];
  assign sig[18] = sig_18_;
  assign sig_17_ = in[17];
  assign sig[17] = sig_17_;
  assign sig_16_ = in[16];
  assign sig[16] = sig_16_;
  assign sig_15_ = in[15];
  assign sig[15] = sig_15_;
  assign sig_14_ = in[14];
  assign sig[14] = sig_14_;
  assign sig_13_ = in[13];
  assign sig[13] = sig_13_;
  assign sig_12_ = in[12];
  assign sig[12] = sig_12_;
  assign sig_11_ = in[11];
  assign sig[11] = sig_11_;
  assign sig_10_ = in[10];
  assign sig[10] = sig_10_;
  assign sig_9_ = in[9];
  assign sig[9] = sig_9_;
  assign sig_8_ = in[8];
  assign sig[8] = sig_8_;
  assign sig_7_ = in[7];
  assign sig[7] = sig_7_;
  assign sig_6_ = in[6];
  assign sig[6] = sig_6_;
  assign sig_5_ = in[5];
  assign sig[5] = sig_5_;
  assign sig_4_ = in[4];
  assign sig[4] = sig_4_;
  assign sig_3_ = in[3];
  assign sig[3] = sig_3_;
  assign sig_2_ = in[2];
  assign sig[2] = sig_2_;
  assign sig_1_ = in[1];
  assign sig[1] = sig_1_;
  assign sig_0_ = in[0];
  assign sig[0] = sig_0_;
  assign N0 = sExp_10_ & sExp_11_;
  assign N1 = sExp_10_ | sExp_11_;
  assign N2 = sExp_9_ | N1;
  assign isZero = ~N2;
  assign isNaN = N0 & sExp_9_;
  assign isInf = N0 & N4;
  assign N4 = ~sExp_9_;
  assign sig[52] = ~isZero;

endmodule



module recFNToFN_expWidth11_sigWidth53
(
  in,
  out
);

  input [64:0] in;
  output [63:0] out;
  wire [63:0] out;
  wire N0,N1,isNaN,isInf,isZero,N2,isSubnormal,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,
  N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,
  N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,
  N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,
  N94,N95,N96,N97,N98,N99,N100,N101,N102,sv2v_dc_1;
  wire [12:0] sExp;
  wire [53:0] sig;
  wire [5:0] denormShiftDist;

  recFNToRawFN_expWidth11_sigWidth53
  recFNToRawFN
  (
    .in(in),
    .isNaN(isNaN),
    .isInf(isInf),
    .isZero(isZero),
    .sign(out[63]),
    .sExp(sExp),
    .sig(sig)
  );

  assign N2 = sExp[8:0] <= 1'b1;
  assign N94 = ~sExp[10];
  assign N95 = sExp[11] | sExp[12];
  assign N96 = N94 | N95;
  assign N97 = sExp[9] | N96;
  assign N98 = ~N97;
  assign N99 = sExp[11] | sExp[12];
  assign N100 = sExp[10] | N99;
  assign N101 = ~N100;
  assign denormShiftDist = 1'b1 - sExp[5:0];
  assign { sv2v_dc_1, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40 } = sig[53:1] >> denormShiftDist;
  assign { N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4 } = sExp[10:0] - { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 };
  assign { N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15 } = { N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4 } + 1'b1;
  assign { N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                     (N1)? { N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15 } : 1'b0;
  assign N0 = isSubnormal;
  assign N1 = N3;
  assign out[51:0] = (N0)? { N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40 } : 
                     (N93)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                     (N39)? sig[51:0] : 1'b0;
  assign isSubnormal = N102 | N101;
  assign N102 = N98 & N2;
  assign N3 = ~isSubnormal;
  assign N37 = isNaN | isInf;
  assign out[62] = N36 | N37;
  assign out[61] = N35 | N37;
  assign out[60] = N34 | N37;
  assign out[59] = N33 | N37;
  assign out[58] = N32 | N37;
  assign out[57] = N31 | N37;
  assign out[56] = N30 | N37;
  assign out[55] = N29 | N37;
  assign out[54] = N28 | N37;
  assign out[53] = N27 | N37;
  assign out[52] = N26 | N37;
  assign N38 = isInf | isSubnormal;
  assign N39 = ~N38;
  assign N92 = ~isSubnormal;
  assign N93 = isInf & N92;

endmodule



module bp_be_fp_unbox_00
(
  reg_i,
  tag_i,
  raw_i,
  val_o
);

  input [65:0] reg_i;
  input [0:0] tag_i;
  output [64:0] val_o;
  input raw_i;
  wire [64:0] val_o;
  wire N0,N1,N2,N3,N4,N5,special,N6,dp2sp_rec_unsafe_exp__8_,dp2sp_rec_unsafe_exp__7_,
  dp2sp_rec_unsafe_exp__6_,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79;
  wire [8:0] adjusted_exp;
  wire [31:0] dp2sp_raw_lo;
  wire [63:0] dp_raw_lo;
  assign N5 = reg_i[63:61] >= { 1'b1, 1'b1, 1'b0 };

  recFNToFN_expWidth8_sigWidth24
  out_sp_rec
  (
    .in({ reg_i[64:64], dp2sp_rec_unsafe_exp__8_, dp2sp_rec_unsafe_exp__7_, dp2sp_rec_unsafe_exp__6_, adjusted_exp[5:0], reg_i[51:29] }),
    .out(dp2sp_raw_lo)
  );


  recFNToFN_expWidth11_sigWidth53
  out_dp_rec
  (
    .in(reg_i[64:0]),
    .out(dp_raw_lo)
  );

  assign N7 = reg_i[65] ^ tag_i[0];
  assign N76 = ~reg_i[65];
  assign N77 = reg_i[62] | reg_i[63];
  assign N78 = reg_i[61] | N77;
  assign N79 = ~N78;
  assign adjusted_exp = reg_i[60:52] + { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign { dp2sp_rec_unsafe_exp__8_, dp2sp_rec_unsafe_exp__7_, dp2sp_rec_unsafe_exp__6_ } = (N0)? reg_i[63:61] : 
                                                                                            (N1)? adjusted_exp[8:6] : 1'b0;
  assign N0 = special;
  assign N1 = N6;
  assign { N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10 } = (N2)? dp_raw_lo : 
                                                                                                                                                                                                                                                                                                                                              (N3)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, dp2sp_raw_lo } : 1'b0;
  assign N2 = N76;
  assign N3 = reg_i[65];
  assign val_o = (N4)? { 1'b0, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10 } : 
                 (N75)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                 (N9)? reg_i[64:0] : 1'b0;
  assign N4 = raw_i;
  assign special = N79 | N5;
  assign N6 = ~special;
  assign N8 = N7 | raw_i;
  assign N9 = ~N8;
  assign N74 = ~raw_i;
  assign N75 = N7 & N74;

endmodule



module bp_be_int_unbox_00
(
  reg_i,
  tag_i,
  unsigned_i,
  val_o
);

  input [65:0] reg_i;
  input [1:0] tag_i;
  output [64:0] val_o;
  input unsigned_i;
  wire [64:0] val_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,val_o_7_,val_o_6_,
  val_o_5_,val_o_4_,val_o_3_,val_o_2_,val_o_1_,val_o_0_,N16,N17,N18,N19,N20,N21,N22,N23,
  sigbox,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61;
  wire [62:8] raw;
  assign val_o_7_ = reg_i[7];
  assign val_o[7] = val_o_7_;
  assign val_o_6_ = reg_i[6];
  assign val_o[6] = val_o_6_;
  assign val_o_5_ = reg_i[5];
  assign val_o[5] = val_o_5_;
  assign val_o_4_ = reg_i[4];
  assign val_o[4] = val_o_4_;
  assign val_o_3_ = reg_i[3];
  assign val_o[3] = val_o_3_;
  assign val_o_2_ = reg_i[2];
  assign val_o[2] = val_o_2_;
  assign val_o_1_ = reg_i[1];
  assign val_o[1] = val_o_1_;
  assign val_o_0_ = reg_i[0];
  assign val_o[0] = val_o_0_;
  assign N16 = reg_i[65] & reg_i[64];
  assign N17 = N21 | reg_i[64];
  assign N19 = reg_i[65] | N22;
  assign N23 = N21 & N22;
  assign sigbox = tag_i >= reg_i[65:64];
  assign N26 = unsigned_i & N24;
  assign N27 = N26 & N25;
  assign N28 = N26 & tag_i[0];
  assign N29 = unsigned_i & tag_i[1];
  assign N30 = N29 & N25;
  assign N31 = N29 & tag_i[0];
  assign N33 = unsigned_i | N32;
  assign N34 = tag_i[1] | tag_i[0];
  assign N35 = N33 | N34;
  assign N37 = unsigned_i | N32;
  assign N38 = tag_i[1] | N25;
  assign N39 = N37 | N38;
  assign N41 = unsigned_i | N32;
  assign N42 = N24 | tag_i[0];
  assign N43 = N41 | N42;
  assign N45 = unsigned_i | N32;
  assign N46 = N24 | N25;
  assign N47 = N45 | N46;
  assign N50 = N49 & N32;
  assign N51 = N24 & N25;
  assign N52 = N50 & N51;
  assign N53 = unsigned_i | sigbox;
  assign N54 = N53 | N38;
  assign N56 = unsigned_i | sigbox;
  assign N57 = N56 | N42;
  assign N59 = unsigned_i | sigbox;
  assign N60 = N59 | N46;
  assign raw = (N0)? { reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63] } : 
               (N1)? { reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[15:8] } : 
               (N2)? { reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[31:8] } : 
               (N3)? reg_i[62:8] : 1'b0;
  assign N0 = N16;
  assign N1 = N18;
  assign N2 = N20;
  assign N3 = N23;
  assign val_o[64:8] = (N4)? { 1'b0, reg_i[63:63], raw } : 
                       (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, raw[31:8] } : 
                       (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, raw[15:8] } : 
                       (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N8)? { reg_i[63:63], reg_i[63:63], raw } : 
                       (N9)? { raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:31], raw[31:8] } : 
                       (N10)? { raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:15], raw[15:8] } : 
                       (N11)? { val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_, val_o_7_ } : 
                       (N12)? { reg_i[63:63], reg_i[63:63], raw } : 
                       (N13)? { reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], raw[31:8] } : 
                       (N14)? { reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], raw[15:8] } : 
                       (N15)? { reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63], reg_i[63:63] } : 1'b0;
  assign N4 = N27;
  assign N5 = N28;
  assign N6 = N30;
  assign N7 = N31;
  assign N8 = N36;
  assign N9 = N40;
  assign N10 = N44;
  assign N11 = N48;
  assign N12 = N52;
  assign N13 = N55;
  assign N14 = N58;
  assign N15 = N61;
  assign N18 = ~N17;
  assign N20 = ~N19;
  assign N21 = ~reg_i[65];
  assign N22 = ~reg_i[64];
  assign N24 = ~tag_i[1];
  assign N25 = ~tag_i[0];
  assign N32 = ~sigbox;
  assign N36 = ~N35;
  assign N40 = ~N39;
  assign N44 = ~N43;
  assign N48 = ~N47;
  assign N49 = ~unsigned_i;
  assign N55 = ~N54;
  assign N58 = ~N57;
  assign N61 = ~N60;

endmodule



module bp_be_reservation_00
(
  clk_i,
  reset_i,
  dispatch_pkt_i,
  bypass_rs_i,
  reservation_o
);

  input [365:0] dispatch_pkt_i;
  input [197:0] bypass_rs_i;
  output [520:0] reservation_o;
  input clk_i;
  input reset_i;
  wire [520:0] reservation_o;
  wire dispatch_pkt_r_queue_v_,dispatch_pkt_r_ispec_v_,dispatch_pkt_r_nspec_v_,
  dispatch_pkt_r_rs1__65_,dispatch_pkt_r_rs1__64_,dispatch_pkt_r_rs1__63_,
  dispatch_pkt_r_rs1__62_,dispatch_pkt_r_rs1__61_,dispatch_pkt_r_rs1__60_,dispatch_pkt_r_rs1__59_,
  dispatch_pkt_r_rs1__58_,dispatch_pkt_r_rs1__57_,dispatch_pkt_r_rs1__56_,
  dispatch_pkt_r_rs1__55_,dispatch_pkt_r_rs1__54_,dispatch_pkt_r_rs1__53_,
  dispatch_pkt_r_rs1__52_,dispatch_pkt_r_rs1__51_,dispatch_pkt_r_rs1__50_,dispatch_pkt_r_rs1__49_,
  dispatch_pkt_r_rs1__48_,dispatch_pkt_r_rs1__47_,dispatch_pkt_r_rs1__46_,
  dispatch_pkt_r_rs1__45_,dispatch_pkt_r_rs1__44_,dispatch_pkt_r_rs1__43_,
  dispatch_pkt_r_rs1__42_,dispatch_pkt_r_rs1__41_,dispatch_pkt_r_rs1__40_,dispatch_pkt_r_rs1__39_,
  dispatch_pkt_r_rs1__38_,dispatch_pkt_r_rs1__37_,dispatch_pkt_r_rs1__36_,
  dispatch_pkt_r_rs1__35_,dispatch_pkt_r_rs1__34_,dispatch_pkt_r_rs1__33_,
  dispatch_pkt_r_rs1__32_,dispatch_pkt_r_rs1__31_,dispatch_pkt_r_rs1__30_,dispatch_pkt_r_rs1__29_,
  dispatch_pkt_r_rs1__28_,dispatch_pkt_r_rs1__27_,dispatch_pkt_r_rs1__26_,
  dispatch_pkt_r_rs1__25_,dispatch_pkt_r_rs1__24_,dispatch_pkt_r_rs1__23_,
  dispatch_pkt_r_rs1__22_,dispatch_pkt_r_rs1__21_,dispatch_pkt_r_rs1__20_,dispatch_pkt_r_rs1__19_,
  dispatch_pkt_r_rs1__18_,dispatch_pkt_r_rs1__17_,dispatch_pkt_r_rs1__16_,
  dispatch_pkt_r_rs1__15_,dispatch_pkt_r_rs1__14_,dispatch_pkt_r_rs1__13_,
  dispatch_pkt_r_rs1__12_,dispatch_pkt_r_rs1__11_,dispatch_pkt_r_rs1__10_,dispatch_pkt_r_rs1__9_,
  dispatch_pkt_r_rs1__8_,dispatch_pkt_r_rs1__7_,dispatch_pkt_r_rs1__6_,
  dispatch_pkt_r_rs1__5_,dispatch_pkt_r_rs1__4_,dispatch_pkt_r_rs1__3_,dispatch_pkt_r_rs1__2_,
  dispatch_pkt_r_rs1__1_,dispatch_pkt_r_rs1__0_,dispatch_pkt_r_rs2__65_,
  dispatch_pkt_r_rs2__64_,dispatch_pkt_r_rs2__63_,dispatch_pkt_r_rs2__62_,
  dispatch_pkt_r_rs2__61_,dispatch_pkt_r_rs2__60_,dispatch_pkt_r_rs2__59_,dispatch_pkt_r_rs2__58_,
  dispatch_pkt_r_rs2__57_,dispatch_pkt_r_rs2__56_,dispatch_pkt_r_rs2__55_,
  dispatch_pkt_r_rs2__54_,dispatch_pkt_r_rs2__53_,dispatch_pkt_r_rs2__52_,
  dispatch_pkt_r_rs2__51_,dispatch_pkt_r_rs2__50_,dispatch_pkt_r_rs2__49_,dispatch_pkt_r_rs2__48_,
  dispatch_pkt_r_rs2__47_,dispatch_pkt_r_rs2__46_,dispatch_pkt_r_rs2__45_,
  dispatch_pkt_r_rs2__44_,dispatch_pkt_r_rs2__43_,dispatch_pkt_r_rs2__42_,
  dispatch_pkt_r_rs2__41_,dispatch_pkt_r_rs2__40_,dispatch_pkt_r_rs2__39_,dispatch_pkt_r_rs2__38_,
  dispatch_pkt_r_rs2__37_,dispatch_pkt_r_rs2__36_,dispatch_pkt_r_rs2__35_,
  dispatch_pkt_r_rs2__34_,dispatch_pkt_r_rs2__33_,dispatch_pkt_r_rs2__32_,
  dispatch_pkt_r_rs2__31_,dispatch_pkt_r_rs2__30_,dispatch_pkt_r_rs2__29_,dispatch_pkt_r_rs2__28_,
  dispatch_pkt_r_rs2__27_,dispatch_pkt_r_rs2__26_,dispatch_pkt_r_rs2__25_,
  dispatch_pkt_r_rs2__24_,dispatch_pkt_r_rs2__23_,dispatch_pkt_r_rs2__22_,
  dispatch_pkt_r_rs2__21_,dispatch_pkt_r_rs2__20_,dispatch_pkt_r_rs2__19_,dispatch_pkt_r_rs2__18_,
  dispatch_pkt_r_rs2__17_,dispatch_pkt_r_rs2__16_,dispatch_pkt_r_rs2__15_,
  dispatch_pkt_r_rs2__14_,dispatch_pkt_r_rs2__13_,dispatch_pkt_r_rs2__12_,
  dispatch_pkt_r_rs2__11_,dispatch_pkt_r_rs2__10_,dispatch_pkt_r_rs2__9_,dispatch_pkt_r_rs2__8_,
  dispatch_pkt_r_rs2__7_,dispatch_pkt_r_rs2__6_,dispatch_pkt_r_rs2__5_,
  dispatch_pkt_r_rs2__4_,dispatch_pkt_r_rs2__3_,dispatch_pkt_r_rs2__2_,dispatch_pkt_r_rs2__1_,
  dispatch_pkt_r_rs2__0_,dispatch_pkt_r_imm__65_,
  dispatch_pkt_r_exception__store_page_fault_,dispatch_pkt_r_exception__load_page_fault_,
  dispatch_pkt_r_exception__instr_page_fault_,dispatch_pkt_r_exception__ecall_m_,
  dispatch_pkt_r_exception__ecall_s_,dispatch_pkt_r_exception__ecall_u_,
  dispatch_pkt_r_exception__store_access_fault_,dispatch_pkt_r_exception__store_misaligned_,
  dispatch_pkt_r_exception__load_access_fault_,dispatch_pkt_r_exception__load_misaligned_,
  dispatch_pkt_r_exception__ebreak_,dispatch_pkt_r_exception__illegal_instr_,
  dispatch_pkt_r_exception__instr_access_fault_,dispatch_pkt_r_exception__instr_misaligned_,
  dispatch_pkt_r_exception__resume_,dispatch_pkt_r_exception__itlb_miss_,
  dispatch_pkt_r_exception__icache_miss_,dispatch_pkt_r_exception__dcache_replay_,
  dispatch_pkt_r_exception__dtlb_load_miss_,dispatch_pkt_r_exception__dtlb_store_miss_,
  dispatch_pkt_r_exception__itlb_fill_,dispatch_pkt_r_exception__dtlb_fill_,
  dispatch_pkt_r_exception___interrupt_,dispatch_pkt_r_exception__cmd_full_,
  dispatch_pkt_r_exception__mispredict_,dispatch_pkt_r_special__dcache_miss_,dispatch_pkt_r_special__fencei_,
  dispatch_pkt_r_special__sfence_vma_,dispatch_pkt_r_special__dbreak_,
  dispatch_pkt_r_special__dret_,dispatch_pkt_r_special__mret_,dispatch_pkt_r_special__sret_,
  dispatch_pkt_r_special__wfi_,dispatch_pkt_r_special__csrw_;

  bsg_dff_0000016e
  dispatch_pkt_reg
  (
    .clk_i(clk_i),
    .data_i({ dispatch_pkt_i[365:232], bypass_rs_i[65:0], bypass_rs_i[131:66], bypass_rs_i[197:132], dispatch_pkt_i[33:0] }),
    .data_o({ reservation_o[520:520], dispatch_pkt_r_queue_v_, dispatch_pkt_r_ispec_v_, dispatch_pkt_r_nspec_v_, reservation_o[519:449], reservation_o[394:390], reservation_o[448:395], dispatch_pkt_r_rs1__65_, dispatch_pkt_r_rs1__64_, dispatch_pkt_r_rs1__63_, dispatch_pkt_r_rs1__62_, dispatch_pkt_r_rs1__61_, dispatch_pkt_r_rs1__60_, dispatch_pkt_r_rs1__59_, dispatch_pkt_r_rs1__58_, dispatch_pkt_r_rs1__57_, dispatch_pkt_r_rs1__56_, dispatch_pkt_r_rs1__55_, dispatch_pkt_r_rs1__54_, dispatch_pkt_r_rs1__53_, dispatch_pkt_r_rs1__52_, dispatch_pkt_r_rs1__51_, dispatch_pkt_r_rs1__50_, dispatch_pkt_r_rs1__49_, dispatch_pkt_r_rs1__48_, dispatch_pkt_r_rs1__47_, dispatch_pkt_r_rs1__46_, dispatch_pkt_r_rs1__45_, dispatch_pkt_r_rs1__44_, dispatch_pkt_r_rs1__43_, dispatch_pkt_r_rs1__42_, dispatch_pkt_r_rs1__41_, dispatch_pkt_r_rs1__40_, dispatch_pkt_r_rs1__39_, dispatch_pkt_r_rs1__38_, dispatch_pkt_r_rs1__37_, dispatch_pkt_r_rs1__36_, dispatch_pkt_r_rs1__35_, dispatch_pkt_r_rs1__34_, dispatch_pkt_r_rs1__33_, dispatch_pkt_r_rs1__32_, dispatch_pkt_r_rs1__31_, dispatch_pkt_r_rs1__30_, dispatch_pkt_r_rs1__29_, dispatch_pkt_r_rs1__28_, dispatch_pkt_r_rs1__27_, dispatch_pkt_r_rs1__26_, dispatch_pkt_r_rs1__25_, dispatch_pkt_r_rs1__24_, dispatch_pkt_r_rs1__23_, dispatch_pkt_r_rs1__22_, dispatch_pkt_r_rs1__21_, dispatch_pkt_r_rs1__20_, dispatch_pkt_r_rs1__19_, dispatch_pkt_r_rs1__18_, dispatch_pkt_r_rs1__17_, dispatch_pkt_r_rs1__16_, dispatch_pkt_r_rs1__15_, dispatch_pkt_r_rs1__14_, dispatch_pkt_r_rs1__13_, dispatch_pkt_r_rs1__12_, dispatch_pkt_r_rs1__11_, dispatch_pkt_r_rs1__10_, dispatch_pkt_r_rs1__9_, dispatch_pkt_r_rs1__8_, dispatch_pkt_r_rs1__7_, dispatch_pkt_r_rs1__6_, dispatch_pkt_r_rs1__5_, dispatch_pkt_r_rs1__4_, dispatch_pkt_r_rs1__3_, dispatch_pkt_r_rs1__2_, dispatch_pkt_r_rs1__1_, dispatch_pkt_r_rs1__0_, dispatch_pkt_r_rs2__65_, dispatch_pkt_r_rs2__64_, dispatch_pkt_r_rs2__63_, dispatch_pkt_r_rs2__62_, dispatch_pkt_r_rs2__61_, dispatch_pkt_r_rs2__60_, dispatch_pkt_r_rs2__59_, dispatch_pkt_r_rs2__58_, dispatch_pkt_r_rs2__57_, dispatch_pkt_r_rs2__56_, dispatch_pkt_r_rs2__55_, dispatch_pkt_r_rs2__54_, dispatch_pkt_r_rs2__53_, dispatch_pkt_r_rs2__52_, dispatch_pkt_r_rs2__51_, dispatch_pkt_r_rs2__50_, dispatch_pkt_r_rs2__49_, dispatch_pkt_r_rs2__48_, dispatch_pkt_r_rs2__47_, dispatch_pkt_r_rs2__46_, dispatch_pkt_r_rs2__45_, dispatch_pkt_r_rs2__44_, dispatch_pkt_r_rs2__43_, dispatch_pkt_r_rs2__42_, dispatch_pkt_r_rs2__41_, dispatch_pkt_r_rs2__40_, dispatch_pkt_r_rs2__39_, dispatch_pkt_r_rs2__38_, dispatch_pkt_r_rs2__37_, dispatch_pkt_r_rs2__36_, dispatch_pkt_r_rs2__35_, dispatch_pkt_r_rs2__34_, dispatch_pkt_r_rs2__33_, dispatch_pkt_r_rs2__32_, dispatch_pkt_r_rs2__31_, dispatch_pkt_r_rs2__30_, dispatch_pkt_r_rs2__29_, dispatch_pkt_r_rs2__28_, dispatch_pkt_r_rs2__27_, dispatch_pkt_r_rs2__26_, dispatch_pkt_r_rs2__25_, dispatch_pkt_r_rs2__24_, dispatch_pkt_r_rs2__23_, dispatch_pkt_r_rs2__22_, dispatch_pkt_r_rs2__21_, dispatch_pkt_r_rs2__20_, dispatch_pkt_r_rs2__19_, dispatch_pkt_r_rs2__18_, dispatch_pkt_r_rs2__17_, dispatch_pkt_r_rs2__16_, dispatch_pkt_r_rs2__15_, dispatch_pkt_r_rs2__14_, dispatch_pkt_r_rs2__13_, dispatch_pkt_r_rs2__12_, dispatch_pkt_r_rs2__11_, dispatch_pkt_r_rs2__10_, dispatch_pkt_r_rs2__9_, dispatch_pkt_r_rs2__8_, dispatch_pkt_r_rs2__7_, dispatch_pkt_r_rs2__6_, dispatch_pkt_r_rs2__5_, dispatch_pkt_r_rs2__4_, dispatch_pkt_r_rs2__3_, dispatch_pkt_r_rs2__2_, dispatch_pkt_r_rs2__1_, dispatch_pkt_r_rs2__0_, dispatch_pkt_r_imm__65_, reservation_o[259:195], dispatch_pkt_r_exception__store_page_fault_, dispatch_pkt_r_exception__load_page_fault_, dispatch_pkt_r_exception__instr_page_fault_, dispatch_pkt_r_exception__ecall_m_, dispatch_pkt_r_exception__ecall_s_, dispatch_pkt_r_exception__ecall_u_, dispatch_pkt_r_exception__store_access_fault_, dispatch_pkt_r_exception__store_misaligned_, dispatch_pkt_r_exception__load_access_fault_, dispatch_pkt_r_exception__load_misaligned_, dispatch_pkt_r_exception__ebreak_, dispatch_pkt_r_exception__illegal_instr_, dispatch_pkt_r_exception__instr_access_fault_, dispatch_pkt_r_exception__instr_misaligned_, dispatch_pkt_r_exception__resume_, dispatch_pkt_r_exception__itlb_miss_, dispatch_pkt_r_exception__icache_miss_, dispatch_pkt_r_exception__dcache_replay_, dispatch_pkt_r_exception__dtlb_load_miss_, dispatch_pkt_r_exception__dtlb_store_miss_, dispatch_pkt_r_exception__itlb_fill_, dispatch_pkt_r_exception__dtlb_fill_, dispatch_pkt_r_exception___interrupt_, dispatch_pkt_r_exception__cmd_full_, dispatch_pkt_r_exception__mispredict_, dispatch_pkt_r_special__dcache_miss_, dispatch_pkt_r_special__fencei_, dispatch_pkt_r_special__sfence_vma_, dispatch_pkt_r_special__dbreak_, dispatch_pkt_r_special__dret_, dispatch_pkt_r_special__mret_, dispatch_pkt_r_special__sret_, dispatch_pkt_r_special__wfi_, dispatch_pkt_r_special__csrw_ })
  );


  bp_be_fp_unbox_00
  frs1_unbox
  (
    .reg_i({ dispatch_pkt_r_rs1__65_, dispatch_pkt_r_rs1__64_, dispatch_pkt_r_rs1__63_, dispatch_pkt_r_rs1__62_, dispatch_pkt_r_rs1__61_, dispatch_pkt_r_rs1__60_, dispatch_pkt_r_rs1__59_, dispatch_pkt_r_rs1__58_, dispatch_pkt_r_rs1__57_, dispatch_pkt_r_rs1__56_, dispatch_pkt_r_rs1__55_, dispatch_pkt_r_rs1__54_, dispatch_pkt_r_rs1__53_, dispatch_pkt_r_rs1__52_, dispatch_pkt_r_rs1__51_, dispatch_pkt_r_rs1__50_, dispatch_pkt_r_rs1__49_, dispatch_pkt_r_rs1__48_, dispatch_pkt_r_rs1__47_, dispatch_pkt_r_rs1__46_, dispatch_pkt_r_rs1__45_, dispatch_pkt_r_rs1__44_, dispatch_pkt_r_rs1__43_, dispatch_pkt_r_rs1__42_, dispatch_pkt_r_rs1__41_, dispatch_pkt_r_rs1__40_, dispatch_pkt_r_rs1__39_, dispatch_pkt_r_rs1__38_, dispatch_pkt_r_rs1__37_, dispatch_pkt_r_rs1__36_, dispatch_pkt_r_rs1__35_, dispatch_pkt_r_rs1__34_, dispatch_pkt_r_rs1__33_, dispatch_pkt_r_rs1__32_, dispatch_pkt_r_rs1__31_, dispatch_pkt_r_rs1__30_, dispatch_pkt_r_rs1__29_, dispatch_pkt_r_rs1__28_, dispatch_pkt_r_rs1__27_, dispatch_pkt_r_rs1__26_, dispatch_pkt_r_rs1__25_, dispatch_pkt_r_rs1__24_, dispatch_pkt_r_rs1__23_, dispatch_pkt_r_rs1__22_, dispatch_pkt_r_rs1__21_, dispatch_pkt_r_rs1__20_, dispatch_pkt_r_rs1__19_, dispatch_pkt_r_rs1__18_, dispatch_pkt_r_rs1__17_, dispatch_pkt_r_rs1__16_, dispatch_pkt_r_rs1__15_, dispatch_pkt_r_rs1__14_, dispatch_pkt_r_rs1__13_, dispatch_pkt_r_rs1__12_, dispatch_pkt_r_rs1__11_, dispatch_pkt_r_rs1__10_, dispatch_pkt_r_rs1__9_, dispatch_pkt_r_rs1__8_, dispatch_pkt_r_rs1__7_, dispatch_pkt_r_rs1__6_, dispatch_pkt_r_rs1__5_, dispatch_pkt_r_rs1__4_, dispatch_pkt_r_rs1__3_, dispatch_pkt_r_rs1__2_, dispatch_pkt_r_rs1__1_, dispatch_pkt_r_rs1__0_ }),
    .tag_i(reservation_o[412]),
    .raw_i(reservation_o[420]),
    .val_o(reservation_o[194:130])
  );


  bp_be_fp_unbox_00
  frs2_unbox
  (
    .reg_i({ dispatch_pkt_r_rs2__65_, dispatch_pkt_r_rs2__64_, dispatch_pkt_r_rs2__63_, dispatch_pkt_r_rs2__62_, dispatch_pkt_r_rs2__61_, dispatch_pkt_r_rs2__60_, dispatch_pkt_r_rs2__59_, dispatch_pkt_r_rs2__58_, dispatch_pkt_r_rs2__57_, dispatch_pkt_r_rs2__56_, dispatch_pkt_r_rs2__55_, dispatch_pkt_r_rs2__54_, dispatch_pkt_r_rs2__53_, dispatch_pkt_r_rs2__52_, dispatch_pkt_r_rs2__51_, dispatch_pkt_r_rs2__50_, dispatch_pkt_r_rs2__49_, dispatch_pkt_r_rs2__48_, dispatch_pkt_r_rs2__47_, dispatch_pkt_r_rs2__46_, dispatch_pkt_r_rs2__45_, dispatch_pkt_r_rs2__44_, dispatch_pkt_r_rs2__43_, dispatch_pkt_r_rs2__42_, dispatch_pkt_r_rs2__41_, dispatch_pkt_r_rs2__40_, dispatch_pkt_r_rs2__39_, dispatch_pkt_r_rs2__38_, dispatch_pkt_r_rs2__37_, dispatch_pkt_r_rs2__36_, dispatch_pkt_r_rs2__35_, dispatch_pkt_r_rs2__34_, dispatch_pkt_r_rs2__33_, dispatch_pkt_r_rs2__32_, dispatch_pkt_r_rs2__31_, dispatch_pkt_r_rs2__30_, dispatch_pkt_r_rs2__29_, dispatch_pkt_r_rs2__28_, dispatch_pkt_r_rs2__27_, dispatch_pkt_r_rs2__26_, dispatch_pkt_r_rs2__25_, dispatch_pkt_r_rs2__24_, dispatch_pkt_r_rs2__23_, dispatch_pkt_r_rs2__22_, dispatch_pkt_r_rs2__21_, dispatch_pkt_r_rs2__20_, dispatch_pkt_r_rs2__19_, dispatch_pkt_r_rs2__18_, dispatch_pkt_r_rs2__17_, dispatch_pkt_r_rs2__16_, dispatch_pkt_r_rs2__15_, dispatch_pkt_r_rs2__14_, dispatch_pkt_r_rs2__13_, dispatch_pkt_r_rs2__12_, dispatch_pkt_r_rs2__11_, dispatch_pkt_r_rs2__10_, dispatch_pkt_r_rs2__9_, dispatch_pkt_r_rs2__8_, dispatch_pkt_r_rs2__7_, dispatch_pkt_r_rs2__6_, dispatch_pkt_r_rs2__5_, dispatch_pkt_r_rs2__4_, dispatch_pkt_r_rs2__3_, dispatch_pkt_r_rs2__2_, dispatch_pkt_r_rs2__1_, dispatch_pkt_r_rs2__0_ }),
    .tag_i(reservation_o[411]),
    .raw_i(reservation_o[420]),
    .val_o(reservation_o[129:65])
  );


  bp_be_fp_unbox_00
  frs3_unbox
  (
    .reg_i({ dispatch_pkt_r_imm__65_, reservation_o[259:195] }),
    .tag_i(reservation_o[410]),
    .raw_i(reservation_o[420]),
    .val_o(reservation_o[64:0])
  );


  bp_be_int_unbox_00
  irs1_unbox
  (
    .reg_i({ dispatch_pkt_r_rs1__65_, dispatch_pkt_r_rs1__64_, dispatch_pkt_r_rs1__63_, dispatch_pkt_r_rs1__62_, dispatch_pkt_r_rs1__61_, dispatch_pkt_r_rs1__60_, dispatch_pkt_r_rs1__59_, dispatch_pkt_r_rs1__58_, dispatch_pkt_r_rs1__57_, dispatch_pkt_r_rs1__56_, dispatch_pkt_r_rs1__55_, dispatch_pkt_r_rs1__54_, dispatch_pkt_r_rs1__53_, dispatch_pkt_r_rs1__52_, dispatch_pkt_r_rs1__51_, dispatch_pkt_r_rs1__50_, dispatch_pkt_r_rs1__49_, dispatch_pkt_r_rs1__48_, dispatch_pkt_r_rs1__47_, dispatch_pkt_r_rs1__46_, dispatch_pkt_r_rs1__45_, dispatch_pkt_r_rs1__44_, dispatch_pkt_r_rs1__43_, dispatch_pkt_r_rs1__42_, dispatch_pkt_r_rs1__41_, dispatch_pkt_r_rs1__40_, dispatch_pkt_r_rs1__39_, dispatch_pkt_r_rs1__38_, dispatch_pkt_r_rs1__37_, dispatch_pkt_r_rs1__36_, dispatch_pkt_r_rs1__35_, dispatch_pkt_r_rs1__34_, dispatch_pkt_r_rs1__33_, dispatch_pkt_r_rs1__32_, dispatch_pkt_r_rs1__31_, dispatch_pkt_r_rs1__30_, dispatch_pkt_r_rs1__29_, dispatch_pkt_r_rs1__28_, dispatch_pkt_r_rs1__27_, dispatch_pkt_r_rs1__26_, dispatch_pkt_r_rs1__25_, dispatch_pkt_r_rs1__24_, dispatch_pkt_r_rs1__23_, dispatch_pkt_r_rs1__22_, dispatch_pkt_r_rs1__21_, dispatch_pkt_r_rs1__20_, dispatch_pkt_r_rs1__19_, dispatch_pkt_r_rs1__18_, dispatch_pkt_r_rs1__17_, dispatch_pkt_r_rs1__16_, dispatch_pkt_r_rs1__15_, dispatch_pkt_r_rs1__14_, dispatch_pkt_r_rs1__13_, dispatch_pkt_r_rs1__12_, dispatch_pkt_r_rs1__11_, dispatch_pkt_r_rs1__10_, dispatch_pkt_r_rs1__9_, dispatch_pkt_r_rs1__8_, dispatch_pkt_r_rs1__7_, dispatch_pkt_r_rs1__6_, dispatch_pkt_r_rs1__5_, dispatch_pkt_r_rs1__4_, dispatch_pkt_r_rs1__3_, dispatch_pkt_r_rs1__2_, dispatch_pkt_r_rs1__1_, dispatch_pkt_r_rs1__0_ }),
    .tag_i(reservation_o[417:416]),
    .unsigned_i(reservation_o[418]),
    .val_o(reservation_o[389:325])
  );


  bp_be_int_unbox_00
  irs2_unbox
  (
    .reg_i({ dispatch_pkt_r_rs2__65_, dispatch_pkt_r_rs2__64_, dispatch_pkt_r_rs2__63_, dispatch_pkt_r_rs2__62_, dispatch_pkt_r_rs2__61_, dispatch_pkt_r_rs2__60_, dispatch_pkt_r_rs2__59_, dispatch_pkt_r_rs2__58_, dispatch_pkt_r_rs2__57_, dispatch_pkt_r_rs2__56_, dispatch_pkt_r_rs2__55_, dispatch_pkt_r_rs2__54_, dispatch_pkt_r_rs2__53_, dispatch_pkt_r_rs2__52_, dispatch_pkt_r_rs2__51_, dispatch_pkt_r_rs2__50_, dispatch_pkt_r_rs2__49_, dispatch_pkt_r_rs2__48_, dispatch_pkt_r_rs2__47_, dispatch_pkt_r_rs2__46_, dispatch_pkt_r_rs2__45_, dispatch_pkt_r_rs2__44_, dispatch_pkt_r_rs2__43_, dispatch_pkt_r_rs2__42_, dispatch_pkt_r_rs2__41_, dispatch_pkt_r_rs2__40_, dispatch_pkt_r_rs2__39_, dispatch_pkt_r_rs2__38_, dispatch_pkt_r_rs2__37_, dispatch_pkt_r_rs2__36_, dispatch_pkt_r_rs2__35_, dispatch_pkt_r_rs2__34_, dispatch_pkt_r_rs2__33_, dispatch_pkt_r_rs2__32_, dispatch_pkt_r_rs2__31_, dispatch_pkt_r_rs2__30_, dispatch_pkt_r_rs2__29_, dispatch_pkt_r_rs2__28_, dispatch_pkt_r_rs2__27_, dispatch_pkt_r_rs2__26_, dispatch_pkt_r_rs2__25_, dispatch_pkt_r_rs2__24_, dispatch_pkt_r_rs2__23_, dispatch_pkt_r_rs2__22_, dispatch_pkt_r_rs2__21_, dispatch_pkt_r_rs2__20_, dispatch_pkt_r_rs2__19_, dispatch_pkt_r_rs2__18_, dispatch_pkt_r_rs2__17_, dispatch_pkt_r_rs2__16_, dispatch_pkt_r_rs2__15_, dispatch_pkt_r_rs2__14_, dispatch_pkt_r_rs2__13_, dispatch_pkt_r_rs2__12_, dispatch_pkt_r_rs2__11_, dispatch_pkt_r_rs2__10_, dispatch_pkt_r_rs2__9_, dispatch_pkt_r_rs2__8_, dispatch_pkt_r_rs2__7_, dispatch_pkt_r_rs2__6_, dispatch_pkt_r_rs2__5_, dispatch_pkt_r_rs2__4_, dispatch_pkt_r_rs2__3_, dispatch_pkt_r_rs2__2_, dispatch_pkt_r_rs2__1_, dispatch_pkt_r_rs2__0_ }),
    .tag_i(reservation_o[414:413]),
    .unsigned_i(reservation_o[415]),
    .val_o(reservation_o[324:260])
  );


endmodule



module bsg_dff_reset_width_p12
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [11:0] data_i;
  output [11:0] data_o;
  input clk_i;
  input reset_i;
  wire [11:0] data_o;
  reg data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,
  data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_width_p40
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [39:0] data_i;
  output [39:0] data_o;
  input clk_i;
  input reset_i;
  wire [39:0] data_o;
  reg data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,
  data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,
  data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,
  data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,
  data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_39_sv2v_reg <= 1'b0;
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_width_p64
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [63:0] data_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  wire [63:0] data_o;
  reg data_o_63_sv2v_reg,data_o_62_sv2v_reg,data_o_61_sv2v_reg,data_o_60_sv2v_reg,
  data_o_59_sv2v_reg,data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,
  data_o_55_sv2v_reg,data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,
  data_o_51_sv2v_reg,data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,
  data_o_47_sv2v_reg,data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,data_o_43_sv2v_reg,
  data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,
  data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,
  data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,
  data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,
  data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,
  data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,
  data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_63_sv2v_reg <= 1'b0;
      data_o_62_sv2v_reg <= 1'b0;
      data_o_61_sv2v_reg <= 1'b0;
      data_o_60_sv2v_reg <= 1'b0;
      data_o_59_sv2v_reg <= 1'b0;
      data_o_58_sv2v_reg <= 1'b0;
      data_o_57_sv2v_reg <= 1'b0;
      data_o_56_sv2v_reg <= 1'b0;
      data_o_55_sv2v_reg <= 1'b0;
      data_o_54_sv2v_reg <= 1'b0;
      data_o_53_sv2v_reg <= 1'b0;
      data_o_52_sv2v_reg <= 1'b0;
      data_o_51_sv2v_reg <= 1'b0;
      data_o_50_sv2v_reg <= 1'b0;
      data_o_49_sv2v_reg <= 1'b0;
      data_o_48_sv2v_reg <= 1'b0;
      data_o_47_sv2v_reg <= 1'b0;
      data_o_46_sv2v_reg <= 1'b0;
      data_o_45_sv2v_reg <= 1'b0;
      data_o_44_sv2v_reg <= 1'b0;
      data_o_43_sv2v_reg <= 1'b0;
      data_o_42_sv2v_reg <= 1'b0;
      data_o_41_sv2v_reg <= 1'b0;
      data_o_40_sv2v_reg <= 1'b0;
      data_o_39_sv2v_reg <= 1'b0;
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_width_p15
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [14:0] data_i;
  output [14:0] data_o;
  input clk_i;
  input reset_i;
  wire [14:0] data_o;
  reg data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_width_p13
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [12:0] data_i;
  output [12:0] data_o;
  input clk_i;
  input reset_i;
  wire [12:0] data_o;
  reg data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,
  data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,
  data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_width_p3
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [2:0] data_i;
  output [2:0] data_o;
  input clk_i;
  input reset_i;
  wire [2:0] data_o;
  reg data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_width_p6
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [5:0] data_i;
  output [5:0] data_o;
  input clk_i;
  input reset_i;
  wire [5:0] data_o;
  reg data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_width_p38
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [37:0] data_i;
  output [37:0] data_o;
  input clk_i;
  input reset_i;
  wire [37:0] data_o;
  reg data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,
  data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,
  data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,
  data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,
  data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,
  data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,
  data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,
  data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_width_p2
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [1:0] data_i;
  output [1:0] data_o;
  input clk_i;
  input reset_i;
  wire [1:0] data_o;
  reg data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_width_p5
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [4:0] data_i;
  output [4:0] data_o;
  input clk_i;
  input reset_i;
  wire [4:0] data_o;
  reg data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_width_p48
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [47:0] data_i;
  output [47:0] data_o;
  input clk_i;
  input reset_i;
  wire [47:0] data_o;
  reg data_o_47_sv2v_reg,data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,
  data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,
  data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,
  data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,
  data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,
  data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,
  data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,
  data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,
  data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_47_sv2v_reg <= 1'b0;
      data_o_46_sv2v_reg <= 1'b0;
      data_o_45_sv2v_reg <= 1'b0;
      data_o_44_sv2v_reg <= 1'b0;
      data_o_43_sv2v_reg <= 1'b0;
      data_o_42_sv2v_reg <= 1'b0;
      data_o_41_sv2v_reg <= 1'b0;
      data_o_40_sv2v_reg <= 1'b0;
      data_o_39_sv2v_reg <= 1'b0;
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_width_p29
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [28:0] data_i;
  output [28:0] data_o;
  input clk_i;
  input reset_i;
  wire [28:0] data_o;
  reg data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,
  data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,
  data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,
  data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,
  data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,
  data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_width_p8
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [7:0] data_i;
  output [7:0] data_o;
  input clk_i;
  input reset_i;
  wire [7:0] data_o;
  reg data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_scan_width_p16_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [15:0] i;
  output [15:0] o;
  wire [15:0] o;
  wire t_3__15_,t_3__14_,t_3__13_,t_3__12_,t_3__11_,t_3__10_,t_3__9_,t_3__8_,t_3__7_,
  t_3__6_,t_3__5_,t_3__4_,t_3__3_,t_3__2_,t_3__1_,t_3__0_,t_2__15_,t_2__14_,
  t_2__13_,t_2__12_,t_2__11_,t_2__10_,t_2__9_,t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,
  t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__15_,t_1__14_,t_1__13_,t_1__12_,t_1__11_,
  t_1__10_,t_1__9_,t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,
  t_1__0_;
  assign t_1__15_ = i[0] | 1'b0;
  assign t_1__14_ = i[1] | i[0];
  assign t_1__13_ = i[2] | i[1];
  assign t_1__12_ = i[3] | i[2];
  assign t_1__11_ = i[4] | i[3];
  assign t_1__10_ = i[5] | i[4];
  assign t_1__9_ = i[6] | i[5];
  assign t_1__8_ = i[7] | i[6];
  assign t_1__7_ = i[8] | i[7];
  assign t_1__6_ = i[9] | i[8];
  assign t_1__5_ = i[10] | i[9];
  assign t_1__4_ = i[11] | i[10];
  assign t_1__3_ = i[12] | i[11];
  assign t_1__2_ = i[13] | i[12];
  assign t_1__1_ = i[14] | i[13];
  assign t_1__0_ = i[15] | i[14];
  assign t_2__15_ = t_1__15_ | 1'b0;
  assign t_2__14_ = t_1__14_ | 1'b0;
  assign t_2__13_ = t_1__13_ | t_1__15_;
  assign t_2__12_ = t_1__12_ | t_1__14_;
  assign t_2__11_ = t_1__11_ | t_1__13_;
  assign t_2__10_ = t_1__10_ | t_1__12_;
  assign t_2__9_ = t_1__9_ | t_1__11_;
  assign t_2__8_ = t_1__8_ | t_1__10_;
  assign t_2__7_ = t_1__7_ | t_1__9_;
  assign t_2__6_ = t_1__6_ | t_1__8_;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign t_3__15_ = t_2__15_ | 1'b0;
  assign t_3__14_ = t_2__14_ | 1'b0;
  assign t_3__13_ = t_2__13_ | 1'b0;
  assign t_3__12_ = t_2__12_ | 1'b0;
  assign t_3__11_ = t_2__11_ | t_2__15_;
  assign t_3__10_ = t_2__10_ | t_2__14_;
  assign t_3__9_ = t_2__9_ | t_2__13_;
  assign t_3__8_ = t_2__8_ | t_2__12_;
  assign t_3__7_ = t_2__7_ | t_2__11_;
  assign t_3__6_ = t_2__6_ | t_2__10_;
  assign t_3__5_ = t_2__5_ | t_2__9_;
  assign t_3__4_ = t_2__4_ | t_2__8_;
  assign t_3__3_ = t_2__3_ | t_2__7_;
  assign t_3__2_ = t_2__2_ | t_2__6_;
  assign t_3__1_ = t_2__1_ | t_2__5_;
  assign t_3__0_ = t_2__0_ | t_2__4_;
  assign o[0] = t_3__15_ | 1'b0;
  assign o[1] = t_3__14_ | 1'b0;
  assign o[2] = t_3__13_ | 1'b0;
  assign o[3] = t_3__12_ | 1'b0;
  assign o[4] = t_3__11_ | 1'b0;
  assign o[5] = t_3__10_ | 1'b0;
  assign o[6] = t_3__9_ | 1'b0;
  assign o[7] = t_3__8_ | 1'b0;
  assign o[8] = t_3__7_ | t_3__15_;
  assign o[9] = t_3__6_ | t_3__14_;
  assign o[10] = t_3__5_ | t_3__13_;
  assign o[11] = t_3__4_ | t_3__12_;
  assign o[12] = t_3__3_ | t_3__11_;
  assign o[13] = t_3__2_ | t_3__10_;
  assign o[14] = t_3__1_ | t_3__9_;
  assign o[15] = t_3__0_ | t_3__8_;

endmodule



module bsg_priority_encode_one_hot_out_width_p16_lo_to_hi_p1
(
  i,
  o,
  v_o
);

  input [15:0] i;
  output [15:0] o;
  output v_o;
  wire [15:0] o;
  wire v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;
  wire [14:1] scan_lo;

  bsg_scan_width_p16_or_p1_lo_to_hi_p1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, scan_lo, o[0:0] })
  );

  assign o[15] = v_o & N0;
  assign N0 = ~scan_lo[14];
  assign o[14] = scan_lo[14] & N1;
  assign N1 = ~scan_lo[13];
  assign o[13] = scan_lo[13] & N2;
  assign N2 = ~scan_lo[12];
  assign o[12] = scan_lo[12] & N3;
  assign N3 = ~scan_lo[11];
  assign o[11] = scan_lo[11] & N4;
  assign N4 = ~scan_lo[10];
  assign o[10] = scan_lo[10] & N5;
  assign N5 = ~scan_lo[9];
  assign o[9] = scan_lo[9] & N6;
  assign N6 = ~scan_lo[8];
  assign o[8] = scan_lo[8] & N7;
  assign N7 = ~scan_lo[7];
  assign o[7] = scan_lo[7] & N8;
  assign N8 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N9;
  assign N9 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N10;
  assign N10 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N11;
  assign N11 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N12;
  assign N12 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N13;
  assign N13 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N14;
  assign N14 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p16_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [15:0] i;
  output [3:0] addr_o;
  output v_o;
  wire [3:0] addr_o;
  wire v_o,v_3__0_,v_2__12_,v_2__8_,v_2__4_,v_2__0_,v_1__14_,v_1__12_,v_1__10_,v_1__8_,
  v_1__6_,v_1__4_,v_1__2_,v_1__0_,addr_3__9_,addr_3__8_,addr_3__1_,addr_3__0_,
  addr_2__12_,addr_2__8_,addr_2__4_,addr_2__0_;
  assign v_1__0_ = i[1] | i[0];
  assign v_1__2_ = i[3] | i[2];
  assign v_1__4_ = i[5] | i[4];
  assign v_1__6_ = i[7] | i[6];
  assign v_1__8_ = i[9] | i[8];
  assign v_1__10_ = i[11] | i[10];
  assign v_1__12_ = i[13] | i[12];
  assign v_1__14_ = i[15] | i[14];
  assign v_2__0_ = v_1__2_ | v_1__0_;
  assign addr_2__0_ = i[1] | i[3];
  assign v_2__4_ = v_1__6_ | v_1__4_;
  assign addr_2__4_ = i[5] | i[7];
  assign v_2__8_ = v_1__10_ | v_1__8_;
  assign addr_2__8_ = i[9] | i[11];
  assign v_2__12_ = v_1__14_ | v_1__12_;
  assign addr_2__12_ = i[13] | i[15];
  assign v_3__0_ = v_2__4_ | v_2__0_;
  assign addr_3__1_ = v_1__2_ | v_1__6_;
  assign addr_3__0_ = addr_2__0_ | addr_2__4_;
  assign addr_o[3] = v_2__12_ | v_2__8_;
  assign addr_3__9_ = v_1__10_ | v_1__14_;
  assign addr_3__8_ = addr_2__8_ | addr_2__12_;
  assign v_o = addr_o[3] | v_3__0_;
  assign addr_o[2] = v_2__4_ | v_2__12_;
  assign addr_o[1] = addr_3__1_ | addr_3__9_;
  assign addr_o[0] = addr_3__0_ | addr_3__8_;

endmodule



module bsg_priority_encode_width_p16_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [15:0] i;
  output [3:0] addr_o;
  output v_o;
  wire [3:0] addr_o;
  wire v_o;
  wire [15:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p16_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_width_p16_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o)
  );


endmodule



module bsg_dff_reset_set_clear_width_p1
(
  clk_i,
  reset_i,
  set_i,
  clear_i,
  data_o
);

  input [0:0] set_i;
  input [0:0] clear_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  wire [0:0] data_o;
  wire N0,N1,N2;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N0 = N2 | set_i[0];
  assign N2 = data_o[0] & N1;
  assign N1 = ~clear_i[0];

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_0_sv2v_reg <= N0;
    end 
  end


endmodule



module bsg_dff_reset_00000027
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [38:0] data_i;
  output [38:0] data_o;
  input clk_i;
  input reset_i;
  wire [38:0] data_o;
  reg data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,
  data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,
  data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,
  data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,
  data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,
  data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_00000027
(
  clk_i,
  data_i,
  data_o
);

  input [38:0] data_i;
  output [38:0] data_o;
  input clk_i;
  wire [38:0] data_o;
  reg data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,
  data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,
  data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,
  data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,
  data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,
  data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_3_3
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [2:0] data_i;
  output [2:0] data_o;
  input clk_i;
  input reset_i;
  wire [2:0] data_o;
  reg data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b1;
      data_o_0_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bp_be_csr_00
(
  clk_i,
  reset_i,
  cfg_bus_i,
  csr_r_v_i,
  csr_r_addr_i,
  csr_r_data_o,
  csr_r_illegal_o,
  retire_pkt_i,
  frf_w_v_i,
  debug_irq_i,
  timer_irq_i,
  software_irq_i,
  m_external_irq_i,
  s_external_irq_i,
  irq_pending_o,
  irq_waiting_o,
  commit_pkt_o,
  decode_info_o,
  trans_info_o,
  frm_dyn_o,
  fflags_acc_i_nv_,
  fflags_acc_i_dz_,
  fflags_acc_i_of_,
  fflags_acc_i_uf_,
  fflags_acc_i_nx_
);

  input [60:0] cfg_bus_i;
  input [11:0] csr_r_addr_i;
  output [63:0] csr_r_data_o;
  input [219:0] retire_pkt_i;
  output [213:0] commit_pkt_o;
  output [12:0] decode_info_o;
  output [32:0] trans_info_o;
  output [2:0] frm_dyn_o;
  input clk_i;
  input reset_i;
  input csr_r_v_i;
  input frf_w_v_i;
  input debug_irq_i;
  input timer_irq_i;
  input software_irq_i;
  input m_external_irq_i;
  input s_external_irq_i;
  input fflags_acc_i_nv_;
  input fflags_acc_i_dz_;
  input fflags_acc_i_of_;
  input fflags_acc_i_uf_;
  input fflags_acc_i_nx_;
  output csr_r_illegal_o;
  output irq_pending_o;
  output irq_waiting_o;
  wire [63:0] csr_r_data_o,dscratch0_n,dscratch0_r,dscratch1_n,dscratch1_r,mscratch_n,
  mscratch_r,sstatus_lo,sie_lo,sscratch_n,sscratch_r,sip_lo;
  wire [213:0] commit_pkt_o;
  wire [12:0] decode_info_o,medeleg_n,medeleg_r;
  wire [32:0] trans_info_o;
  wire [2:0] frm_dyn_o;
  wire csr_r_illegal_o,irq_pending_o,irq_waiting_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,
  N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,
  N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,
  N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,
  N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,
  N91,N92,N93,N94,N95,N96,N97,N98,commit_pkt_o_211_,commit_pkt_o_210_,
  commit_pkt_o_209_,commit_pkt_o_208_,commit_pkt_o_207_,commit_pkt_o_206_,commit_pkt_o_127_,
  commit_pkt_o_126_,commit_pkt_o_125_,commit_pkt_o_124_,commit_pkt_o_123_,
  commit_pkt_o_122_,commit_pkt_o_121_,commit_pkt_o_120_,commit_pkt_o_119_,commit_pkt_o_118_,
  commit_pkt_o_117_,commit_pkt_o_116_,commit_pkt_o_115_,commit_pkt_o_114_,
  commit_pkt_o_113_,commit_pkt_o_112_,commit_pkt_o_111_,commit_pkt_o_110_,commit_pkt_o_109_,
  commit_pkt_o_108_,commit_pkt_o_107_,commit_pkt_o_106_,commit_pkt_o_105_,
  commit_pkt_o_104_,commit_pkt_o_103_,commit_pkt_o_102_,commit_pkt_o_101_,
  commit_pkt_o_100_,commit_pkt_o_99_,commit_pkt_o_98_,commit_pkt_o_97_,commit_pkt_o_96_,
  commit_pkt_o_95_,commit_pkt_o_94_,commit_pkt_o_93_,commit_pkt_o_92_,commit_pkt_o_91_,
  commit_pkt_o_90_,commit_pkt_o_89_,commit_pkt_o_88_,commit_pkt_o_87_,commit_pkt_o_86_,
  commit_pkt_o_85_,commit_pkt_o_84_,commit_pkt_o_83_,commit_pkt_o_82_,
  commit_pkt_o_81_,commit_pkt_o_80_,commit_pkt_o_79_,commit_pkt_o_78_,commit_pkt_o_77_,
  commit_pkt_o_76_,commit_pkt_o_75_,commit_pkt_o_74_,commit_pkt_o_73_,commit_pkt_o_72_,
  commit_pkt_o_71_,commit_pkt_o_70_,commit_pkt_o_69_,commit_pkt_o_68_,
  commit_pkt_o_67_,commit_pkt_o_66_,commit_pkt_o_65_,commit_pkt_o_64_,commit_pkt_o_63_,
  commit_pkt_o_62_,commit_pkt_o_61_,commit_pkt_o_60_,commit_pkt_o_59_,commit_pkt_o_58_,
  commit_pkt_o_57_,commit_pkt_o_56_,commit_pkt_o_55_,commit_pkt_o_54_,
  commit_pkt_o_53_,commit_pkt_o_52_,commit_pkt_o_51_,commit_pkt_o_50_,commit_pkt_o_49_,
  commit_pkt_o_48_,commit_pkt_o_47_,commit_pkt_o_46_,commit_pkt_o_45_,commit_pkt_o_44_,
  commit_pkt_o_43_,commit_pkt_o_42_,commit_pkt_o_41_,commit_pkt_o_40_,commit_pkt_o_39_,
  commit_pkt_o_38_,commit_pkt_o_37_,commit_pkt_o_36_,commit_pkt_o_35_,
  commit_pkt_o_34_,commit_pkt_o_33_,commit_pkt_o_32_,commit_pkt_o_31_,commit_pkt_o_30_,
  commit_pkt_o_29_,commit_pkt_o_28_,commit_pkt_o_27_,commit_pkt_o_26_,commit_pkt_o_25_,
  commit_pkt_o_24_,commit_pkt_o_23_,commit_pkt_o_22_,commit_pkt_o_21_,
  commit_pkt_o_15_,commit_pkt_o_13_,commit_pkt_o_12_,commit_pkt_o_11_,commit_pkt_o_10_,
  commit_pkt_o_9_,commit_pkt_o_8_,commit_pkt_o_7_,commit_pkt_o_6_,commit_pkt_o_5_,
  commit_pkt_o_4_,commit_pkt_o_3_,commit_pkt_o_2_,commit_pkt_o_1_,commit_pkt_o_0_,
  decode_info_o_5_,dcsr_r_ebreaks_,dcsr_r_ebreaku_,dcsr_r_stepie_,dcsr_r_cause__3_,
  dcsr_r_cause__2_,dcsr_r_cause__1_,dcsr_r_cause__0_,dcsr_r_prv__1_,dcsr_r_prv__0_,
  dcsr_r_mprven_,dcsr_r_step_,mstatus_r_mprv_,mstatus_r_fs__1_,mstatus_r_fs__0_,
  mstatus_r_mpp__1_,mstatus_r_mpp__0_,mstatus_r_spp_,mstatus_r_mpie_,mstatus_r_spie_,
  mstatus_r_mie_,mstatus_r_sie_,mideleg_n_sei_,mideleg_n_sti_,mideleg_n_ssi_,
  mideleg_r_sei_,mideleg_r_sti_,mideleg_r_ssi_,mie_n_meie_,mie_n_seie_,mie_n_mtie_,
  mie_n_stie_,mie_n_msie_,mie_n_ssie_,mie_r_meie_,mie_r_seie_,mie_r_mtie_,mie_r_stie_,
  mie_r_msie_,mie_r_ssie_,mcounteren_n_ir_,mcounteren_n_cy_,mcounteren_r_ir_,
  mcounteren_r_cy_,mip_n_seip_,mip_n_stip_,mip_n_ssip_,mip_r_meip_,mip_r_seip_,mip_r_mtip_,
  mip_r_stip_,mip_r_msip_,mip_r_ssip_,mcountinhibit_n_ir_,mcountinhibit_n_cy_,
  mcountinhibit_r_ir_,mcountinhibit_r_cy_,scounteren_n_ir_,scounteren_n_cy_,
  scounteren_r_ir_,scounteren_r_cy_,satp_r_mode_,satp_li_mode__2_,satp_li_mode__1_,
  satp_li_mode__0_,fcsr_r_fflags__4_,fcsr_r_fflags__3_,fcsr_r_fflags__2_,fcsr_r_fflags__1_,
  fcsr_r_fflags__0_,dgie,mgie,sgie,interrupt_icode_dec_li_9,interrupt_icode_dec_li_7,
  interrupt_icode_dec_li_5,interrupt_icode_dec_li_3,interrupt_icode_dec_li_1,
  exception_ecode_v_li,_0_net__15_,_0_net__14_,_0_net__13_,_0_net__12_,_0_net__11_,
  _0_net__10_,_0_net__9_,_0_net__8_,_0_net__7_,_0_net__6_,_0_net__5_,_0_net__4_,
  _0_net__3_,_0_net__2_,_0_net__1_,_0_net__0_,m_interrupt_icode_v_li,_1_net__15_,
  _1_net__14_,_1_net__13_,_1_net__12_,_1_net__11_,_1_net__10_,_1_net__9_,_1_net__8_,
  _1_net__7_,_1_net__6_,_1_net__5_,_1_net__4_,_1_net__3_,_1_net__2_,_1_net__1_,
  _1_net__0_,s_interrupt_icode_v_li,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,
  N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,
  N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,csr_fany_li,N138,
  N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,
  N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,
  N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,instr_fany_li,enter_debug,
  exit_debug,N182,N183,N184,N185,N186,N187,N188,N189,interrupt_v_lo,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,translation_en_r,N202,N203,N204,
  N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,
  N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,
  N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,
  N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,
  N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,
  N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,
  N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,
  N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,
  N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
  N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,
  N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,
  N381,N382,csr_data_lo_9,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,
  N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,
  N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,
  N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,
  N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,
  N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,
  N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,
  N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,
  N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,
  N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,
  N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,
  N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,
  N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,
  N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,
  N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,
  N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,
  N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,
  N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,
  N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,
  N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,
  N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,
  N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,
  N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,
  N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,
  N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,
  N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,
  N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,
  N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,
  N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,
  N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,
  N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,
  N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,
  N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,
  N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,
  N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,
  N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,
  N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,
  N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,
  N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,
  N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,
  N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,
  N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,
  N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,
  N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,
  N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,
  N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,
  N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,
  N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,
  N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,
  N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,
  N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,
  N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,
  N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,
  N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,
  N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,
  N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,
  N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,
  N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,
  N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,
  N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,
  N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,
  N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,
  N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,
  N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,
  N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,
  N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,
  N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,
  N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,
  N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,
  N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,
  N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,
  N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,
  N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,
  N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,
  N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,
  N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,
  N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,
  N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,
  N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,
  N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,
  N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,
  N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,
  N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,
  N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,
  N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,
  N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,
  N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,
  N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,
  N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,
  N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,
  N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,
  N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,
  N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,
  N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734,
  N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,
  N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760,N1761,
  N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,N1771,N1772,N1773,N1774,
  N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,
  N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,
  N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814,
  N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,
  N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,N1838,N1839,N1840,N1841,
  N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,
  N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,
  N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,
  N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,N1891,N1892,N1893,N1894,
  N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,
  N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,N1919,N1920,N1921,
  N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,
  N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,
  N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,N1958,N1959,N1960,N1961,
  N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,
  N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,
  N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,N1998,N1999,N2000,N2001,
  N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,
  N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,
  N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,N2038,N2039,N2040,N2041,
  N2042,N2043,N2044,N2045,N2046,N2048,N2049,N2050,N2051,N2052,N2053,N2054,N2055,
  N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2069,N2071,
  N2072,N2073,N2074,N2075,N2076,N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,
  N2085,N2086,N2087,N2088,N2089,N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,
  N2098,N2099,N2100,N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,
  N2112,N2113,N2114,N2115,N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,
  N2125,N2126,N2127,N2128,N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,
  N2138,N2139,N2140,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,
  N2152,N2153,N2154,N2155,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,
  N2165,N2166,N2167,N2168,N2169,N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,
  N2178,N2179,N2180,N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,
  N2192,N2193,N2194,N2195,N2196,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,
  N2205,N2206,N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,
  N2218,N2219,N2220,N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,
  N2232,N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,
  N2245,N2246,N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,
  N2258,N2259,N2260,N2261;
  wire [11:0] dcsr_n;
  wire [39:0] dpc_n,dpc_r,mepc_n,mepc_r,mtval_n,mtval_r,sepc_n,sepc_r,stval_n,stval_r;
  wire [14:0] mstatus_n;
  wire [37:0] mtvec_n,mtvec_r,stvec_n,stvec_r;
  wire [4:0] mcause_n,mcause_r,scause_n,scause_r,csr_data_lo;
  wire [47:0] mcycle_n,mcycle_r,minstret_n,minstret_r;
  wire [28:0] satp_n;
  wire [7:0] fcsr_n;
  wire [11:11] interrupt_icode_dec_li;
  wire [3:0] exception_ecode_li,m_interrupt_icode_li,s_interrupt_icode_li;
  wire [38:0] cfg_npc_r,ret_pc,core_npc;
  wire [38:2] tvec_pc;
  assign commit_pkt_o_211_ = retire_pkt_i[217];
  assign commit_pkt_o[211] = commit_pkt_o_211_;
  assign commit_pkt_o_210_ = retire_pkt_i[40];
  assign commit_pkt_o[210] = commit_pkt_o_210_;
  assign commit_pkt_o_209_ = retire_pkt_i[39];
  assign commit_pkt_o[209] = commit_pkt_o_209_;
  assign commit_pkt_o_208_ = retire_pkt_i[38];
  assign commit_pkt_o[208] = commit_pkt_o_208_;
  assign commit_pkt_o_207_ = retire_pkt_i[37];
  assign commit_pkt_o[207] = commit_pkt_o_207_;
  assign commit_pkt_o_206_ = retire_pkt_i[36];
  assign commit_pkt_o[206] = commit_pkt_o_206_;
  assign commit_pkt_o_127_ = retire_pkt_i[177];
  assign commit_pkt_o[127] = commit_pkt_o_127_;
  assign commit_pkt_o_126_ = retire_pkt_i[176];
  assign commit_pkt_o[126] = commit_pkt_o_126_;
  assign commit_pkt_o_125_ = retire_pkt_i[175];
  assign commit_pkt_o[125] = commit_pkt_o_125_;
  assign commit_pkt_o_124_ = retire_pkt_i[174];
  assign commit_pkt_o[124] = commit_pkt_o_124_;
  assign commit_pkt_o_123_ = retire_pkt_i[173];
  assign commit_pkt_o[123] = commit_pkt_o_123_;
  assign commit_pkt_o_122_ = retire_pkt_i[172];
  assign commit_pkt_o[122] = commit_pkt_o_122_;
  assign commit_pkt_o_121_ = retire_pkt_i[171];
  assign commit_pkt_o[121] = commit_pkt_o_121_;
  assign commit_pkt_o_120_ = retire_pkt_i[170];
  assign commit_pkt_o[120] = commit_pkt_o_120_;
  assign commit_pkt_o_119_ = retire_pkt_i[169];
  assign commit_pkt_o[119] = commit_pkt_o_119_;
  assign commit_pkt_o_118_ = retire_pkt_i[168];
  assign commit_pkt_o[118] = commit_pkt_o_118_;
  assign commit_pkt_o_117_ = retire_pkt_i[167];
  assign commit_pkt_o[117] = commit_pkt_o_117_;
  assign commit_pkt_o_116_ = retire_pkt_i[166];
  assign commit_pkt_o[116] = commit_pkt_o_116_;
  assign commit_pkt_o_115_ = retire_pkt_i[165];
  assign commit_pkt_o[115] = commit_pkt_o_115_;
  assign commit_pkt_o_114_ = retire_pkt_i[164];
  assign commit_pkt_o[114] = commit_pkt_o_114_;
  assign commit_pkt_o_113_ = retire_pkt_i[163];
  assign commit_pkt_o[113] = commit_pkt_o_113_;
  assign commit_pkt_o_112_ = retire_pkt_i[162];
  assign commit_pkt_o[112] = commit_pkt_o_112_;
  assign commit_pkt_o_111_ = retire_pkt_i[161];
  assign commit_pkt_o[111] = commit_pkt_o_111_;
  assign commit_pkt_o_110_ = retire_pkt_i[160];
  assign commit_pkt_o[110] = commit_pkt_o_110_;
  assign commit_pkt_o_109_ = retire_pkt_i[159];
  assign commit_pkt_o[109] = commit_pkt_o_109_;
  assign commit_pkt_o_108_ = retire_pkt_i[158];
  assign commit_pkt_o[108] = commit_pkt_o_108_;
  assign commit_pkt_o_107_ = retire_pkt_i[157];
  assign commit_pkt_o[107] = commit_pkt_o_107_;
  assign commit_pkt_o_106_ = retire_pkt_i[156];
  assign commit_pkt_o[106] = commit_pkt_o_106_;
  assign commit_pkt_o_105_ = retire_pkt_i[155];
  assign commit_pkt_o[105] = commit_pkt_o_105_;
  assign commit_pkt_o_104_ = retire_pkt_i[154];
  assign commit_pkt_o[104] = commit_pkt_o_104_;
  assign commit_pkt_o_103_ = retire_pkt_i[153];
  assign commit_pkt_o[103] = commit_pkt_o_103_;
  assign commit_pkt_o_102_ = retire_pkt_i[152];
  assign commit_pkt_o[102] = commit_pkt_o_102_;
  assign commit_pkt_o_101_ = retire_pkt_i[151];
  assign commit_pkt_o[101] = commit_pkt_o_101_;
  assign commit_pkt_o_100_ = retire_pkt_i[150];
  assign commit_pkt_o[100] = commit_pkt_o_100_;
  assign commit_pkt_o_99_ = retire_pkt_i[149];
  assign commit_pkt_o[99] = commit_pkt_o_99_;
  assign commit_pkt_o_98_ = retire_pkt_i[148];
  assign commit_pkt_o[98] = commit_pkt_o_98_;
  assign commit_pkt_o_97_ = retire_pkt_i[147];
  assign commit_pkt_o[97] = commit_pkt_o_97_;
  assign commit_pkt_o_96_ = retire_pkt_i[146];
  assign commit_pkt_o[96] = commit_pkt_o_96_;
  assign commit_pkt_o_95_ = retire_pkt_i[145];
  assign commit_pkt_o[95] = commit_pkt_o_95_;
  assign commit_pkt_o_94_ = retire_pkt_i[144];
  assign commit_pkt_o[94] = commit_pkt_o_94_;
  assign commit_pkt_o_93_ = retire_pkt_i[143];
  assign commit_pkt_o[93] = commit_pkt_o_93_;
  assign commit_pkt_o_92_ = retire_pkt_i[142];
  assign commit_pkt_o[92] = commit_pkt_o_92_;
  assign commit_pkt_o_91_ = retire_pkt_i[141];
  assign commit_pkt_o[91] = commit_pkt_o_91_;
  assign commit_pkt_o_90_ = retire_pkt_i[140];
  assign commit_pkt_o[90] = commit_pkt_o_90_;
  assign commit_pkt_o_89_ = retire_pkt_i[139];
  assign commit_pkt_o[89] = commit_pkt_o_89_;
  assign commit_pkt_o_88_ = retire_pkt_i[72];
  assign commit_pkt_o[88] = commit_pkt_o_88_;
  assign commit_pkt_o_87_ = retire_pkt_i[71];
  assign commit_pkt_o[87] = commit_pkt_o_87_;
  assign commit_pkt_o_86_ = retire_pkt_i[70];
  assign commit_pkt_o[86] = commit_pkt_o_86_;
  assign commit_pkt_o_85_ = retire_pkt_i[69];
  assign commit_pkt_o[85] = commit_pkt_o_85_;
  assign commit_pkt_o_84_ = retire_pkt_i[68];
  assign commit_pkt_o[84] = commit_pkt_o_84_;
  assign commit_pkt_o_83_ = retire_pkt_i[67];
  assign commit_pkt_o[83] = commit_pkt_o_83_;
  assign commit_pkt_o_82_ = retire_pkt_i[66];
  assign commit_pkt_o[82] = commit_pkt_o_82_;
  assign commit_pkt_o_81_ = retire_pkt_i[65];
  assign commit_pkt_o[81] = commit_pkt_o_81_;
  assign commit_pkt_o_80_ = retire_pkt_i[64];
  assign commit_pkt_o[80] = commit_pkt_o_80_;
  assign commit_pkt_o_79_ = retire_pkt_i[63];
  assign commit_pkt_o[79] = commit_pkt_o_79_;
  assign commit_pkt_o_78_ = retire_pkt_i[62];
  assign commit_pkt_o[78] = commit_pkt_o_78_;
  assign commit_pkt_o_77_ = retire_pkt_i[61];
  assign commit_pkt_o[77] = commit_pkt_o_77_;
  assign commit_pkt_o_76_ = retire_pkt_i[60];
  assign commit_pkt_o[76] = commit_pkt_o_76_;
  assign commit_pkt_o_75_ = retire_pkt_i[59];
  assign commit_pkt_o[75] = commit_pkt_o_75_;
  assign commit_pkt_o_74_ = retire_pkt_i[58];
  assign commit_pkt_o[74] = commit_pkt_o_74_;
  assign commit_pkt_o_73_ = retire_pkt_i[57];
  assign commit_pkt_o[73] = commit_pkt_o_73_;
  assign commit_pkt_o_72_ = retire_pkt_i[56];
  assign commit_pkt_o[72] = commit_pkt_o_72_;
  assign commit_pkt_o_71_ = retire_pkt_i[55];
  assign commit_pkt_o[71] = commit_pkt_o_71_;
  assign commit_pkt_o_70_ = retire_pkt_i[54];
  assign commit_pkt_o[70] = commit_pkt_o_70_;
  assign commit_pkt_o_69_ = retire_pkt_i[53];
  assign commit_pkt_o[69] = commit_pkt_o_69_;
  assign commit_pkt_o_68_ = retire_pkt_i[52];
  assign commit_pkt_o[68] = commit_pkt_o_68_;
  assign commit_pkt_o_67_ = retire_pkt_i[51];
  assign commit_pkt_o[67] = commit_pkt_o_67_;
  assign commit_pkt_o_66_ = retire_pkt_i[50];
  assign commit_pkt_o[66] = commit_pkt_o_66_;
  assign commit_pkt_o_65_ = retire_pkt_i[49];
  assign commit_pkt_o[65] = commit_pkt_o_65_;
  assign commit_pkt_o_64_ = retire_pkt_i[48];
  assign commit_pkt_o[64] = commit_pkt_o_64_;
  assign commit_pkt_o_63_ = retire_pkt_i[47];
  assign commit_pkt_o[63] = commit_pkt_o_63_;
  assign commit_pkt_o_62_ = retire_pkt_i[46];
  assign commit_pkt_o[62] = commit_pkt_o_62_;
  assign commit_pkt_o_61_ = retire_pkt_i[45];
  assign commit_pkt_o[61] = commit_pkt_o_61_;
  assign commit_pkt_o_60_ = retire_pkt_i[44];
  assign commit_pkt_o[60] = commit_pkt_o_60_;
  assign commit_pkt_o_59_ = retire_pkt_i[43];
  assign commit_pkt_o[59] = commit_pkt_o_59_;
  assign commit_pkt_o_58_ = retire_pkt_i[42];
  assign commit_pkt_o[58] = commit_pkt_o_58_;
  assign commit_pkt_o_57_ = retire_pkt_i[41];
  assign commit_pkt_o[57] = commit_pkt_o_57_;
  assign commit_pkt_o_56_ = retire_pkt_i[108];
  assign commit_pkt_o[56] = commit_pkt_o_56_;
  assign commit_pkt_o_55_ = retire_pkt_i[107];
  assign commit_pkt_o[55] = commit_pkt_o_55_;
  assign commit_pkt_o_54_ = retire_pkt_i[106];
  assign commit_pkt_o[54] = commit_pkt_o_54_;
  assign commit_pkt_o_53_ = retire_pkt_i[105];
  assign commit_pkt_o[53] = commit_pkt_o_53_;
  assign commit_pkt_o_52_ = retire_pkt_i[104];
  assign commit_pkt_o[52] = commit_pkt_o_52_;
  assign commit_pkt_o_51_ = retire_pkt_i[103];
  assign commit_pkt_o[51] = commit_pkt_o_51_;
  assign commit_pkt_o_50_ = retire_pkt_i[102];
  assign commit_pkt_o[50] = commit_pkt_o_50_;
  assign commit_pkt_o_49_ = retire_pkt_i[101];
  assign commit_pkt_o[49] = commit_pkt_o_49_;
  assign commit_pkt_o_48_ = retire_pkt_i[100];
  assign commit_pkt_o[48] = commit_pkt_o_48_;
  assign commit_pkt_o_47_ = retire_pkt_i[99];
  assign commit_pkt_o[47] = commit_pkt_o_47_;
  assign commit_pkt_o_46_ = retire_pkt_i[98];
  assign commit_pkt_o[46] = commit_pkt_o_46_;
  assign commit_pkt_o_45_ = retire_pkt_i[97];
  assign commit_pkt_o[45] = commit_pkt_o_45_;
  assign commit_pkt_o_44_ = retire_pkt_i[96];
  assign commit_pkt_o[44] = commit_pkt_o_44_;
  assign commit_pkt_o_43_ = retire_pkt_i[95];
  assign commit_pkt_o[43] = commit_pkt_o_43_;
  assign commit_pkt_o_42_ = retire_pkt_i[94];
  assign commit_pkt_o[42] = commit_pkt_o_42_;
  assign commit_pkt_o_41_ = retire_pkt_i[93];
  assign commit_pkt_o[41] = commit_pkt_o_41_;
  assign commit_pkt_o_40_ = retire_pkt_i[92];
  assign commit_pkt_o[40] = commit_pkt_o_40_;
  assign commit_pkt_o_39_ = retire_pkt_i[91];
  assign commit_pkt_o[39] = commit_pkt_o_39_;
  assign commit_pkt_o_38_ = retire_pkt_i[90];
  assign commit_pkt_o[38] = commit_pkt_o_38_;
  assign commit_pkt_o_37_ = retire_pkt_i[89];
  assign commit_pkt_o[37] = commit_pkt_o_37_;
  assign commit_pkt_o_36_ = retire_pkt_i[88];
  assign commit_pkt_o[36] = commit_pkt_o_36_;
  assign commit_pkt_o_35_ = retire_pkt_i[87];
  assign commit_pkt_o[35] = commit_pkt_o_35_;
  assign commit_pkt_o_34_ = retire_pkt_i[86];
  assign commit_pkt_o[34] = commit_pkt_o_34_;
  assign commit_pkt_o_33_ = retire_pkt_i[85];
  assign commit_pkt_o[33] = commit_pkt_o_33_;
  assign commit_pkt_o_32_ = retire_pkt_i[84];
  assign commit_pkt_o[32] = commit_pkt_o_32_;
  assign commit_pkt_o_31_ = retire_pkt_i[83];
  assign commit_pkt_o[31] = commit_pkt_o_31_;
  assign commit_pkt_o_30_ = retire_pkt_i[82];
  assign commit_pkt_o[30] = commit_pkt_o_30_;
  assign commit_pkt_o_29_ = retire_pkt_i[81];
  assign commit_pkt_o[29] = commit_pkt_o_29_;
  assign commit_pkt_o_28_ = retire_pkt_i[80];
  assign commit_pkt_o[28] = commit_pkt_o_28_;
  assign commit_pkt_o_27_ = retire_pkt_i[79];
  assign commit_pkt_o[27] = commit_pkt_o_27_;
  assign commit_pkt_o_26_ = retire_pkt_i[78];
  assign commit_pkt_o[26] = commit_pkt_o_26_;
  assign commit_pkt_o_25_ = retire_pkt_i[77];
  assign commit_pkt_o[25] = commit_pkt_o_25_;
  assign commit_pkt_o_24_ = retire_pkt_i[76];
  assign commit_pkt_o[24] = commit_pkt_o_24_;
  assign commit_pkt_o_23_ = retire_pkt_i[75];
  assign commit_pkt_o[23] = commit_pkt_o_23_;
  assign commit_pkt_o_22_ = retire_pkt_i[74];
  assign commit_pkt_o[22] = commit_pkt_o_22_;
  assign commit_pkt_o_21_ = retire_pkt_i[73];
  assign commit_pkt_o[21] = commit_pkt_o_21_;
  assign commit_pkt_o_15_ = retire_pkt_i[21];
  assign commit_pkt_o[15] = commit_pkt_o_15_;
  assign commit_pkt_o_13_ = retire_pkt_i[9];
  assign commit_pkt_o[13] = commit_pkt_o_13_;
  assign commit_pkt_o_12_ = retire_pkt_i[8];
  assign commit_pkt_o[12] = commit_pkt_o_12_;
  assign commit_pkt_o_11_ = retire_pkt_i[2];
  assign commit_pkt_o[11] = commit_pkt_o_11_;
  assign commit_pkt_o_10_ = retire_pkt_i[3];
  assign commit_pkt_o[10] = commit_pkt_o_10_;
  assign commit_pkt_o_9_ = retire_pkt_i[20];
  assign commit_pkt_o[9] = commit_pkt_o_9_;
  assign commit_pkt_o_8_ = retire_pkt_i[19];
  assign commit_pkt_o[8] = commit_pkt_o_8_;
  assign commit_pkt_o_7_ = retire_pkt_i[16];
  assign commit_pkt_o[7] = commit_pkt_o_7_;
  assign commit_pkt_o_6_ = retire_pkt_i[17];
  assign commit_pkt_o[6] = commit_pkt_o_6_;
  assign commit_pkt_o_5_ = retire_pkt_i[10];
  assign commit_pkt_o[5] = commit_pkt_o_5_;
  assign commit_pkt_o_4_ = retire_pkt_i[18];
  assign commit_pkt_o[4] = commit_pkt_o_4_;
  assign commit_pkt_o_3_ = retire_pkt_i[15];
  assign commit_pkt_o[3] = commit_pkt_o_3_;
  assign commit_pkt_o_2_ = retire_pkt_i[14];
  assign commit_pkt_o[2] = commit_pkt_o_2_;
  assign commit_pkt_o_1_ = retire_pkt_i[1];
  assign commit_pkt_o[1] = commit_pkt_o_1_;
  assign commit_pkt_o_0_ = retire_pkt_i[0];
  assign commit_pkt_o[0] = commit_pkt_o_0_;
  assign decode_info_o[3] = decode_info_o_5_;
  assign decode_info_o[4] = decode_info_o_5_;
  assign decode_info_o[5] = decode_info_o_5_;

  bsg_dff_reset_width_p12
  dcsr_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(dcsr_n),
    .data_o({ decode_info_o_5_, dcsr_r_ebreaks_, dcsr_r_ebreaku_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_prv__1_, dcsr_r_prv__0_, dcsr_r_mprven_, dcsr_r_step_ })
  );


  bsg_dff_reset_width_p40
  dpc_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(dpc_n),
    .data_o(dpc_r)
  );


  bsg_dff_reset_width_p64
  dscratch0_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(dscratch0_n),
    .data_o(dscratch0_r)
  );


  bsg_dff_reset_width_p64
  dscratch1_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(dscratch1_n),
    .data_o(dscratch1_r)
  );


  bsg_dff_reset_width_p15
  mstatus_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(mstatus_n),
    .data_o({ decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ })
  );


  bsg_dff_reset_width_p13
  medeleg_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(medeleg_n),
    .data_o(medeleg_r)
  );


  bsg_dff_reset_width_p3
  mideleg_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ mideleg_n_sei_, mideleg_n_sti_, mideleg_n_ssi_ }),
    .data_o({ mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ })
  );


  bsg_dff_reset_width_p6
  mie_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ mie_n_meie_, mie_n_seie_, mie_n_mtie_, mie_n_stie_, mie_n_msie_, mie_n_ssie_ }),
    .data_o({ mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ })
  );


  bsg_dff_reset_width_p38
  mtvec_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(mtvec_n),
    .data_o(mtvec_r)
  );


  bsg_dff_reset_width_p2
  mcounteren_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ mcounteren_n_ir_, mcounteren_n_cy_ }),
    .data_o({ mcounteren_r_ir_, mcounteren_r_cy_ })
  );


  bsg_dff_reset_width_p64
  mscratch_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(mscratch_n),
    .data_o(mscratch_r)
  );


  bsg_dff_reset_width_p40
  mepc_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(mepc_n),
    .data_o(mepc_r)
  );


  bsg_dff_reset_width_p5
  mcause_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(mcause_n),
    .data_o(mcause_r)
  );


  bsg_dff_reset_width_p40
  mtval_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(mtval_n),
    .data_o(mtval_r)
  );


  bsg_dff_reset_width_p6
  mip_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ m_external_irq_i, mip_n_seip_, timer_irq_i, mip_n_stip_, software_irq_i, mip_n_ssip_ }),
    .data_o({ mip_r_meip_, mip_r_seip_, mip_r_mtip_, mip_r_stip_, mip_r_msip_, mip_r_ssip_ })
  );


  bsg_dff_reset_width_p48
  mcycle_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(mcycle_n),
    .data_o(mcycle_r)
  );


  bsg_dff_reset_width_p48
  minstret_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(minstret_n),
    .data_o(minstret_r)
  );


  bsg_dff_reset_width_p2
  mcountinhibit_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ mcountinhibit_n_ir_, mcountinhibit_n_cy_ }),
    .data_o({ mcountinhibit_r_ir_, mcountinhibit_r_cy_ })
  );


  bsg_dff_reset_width_p38
  stvec_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(stvec_n),
    .data_o(stvec_r)
  );


  bsg_dff_reset_width_p2
  scounteren_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ scounteren_n_ir_, scounteren_n_cy_ }),
    .data_o({ scounteren_r_ir_, scounteren_r_cy_ })
  );


  bsg_dff_reset_width_p64
  sscratch_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(sscratch_n),
    .data_o(sscratch_r)
  );


  bsg_dff_reset_width_p40
  sepc_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(sepc_n),
    .data_o(sepc_r)
  );


  bsg_dff_reset_width_p5
  scause_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(scause_n),
    .data_o(scause_r)
  );


  bsg_dff_reset_width_p40
  stval_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(stval_n),
    .data_o(stval_r)
  );


  bsg_dff_reset_width_p29
  satp_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(satp_n),
    .data_o({ satp_r_mode_, trans_info_o[30:3] })
  );


  bsg_dff_reset_width_p8
  fcsr_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(fcsr_n),
    .data_o({ frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ })
  );


  bsg_priority_encode_width_p16_lo_to_hi_p1
  mcause_exception_enc
  (
    .i({ retire_pkt_i[35:35], 1'b0, retire_pkt_i[34:32], 1'b0, retire_pkt_i[31:22] }),
    .addr_o(exception_ecode_li),
    .v_o(exception_ecode_v_li)
  );


  bsg_priority_encode_width_p16_lo_to_hi_p1
  m_interrupt_enc
  (
    .i({ _0_net__15_, _0_net__14_, _0_net__13_, _0_net__12_, _0_net__11_, _0_net__10_, _0_net__9_, _0_net__8_, _0_net__7_, _0_net__6_, _0_net__5_, _0_net__4_, _0_net__3_, _0_net__2_, _0_net__1_, _0_net__0_ }),
    .addr_o(m_interrupt_icode_li),
    .v_o(m_interrupt_icode_v_li)
  );


  bsg_priority_encode_width_p16_lo_to_hi_p1
  s_interrupt_enc
  (
    .i({ _1_net__15_, _1_net__14_, _1_net__13_, _1_net__12_, _1_net__11_, _1_net__10_, _1_net__9_, _1_net__8_, _1_net__7_, _1_net__6_, _1_net__5_, _1_net__4_, _1_net__3_, _1_net__2_, _1_net__1_, _1_net__0_ }),
    .addr_o(s_interrupt_icode_li),
    .v_o(s_interrupt_icode_v_li)
  );

  assign N99 = ~commit_pkt_o_78_;
  assign N100 = ~commit_pkt_o_77_;
  assign N101 = commit_pkt_o_87_ | commit_pkt_o_88_;
  assign N102 = commit_pkt_o_86_ | N101;
  assign N103 = commit_pkt_o_85_ | N102;
  assign N104 = commit_pkt_o_84_ | N103;
  assign N105 = commit_pkt_o_83_ | N104;
  assign N106 = commit_pkt_o_82_ | N105;
  assign N107 = commit_pkt_o_81_ | N106;
  assign N108 = commit_pkt_o_80_ | N107;
  assign N109 = commit_pkt_o_79_ | N108;
  assign N110 = N99 | N109;
  assign N111 = N100 | N110;
  assign N112 = ~N111;
  assign N113 = commit_pkt_o_87_ | commit_pkt_o_88_;
  assign N114 = commit_pkt_o_86_ | N113;
  assign N115 = commit_pkt_o_85_ | N114;
  assign N116 = commit_pkt_o_84_ | N115;
  assign N117 = commit_pkt_o_83_ | N116;
  assign N118 = commit_pkt_o_82_ | N117;
  assign N119 = commit_pkt_o_81_ | N118;
  assign N120 = commit_pkt_o_80_ | N119;
  assign N121 = commit_pkt_o_79_ | N120;
  assign N122 = commit_pkt_o_78_ | N121;
  assign N123 = N100 | N122;
  assign N124 = ~N123;
  assign N125 = N112 | N124;
  assign N126 = commit_pkt_o_87_ | commit_pkt_o_88_;
  assign N127 = commit_pkt_o_86_ | N126;
  assign N128 = commit_pkt_o_85_ | N127;
  assign N129 = commit_pkt_o_84_ | N128;
  assign N130 = commit_pkt_o_83_ | N129;
  assign N131 = commit_pkt_o_82_ | N130;
  assign N132 = commit_pkt_o_81_ | N131;
  assign N133 = commit_pkt_o_80_ | N132;
  assign N134 = commit_pkt_o_79_ | N133;
  assign N135 = N99 | N134;
  assign N136 = commit_pkt_o_77_ | N135;
  assign N137 = ~N136;
  assign csr_fany_li = N125 | N137;
  assign N138 = ~commit_pkt_o_59_;
  assign N139 = ~commit_pkt_o_58_;
  assign N140 = ~commit_pkt_o_57_;
  assign N141 = commit_pkt_o_62_ | commit_pkt_o_63_;
  assign N142 = commit_pkt_o_61_ | N141;
  assign N143 = commit_pkt_o_60_ | N142;
  assign N144 = N138 | N143;
  assign N145 = N139 | N144;
  assign N146 = N140 | N145;
  assign N147 = ~N146;
  assign N148 = ~commit_pkt_o_63_;
  assign N149 = commit_pkt_o_62_ | N148;
  assign N150 = commit_pkt_o_61_ | N149;
  assign N151 = commit_pkt_o_60_ | N150;
  assign N152 = commit_pkt_o_59_ | N151;
  assign N153 = N139 | N152;
  assign N154 = N140 | N153;
  assign N155 = ~N154;
  assign N156 = N147 | N155;
  assign N157 = commit_pkt_o_62_ | N148;
  assign N158 = commit_pkt_o_61_ | N157;
  assign N159 = commit_pkt_o_60_ | N158;
  assign N160 = N138 | N159;
  assign N161 = N139 | N160;
  assign N162 = N140 | N161;
  assign N163 = ~N162;
  assign N164 = N156 | N163;
  assign N165 = ~commit_pkt_o_60_;
  assign N166 = commit_pkt_o_62_ | N148;
  assign N167 = commit_pkt_o_61_ | N166;
  assign N168 = N165 | N167;
  assign N169 = commit_pkt_o_59_ | N168;
  assign N170 = N139 | N169;
  assign N171 = N140 | N170;
  assign N172 = ~N171;
  assign N173 = N164 | N172;
  assign N174 = ~commit_pkt_o_61_;
  assign N175 = commit_pkt_o_62_ | N148;
  assign N176 = N174 | N175;
  assign N177 = commit_pkt_o_60_ | N176;
  assign N178 = commit_pkt_o_59_ | N177;
  assign N179 = N139 | N178;
  assign N180 = N140 | N179;
  assign N181 = ~N180;
  assign instr_fany_li = N173 | N181;

  bsg_dff_reset_set_clear_width_p1
  debug_mode_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .set_i(enter_debug),
    .clear_i(exit_debug),
    .data_o(decode_info_o[9])
  );


  bsg_dff_reset_00000027
  apc_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(commit_pkt_o[166:128]),
    .data_o(commit_pkt_o[205:167])
  );


  bsg_dff_00000027
  cfg_npc_reg
  (
    .clk_i(clk_i),
    .data_i(cfg_bus_i[59:21]),
    .data_o(cfg_npc_r)
  );

  assign N201 = commit_pkt_o[20:19] < { 1'b1, 1'b1 };

  bsg_dff_reset_3_3
  priv_mode_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ commit_pkt_o[18:18], commit_pkt_o[20:19] }),
    .data_o({ translation_en_r, trans_info_o[32:31] })
  );

  assign N203 = N208 | N318;
  assign N205 = N208 | N321;
  assign N207 = N306 | N213;
  assign N208 = N207 | N302;
  assign N209 = N208 | N339;
  assign N211 = N215 | N314;
  assign N213 = csr_r_addr_i[9] | csr_r_addr_i[8];
  assign N214 = N254 | N213;
  assign N215 = N214 | N302;
  assign N216 = N215 | N321;
  assign N218 = N228 | N314;
  assign N220 = N228 | N321;
  assign N222 = N228 | N339;
  assign N224 = N228 | N281;
  assign N226 = N228 | N271;
  assign N228 = N243 | N302;
  assign N229 = N228 | N275;
  assign N231 = N239 | N314;
  assign N233 = N239 | N318;
  assign N235 = N239 | N321;
  assign N237 = N239 | N339;
  assign N239 = N243 | N292;
  assign N240 = N239 | N281;
  assign N242 = csr_r_addr_i[9] | N326;
  assign N243 = N306 | N242;
  assign N244 = N334 | N300;
  assign N245 = N243 | N244;
  assign N246 = N245 | N314;
  assign N248 = N258 | N318;
  assign N250 = N258 | N321;
  assign N252 = N258 | N339;
  assign N254 = N298 | N324;
  assign N255 = csr_r_addr_i[5] | N329;
  assign N256 = N254 | N333;
  assign N257 = N307 | N255;
  assign N258 = N256 | N257;
  assign N259 = N258 | N281;
  assign N261 = N276 | N314;
  assign N263 = N276 | N318;
  assign N265 = N276 | N321;
  assign N267 = N276 | N339;
  assign N269 = N276 | N281;
  assign N271 = N280 | N331;
  assign N272 = N276 | N271;
  assign N274 = N279 | N330;
  assign N275 = N274 | csr_r_addr_i[0];
  assign N276 = N309 | N302;
  assign N277 = N276 | N275;
  assign N280 = N279 | csr_r_addr_i[1];
  assign N281 = N280 | csr_r_addr_i[0];
  assign N282 = N293 | N281;
  assign N284 = N293 | N314;
  assign N286 = N293 | N318;
  assign N288 = N293 | N321;
  assign N291 = csr_r_addr_i[7] | N290;
  assign N292 = N291 | N300;
  assign N293 = N309 | N292;
  assign N294 = N293 | N339;
  assign N296 = N303 | N314;
  assign N299 = N298 | csr_r_addr_i[10];
  assign N300 = csr_r_addr_i[5] | csr_r_addr_i[4];
  assign N301 = N299 | N333;
  assign N302 = N307 | N300;
  assign N303 = N301 | N302;
  assign N304 = N303 | N321;
  assign N306 = csr_r_addr_i[11] | csr_r_addr_i[10];
  assign N307 = csr_r_addr_i[7] | csr_r_addr_i[6];
  assign N308 = N328 | csr_r_addr_i[4];
  assign N309 = N306 | N333;
  assign N310 = N307 | N308;
  assign N311 = N309 | N310;
  assign N312 = N311 | N314;
  assign N314 = N317 | csr_r_addr_i[0];
  assign N315 = N340 | N314;
  assign N317 = csr_r_addr_i[2] | csr_r_addr_i[1];
  assign N318 = N317 | N331;
  assign N319 = N340 | N318;
  assign N321 = N336 | csr_r_addr_i[0];
  assign N322 = N340 | N321;
  assign N332 = csr_r_addr_i[11] | N324;
  assign N333 = N325 | N326;
  assign N334 = N327 | csr_r_addr_i[6];
  assign N335 = N328 | N329;
  assign N336 = csr_r_addr_i[2] | N330;
  assign N337 = N332 | N333;
  assign N338 = N334 | N335;
  assign N339 = N336 | N331;
  assign N340 = N337 | N338;
  assign N341 = N340 | N339;
  assign N449 = N448 | commit_pkt_o_88_;
  assign N450 = commit_pkt_o_87_ | commit_pkt_o_86_;
  assign N451 = commit_pkt_o_85_ | commit_pkt_o_84_;
  assign N452 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N453 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N454 = commit_pkt_o_79_ | commit_pkt_o_78_;
  assign N455 = N449 | N450;
  assign N456 = N451 | N452;
  assign N457 = N453 | N454;
  assign N458 = N455 | N456;
  assign N459 = N457 | N100;
  assign N460 = N458 | N459;
  assign N462 = N448 | commit_pkt_o_88_;
  assign N463 = commit_pkt_o_87_ | commit_pkt_o_86_;
  assign N464 = commit_pkt_o_85_ | commit_pkt_o_84_;
  assign N465 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N466 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N467 = commit_pkt_o_79_ | N99;
  assign N468 = N462 | N463;
  assign N469 = N464 | N465;
  assign N470 = N466 | N467;
  assign N471 = N468 | N469;
  assign N472 = N470 | commit_pkt_o_77_;
  assign N473 = N471 | N472;
  assign N475 = N448 | commit_pkt_o_88_;
  assign N476 = commit_pkt_o_87_ | commit_pkt_o_86_;
  assign N477 = commit_pkt_o_85_ | commit_pkt_o_84_;
  assign N478 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N479 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N480 = commit_pkt_o_79_ | N99;
  assign N481 = N475 | N476;
  assign N482 = N477 | N478;
  assign N483 = N479 | N480;
  assign N484 = N481 | N482;
  assign N485 = N483 | N100;
  assign N486 = N484 | N485;
  assign N488 = N448 | N1834;
  assign N489 = N1835 | commit_pkt_o_86_;
  assign N490 = commit_pkt_o_85_ | commit_pkt_o_84_;
  assign N491 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N492 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N493 = commit_pkt_o_79_ | N99;
  assign N494 = N488 | N489;
  assign N495 = N490 | N491;
  assign N496 = N492 | N493;
  assign N497 = N494 | N495;
  assign N498 = N496 | commit_pkt_o_77_;
  assign N499 = N497 | N498;
  assign N501 = N448 | commit_pkt_o_88_;
  assign N502 = commit_pkt_o_87_ | commit_pkt_o_86_;
  assign N503 = N1849 | commit_pkt_o_84_;
  assign N504 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N505 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N506 = commit_pkt_o_79_ | commit_pkt_o_78_;
  assign N507 = N501 | N502;
  assign N508 = N503 | N504;
  assign N509 = N505 | N506;
  assign N510 = N507 | N508;
  assign N511 = N509 | commit_pkt_o_77_;
  assign N512 = N510 | N511;
  assign N514 = N448 | commit_pkt_o_88_;
  assign N515 = commit_pkt_o_87_ | commit_pkt_o_86_;
  assign N516 = N1849 | commit_pkt_o_84_;
  assign N517 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N518 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N519 = commit_pkt_o_79_ | N99;
  assign N520 = N514 | N515;
  assign N521 = N516 | N517;
  assign N522 = N518 | N519;
  assign N523 = N520 | N521;
  assign N524 = N522 | commit_pkt_o_77_;
  assign N525 = N523 | N524;
  assign N527 = N448 | commit_pkt_o_88_;
  assign N528 = commit_pkt_o_87_ | commit_pkt_o_86_;
  assign N529 = N1849 | commit_pkt_o_84_;
  assign N530 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N531 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N532 = commit_pkt_o_79_ | N99;
  assign N533 = N527 | N528;
  assign N534 = N529 | N530;
  assign N535 = N531 | N532;
  assign N536 = N533 | N534;
  assign N537 = N535 | N100;
  assign N538 = N536 | N537;
  assign N541 = N448 | commit_pkt_o_88_;
  assign N542 = commit_pkt_o_87_ | commit_pkt_o_86_;
  assign N543 = N1849 | commit_pkt_o_84_;
  assign N544 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N545 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N546 = N540 | commit_pkt_o_78_;
  assign N547 = N541 | N542;
  assign N548 = N543 | N544;
  assign N549 = N545 | N546;
  assign N550 = N547 | N548;
  assign N551 = N549 | commit_pkt_o_77_;
  assign N552 = N550 | N551;
  assign N554 = N448 | commit_pkt_o_88_;
  assign N555 = commit_pkt_o_87_ | commit_pkt_o_86_;
  assign N556 = N1849 | commit_pkt_o_84_;
  assign N557 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N558 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N559 = N540 | commit_pkt_o_78_;
  assign N560 = N554 | N555;
  assign N561 = N556 | N557;
  assign N562 = N558 | N559;
  assign N563 = N560 | N561;
  assign N564 = N562 | N100;
  assign N565 = N563 | N564;
  assign N567 = N448 | commit_pkt_o_88_;
  assign N568 = commit_pkt_o_87_ | commit_pkt_o_86_;
  assign N569 = N1849 | commit_pkt_o_84_;
  assign N570 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N571 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N572 = N540 | N99;
  assign N573 = N567 | N568;
  assign N574 = N569 | N570;
  assign N575 = N571 | N572;
  assign N576 = N573 | N574;
  assign N577 = N575 | commit_pkt_o_77_;
  assign N578 = N576 | N577;
  assign N581 = N448 | commit_pkt_o_88_;
  assign N582 = commit_pkt_o_87_ | commit_pkt_o_86_;
  assign N583 = N1849 | commit_pkt_o_84_;
  assign N584 = N580 | commit_pkt_o_82_;
  assign N585 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N586 = commit_pkt_o_79_ | commit_pkt_o_78_;
  assign N587 = N581 | N582;
  assign N588 = N583 | N584;
  assign N589 = N585 | N586;
  assign N590 = N587 | N588;
  assign N591 = N589 | commit_pkt_o_77_;
  assign N592 = N590 | N591;
  assign N594 = N448 | commit_pkt_o_88_;
  assign N595 = commit_pkt_o_87_ | commit_pkt_o_86_;
  assign N596 = N1849 | commit_pkt_o_84_;
  assign N597 = N580 | commit_pkt_o_82_;
  assign N598 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N599 = commit_pkt_o_79_ | commit_pkt_o_78_;
  assign N600 = N594 | N595;
  assign N601 = N596 | N597;
  assign N602 = N598 | N599;
  assign N603 = N600 | N601;
  assign N604 = N602 | N100;
  assign N605 = N603 | N604;
  assign N607 = N448 | commit_pkt_o_88_;
  assign N608 = commit_pkt_o_87_ | commit_pkt_o_86_;
  assign N609 = N1849 | commit_pkt_o_84_;
  assign N610 = N580 | commit_pkt_o_82_;
  assign N611 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N612 = commit_pkt_o_79_ | N99;
  assign N613 = N607 | N608;
  assign N614 = N609 | N610;
  assign N615 = N611 | N612;
  assign N616 = N613 | N614;
  assign N617 = N615 | commit_pkt_o_77_;
  assign N618 = N616 | N617;
  assign N620 = N448 | commit_pkt_o_88_;
  assign N621 = commit_pkt_o_87_ | commit_pkt_o_86_;
  assign N622 = N1849 | commit_pkt_o_84_;
  assign N623 = N580 | commit_pkt_o_82_;
  assign N624 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N625 = commit_pkt_o_79_ | N99;
  assign N626 = N620 | N621;
  assign N627 = N622 | N623;
  assign N628 = N624 | N625;
  assign N629 = N626 | N627;
  assign N630 = N628 | N100;
  assign N631 = N629 | N630;
  assign N633 = N448 | commit_pkt_o_88_;
  assign N634 = commit_pkt_o_87_ | commit_pkt_o_86_;
  assign N635 = N1849 | commit_pkt_o_84_;
  assign N636 = N580 | commit_pkt_o_82_;
  assign N637 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N638 = N540 | commit_pkt_o_78_;
  assign N639 = N633 | N634;
  assign N640 = N635 | N636;
  assign N641 = N637 | N638;
  assign N642 = N639 | N640;
  assign N643 = N641 | commit_pkt_o_77_;
  assign N644 = N642 | N643;
  assign N647 = N448 | commit_pkt_o_88_;
  assign N648 = commit_pkt_o_87_ | commit_pkt_o_86_;
  assign N649 = N1849 | N646;
  assign N650 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N651 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N652 = commit_pkt_o_79_ | commit_pkt_o_78_;
  assign N653 = N647 | N648;
  assign N654 = N649 | N650;
  assign N655 = N651 | N652;
  assign N656 = N653 | N654;
  assign N657 = N655 | commit_pkt_o_77_;
  assign N658 = N656 | N657;
  assign N660 = N448 | commit_pkt_o_88_;
  assign N661 = commit_pkt_o_87_ | N1848;
  assign N662 = N1849 | commit_pkt_o_84_;
  assign N663 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N664 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N665 = commit_pkt_o_79_ | commit_pkt_o_78_;
  assign N666 = N660 | N661;
  assign N667 = N662 | N663;
  assign N668 = N664 | N665;
  assign N669 = N666 | N667;
  assign N670 = N668 | commit_pkt_o_77_;
  assign N671 = N669 | N670;
  assign N673 = N448 | commit_pkt_o_88_;
  assign N674 = commit_pkt_o_87_ | N1848;
  assign N675 = N1849 | commit_pkt_o_84_;
  assign N676 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N677 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N678 = commit_pkt_o_79_ | commit_pkt_o_78_;
  assign N679 = N673 | N674;
  assign N680 = N675 | N676;
  assign N681 = N677 | N678;
  assign N682 = N679 | N680;
  assign N683 = N681 | N100;
  assign N684 = N682 | N683;
  assign N686 = N448 | commit_pkt_o_88_;
  assign N687 = commit_pkt_o_87_ | N1848;
  assign N688 = N1849 | commit_pkt_o_84_;
  assign N689 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N690 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N691 = commit_pkt_o_79_ | N99;
  assign N692 = N686 | N687;
  assign N693 = N688 | N689;
  assign N694 = N690 | N691;
  assign N695 = N692 | N693;
  assign N696 = N694 | commit_pkt_o_77_;
  assign N697 = N695 | N696;
  assign N699 = N448 | commit_pkt_o_88_;
  assign N700 = commit_pkt_o_87_ | N1848;
  assign N701 = N1849 | commit_pkt_o_84_;
  assign N702 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N703 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N704 = commit_pkt_o_79_ | N99;
  assign N705 = N699 | N700;
  assign N706 = N701 | N702;
  assign N707 = N703 | N704;
  assign N708 = N705 | N706;
  assign N709 = N707 | N100;
  assign N710 = N708 | N709;
  assign N712 = N448 | commit_pkt_o_88_;
  assign N713 = commit_pkt_o_87_ | N1848;
  assign N714 = N1849 | commit_pkt_o_84_;
  assign N715 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N716 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N717 = N540 | commit_pkt_o_78_;
  assign N718 = N712 | N713;
  assign N719 = N714 | N715;
  assign N720 = N716 | N717;
  assign N721 = N718 | N719;
  assign N722 = N720 | commit_pkt_o_77_;
  assign N723 = N721 | N722;
  assign N725 = N448 | commit_pkt_o_88_;
  assign N726 = commit_pkt_o_87_ | N1848;
  assign N727 = N1849 | commit_pkt_o_84_;
  assign N728 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N729 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N730 = N540 | commit_pkt_o_78_;
  assign N731 = N725 | N726;
  assign N732 = N727 | N728;
  assign N733 = N729 | N730;
  assign N734 = N731 | N732;
  assign N735 = N733 | N100;
  assign N736 = N734 | N735;
  assign N738 = N448 | commit_pkt_o_88_;
  assign N739 = commit_pkt_o_87_ | N1848;
  assign N740 = N1849 | commit_pkt_o_84_;
  assign N741 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N742 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N743 = N540 | N99;
  assign N744 = N738 | N739;
  assign N745 = N740 | N741;
  assign N746 = N742 | N743;
  assign N747 = N744 | N745;
  assign N748 = N746 | commit_pkt_o_77_;
  assign N749 = N747 | N748;
  assign N751 = N448 | commit_pkt_o_88_;
  assign N752 = commit_pkt_o_87_ | N1848;
  assign N753 = N1849 | commit_pkt_o_84_;
  assign N754 = N580 | commit_pkt_o_82_;
  assign N755 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N756 = N540 | commit_pkt_o_78_;
  assign N757 = N751 | N752;
  assign N758 = N753 | N754;
  assign N759 = N755 | N756;
  assign N760 = N757 | N758;
  assign N761 = N759 | commit_pkt_o_77_;
  assign N762 = N760 | N761;
  assign N764 = N448 | commit_pkt_o_88_;
  assign N765 = commit_pkt_o_87_ | N1848;
  assign N766 = N1849 | commit_pkt_o_84_;
  assign N767 = N580 | commit_pkt_o_82_;
  assign N768 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N769 = commit_pkt_o_79_ | commit_pkt_o_78_;
  assign N770 = N764 | N765;
  assign N771 = N766 | N767;
  assign N772 = N768 | N769;
  assign N773 = N770 | N771;
  assign N774 = N772 | commit_pkt_o_77_;
  assign N775 = N773 | N774;
  assign N777 = N448 | commit_pkt_o_88_;
  assign N778 = commit_pkt_o_87_ | N1848;
  assign N779 = N1849 | commit_pkt_o_84_;
  assign N780 = N580 | commit_pkt_o_82_;
  assign N781 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N782 = commit_pkt_o_79_ | commit_pkt_o_78_;
  assign N783 = N777 | N778;
  assign N784 = N779 | N780;
  assign N785 = N781 | N782;
  assign N786 = N783 | N784;
  assign N787 = N785 | N100;
  assign N788 = N786 | N787;
  assign N790 = N448 | commit_pkt_o_88_;
  assign N791 = commit_pkt_o_87_ | N1848;
  assign N792 = N1849 | commit_pkt_o_84_;
  assign N793 = N580 | commit_pkt_o_82_;
  assign N794 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N795 = commit_pkt_o_79_ | N99;
  assign N796 = N790 | N791;
  assign N797 = N792 | N793;
  assign N798 = N794 | N795;
  assign N799 = N796 | N797;
  assign N800 = N798 | commit_pkt_o_77_;
  assign N801 = N799 | N800;
  assign N803 = N448 | commit_pkt_o_88_;
  assign N804 = commit_pkt_o_87_ | N1848;
  assign N805 = N1849 | commit_pkt_o_84_;
  assign N806 = N580 | commit_pkt_o_82_;
  assign N807 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N808 = commit_pkt_o_79_ | N99;
  assign N809 = N803 | N804;
  assign N810 = N805 | N806;
  assign N811 = N807 | N808;
  assign N812 = N809 | N810;
  assign N813 = N811 | N100;
  assign N814 = N812 | N813;
  assign N816 = N448 | N1834;
  assign N817 = commit_pkt_o_87_ | N1848;
  assign N818 = N1849 | commit_pkt_o_84_;
  assign N819 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N820 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N821 = commit_pkt_o_79_ | commit_pkt_o_78_;
  assign N822 = N816 | N817;
  assign N823 = N818 | N819;
  assign N824 = N820 | N821;
  assign N825 = N822 | N823;
  assign N826 = N824 | commit_pkt_o_77_;
  assign N827 = N825 | N826;
  assign N829 = N448 | N1834;
  assign N830 = commit_pkt_o_87_ | N1848;
  assign N831 = N1849 | commit_pkt_o_84_;
  assign N832 = commit_pkt_o_83_ | commit_pkt_o_82_;
  assign N833 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N834 = commit_pkt_o_79_ | N99;
  assign N835 = N829 | N830;
  assign N836 = N831 | N832;
  assign N837 = N833 | N834;
  assign N838 = N835 | N836;
  assign N839 = N837 | commit_pkt_o_77_;
  assign N840 = N838 | N839;
  assign N843 = N448 | commit_pkt_o_88_;
  assign N844 = commit_pkt_o_87_ | N1848;
  assign N845 = N1849 | commit_pkt_o_84_;
  assign N846 = commit_pkt_o_83_ | N842;
  assign N847 = commit_pkt_o_81_ | commit_pkt_o_80_;
  assign N848 = commit_pkt_o_79_ | commit_pkt_o_78_;
  assign N849 = N843 | N844;
  assign N850 = N845 | N846;
  assign N851 = N847 | N848;
  assign N852 = N849 | N850;
  assign N853 = N851 | commit_pkt_o_77_;
  assign N854 = N852 | N853;
  assign N857 = N448 | commit_pkt_o_88_;
  assign N858 = N1835 | N1848;
  assign N859 = N1849 | N646;
  assign N860 = commit_pkt_o_83_ | N842;
  assign N861 = N856 | commit_pkt_o_80_;
  assign N862 = commit_pkt_o_79_ | commit_pkt_o_78_;
  assign N863 = N857 | N858;
  assign N864 = N859 | N860;
  assign N865 = N861 | N862;
  assign N866 = N863 | N864;
  assign N867 = N865 | commit_pkt_o_77_;
  assign N868 = N866 | N867;
  assign N870 = N448 | commit_pkt_o_88_;
  assign N871 = N1835 | N1848;
  assign N872 = N1849 | N646;
  assign N873 = commit_pkt_o_83_ | N842;
  assign N874 = N856 | commit_pkt_o_80_;
  assign N875 = commit_pkt_o_79_ | commit_pkt_o_78_;
  assign N876 = N870 | N871;
  assign N877 = N872 | N873;
  assign N878 = N874 | N875;
  assign N879 = N876 | N877;
  assign N880 = N878 | N100;
  assign N881 = N879 | N880;
  assign N883 = N448 | commit_pkt_o_88_;
  assign N884 = N1835 | N1848;
  assign N885 = N1849 | N646;
  assign N886 = commit_pkt_o_83_ | N842;
  assign N887 = N856 | commit_pkt_o_80_;
  assign N888 = commit_pkt_o_79_ | N99;
  assign N889 = N883 | N884;
  assign N890 = N885 | N886;
  assign N891 = N887 | N888;
  assign N892 = N889 | N890;
  assign N893 = N891 | commit_pkt_o_77_;
  assign N894 = N892 | N893;
  assign N896 = N448 | commit_pkt_o_88_;
  assign N897 = N1835 | N1848;
  assign N898 = N1849 | N646;
  assign N899 = commit_pkt_o_83_ | N842;
  assign N900 = N856 | commit_pkt_o_80_;
  assign N901 = commit_pkt_o_79_ | N99;
  assign N902 = N896 | N897;
  assign N903 = N898 | N899;
  assign N904 = N900 | N901;
  assign N905 = N902 | N903;
  assign N906 = N904 | N100;
  assign N907 = N905 | N906;
  assign N1514 = (N1498)? medeleg_r[0] : 
                 (N1500)? medeleg_r[1] : 
                 (N1502)? medeleg_r[2] : 
                 (N1504)? medeleg_r[3] : 
                 (N1506)? medeleg_r[4] : 
                 (N1508)? medeleg_r[5] : 
                 (N1510)? medeleg_r[6] : 
                 (N1512)? medeleg_r[7] : 
                 (N1499)? medeleg_r[8] : 
                 (N1501)? medeleg_r[9] : 
                 (N1503)? 1'b0 : 
                 (N1505)? 1'b0 : 
                 (N1507)? medeleg_r[10] : 
                 (N1509)? medeleg_r[11] : 
                 (N1511)? 1'b0 : 
                 (N1513)? medeleg_r[12] : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 
                 (N0)? 1'b0 : 1'b0;
  assign N0 = 1'b0;
  assign N1797 = { mstatus_r_mpp__1_, mstatus_r_mpp__0_ } < { 1'b1, 1'b1 };
  assign N1803 = commit_pkt_o_87_ | commit_pkt_o_88_;
  assign N1804 = commit_pkt_o_86_ | N1803;
  assign N1805 = commit_pkt_o_85_ | N1804;
  assign N1806 = commit_pkt_o_84_ | N1805;
  assign N1807 = commit_pkt_o_83_ | N1806;
  assign N1808 = commit_pkt_o_82_ | N1807;
  assign N1809 = commit_pkt_o_81_ | N1808;
  assign N1810 = commit_pkt_o_80_ | N1809;
  assign N1811 = commit_pkt_o_79_ | N1810;
  assign N1812 = commit_pkt_o_78_ | N1811;
  assign N1813 = N100 | N1812;
  assign N1814 = ~N1813;
  assign N1815 = commit_pkt_o_87_ | commit_pkt_o_88_;
  assign N1816 = commit_pkt_o_86_ | N1815;
  assign N1817 = commit_pkt_o_85_ | N1816;
  assign N1818 = commit_pkt_o_84_ | N1817;
  assign N1819 = commit_pkt_o_83_ | N1818;
  assign N1820 = commit_pkt_o_82_ | N1819;
  assign N1821 = commit_pkt_o_81_ | N1820;
  assign N1822 = commit_pkt_o_80_ | N1821;
  assign N1823 = commit_pkt_o_79_ | N1822;
  assign N1824 = N99 | N1823;
  assign N1825 = N100 | N1824;
  assign N1826 = ~N1825;
  assign N1827 = N1814 | N1826;
  assign N1834 = ~commit_pkt_o_88_;
  assign N1835 = ~commit_pkt_o_87_;
  assign N1836 = N1835 | N1834;
  assign N1837 = commit_pkt_o_86_ | N1836;
  assign N1838 = commit_pkt_o_85_ | N1837;
  assign N1839 = commit_pkt_o_84_ | N1838;
  assign N1840 = commit_pkt_o_83_ | N1839;
  assign N1841 = commit_pkt_o_82_ | N1840;
  assign N1842 = commit_pkt_o_81_ | N1841;
  assign N1843 = commit_pkt_o_80_ | N1842;
  assign N1844 = commit_pkt_o_79_ | N1843;
  assign N1845 = commit_pkt_o_78_ | N1844;
  assign N1846 = commit_pkt_o_77_ | N1845;
  assign N1847 = ~N1846;
  assign N1848 = ~commit_pkt_o_86_;
  assign N1849 = ~commit_pkt_o_85_;
  assign N1850 = commit_pkt_o_87_ | N1834;
  assign N1851 = N1848 | N1850;
  assign N1852 = N1849 | N1851;
  assign N1853 = commit_pkt_o_84_ | N1852;
  assign N1854 = commit_pkt_o_83_ | N1853;
  assign N1855 = commit_pkt_o_82_ | N1854;
  assign N1856 = commit_pkt_o_81_ | N1855;
  assign N1857 = commit_pkt_o_80_ | N1856;
  assign N1858 = commit_pkt_o_79_ | N1857;
  assign N1859 = commit_pkt_o_78_ | N1858;
  assign N1860 = commit_pkt_o_77_ | N1859;
  assign N1861 = ~N1860;
  assign N1862 = N1847 | N1861;
  assign N1913 = N1835 | N1834;
  assign N1914 = commit_pkt_o_86_ | N1913;
  assign N1915 = commit_pkt_o_85_ | N1914;
  assign N1916 = commit_pkt_o_84_ | N1915;
  assign N1917 = commit_pkt_o_83_ | N1916;
  assign N1918 = commit_pkt_o_82_ | N1917;
  assign N1919 = commit_pkt_o_81_ | N1918;
  assign N1920 = commit_pkt_o_80_ | N1919;
  assign N1921 = commit_pkt_o_79_ | N1920;
  assign N1922 = N99 | N1921;
  assign N1923 = commit_pkt_o_77_ | N1922;
  assign N1924 = ~N1923;
  assign N1925 = commit_pkt_o_87_ | N1834;
  assign N1926 = N1848 | N1925;
  assign N1927 = N1849 | N1926;
  assign N1928 = commit_pkt_o_84_ | N1927;
  assign N1929 = commit_pkt_o_83_ | N1928;
  assign N1930 = commit_pkt_o_82_ | N1929;
  assign N1931 = commit_pkt_o_81_ | N1930;
  assign N1932 = commit_pkt_o_80_ | N1931;
  assign N1933 = commit_pkt_o_79_ | N1932;
  assign N1934 = N99 | N1933;
  assign N1935 = commit_pkt_o_77_ | N1934;
  assign N1936 = ~N1935;
  assign N1937 = N1924 | N1936;
  assign N2001 = N1834 & N1835;
  assign N2002 = N646 & N842;
  assign N2003 = N856 & N2000;
  assign N2004 = N2001 & N2002;
  assign N2005 = N2004 & N2003;
  assign N2007 = commit_pkt_o_86_ | N1849;
  assign N2008 = N580 | N540;
  assign N2009 = commit_pkt_o_78_ | commit_pkt_o_77_;
  assign N2010 = N2007 | N2008;
  assign N2011 = N2010 | N2009;
  assign N2013 = N1848 | N1849;
  assign N2014 = N580 | N540;
  assign N2015 = commit_pkt_o_78_ | commit_pkt_o_77_;
  assign N2016 = N2013 | N2014;
  assign N2017 = N2016 | N2015;
  assign N2019 = commit_pkt_o_86_ | commit_pkt_o_85_;
  assign N2020 = commit_pkt_o_83_ | commit_pkt_o_79_;
  assign N2021 = commit_pkt_o_78_ | N100;
  assign N2022 = N2019 | N2020;
  assign N2023 = N2022 | N2021;
  assign N2024 = commit_pkt_o_86_ | commit_pkt_o_85_;
  assign N2025 = commit_pkt_o_83_ | commit_pkt_o_79_;
  assign N2026 = N99 | N100;
  assign N2027 = N2024 | N2025;
  assign N2028 = N2027 | N2026;
  assign N2046 = { mstatus_r_mpp__1_, mstatus_r_mpp__0_ } < { 1'b1, 1'b1 };
  assign decode_info_o[2] = mstatus_r_fs__0_ | mstatus_r_fs__1_;
  assign N2048 = ~satp_n[28];
  assign N2049 = satp_li_mode__2_ | N2048;
  assign N2050 = satp_li_mode__1_ | N2049;
  assign N2051 = satp_li_mode__0_ | N2050;
  assign N2052 = ~N2051;
  assign N2053 = mstatus_r_fs__0_ & mstatus_r_fs__1_;
  assign N2054 = ~exception_ecode_li[1];
  assign N2055 = exception_ecode_li[2] | exception_ecode_li[3];
  assign N2056 = N2054 | N2055;
  assign N2057 = exception_ecode_li[0] | N2056;
  assign N2058 = ~N2057;
  assign N2059 = exception_ecode_li[2] | exception_ecode_li[3];
  assign N2060 = N2054 | N2059;
  assign N2061 = exception_ecode_li[0] | N2060;
  assign N2062 = ~N2061;
  assign N2063 = ~commit_pkt_o[19];
  assign N2064 = N2063 | commit_pkt_o[20];
  assign N2065 = ~N2064;
  assign N2066 = ~trans_info_o[31];
  assign N2067 = N2066 | trans_info_o[32];
  assign decode_info_o[11] = ~N2067;
  assign N2069 = trans_info_o[31] | trans_info_o[32];
  assign decode_info_o[12] = ~N2069;
  assign N2071 = trans_info_o[31] & trans_info_o[32];
  assign { N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865 } = mcycle_r + 1'b1;
  assign { N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940 } = minstret_r + commit_pkt_o_211_;
  assign ret_pc = (N1)? { sepc_r[37:0], 1'b0 } : 
                  (N185)? { mepc_r[37:0], 1'b0 } : 
                  (N183)? dpc_r[38:0] : 1'b0;
  assign N1 = retire_pkt_i[4];
  assign tvec_pc = (N2)? { cfg_npc_r[38:4], 1'b1, 1'b0 } : 
                   (N189)? stvec_r[36:0] : 
                   (N187)? mtvec_r[36:0] : 1'b0;
  assign N2 = decode_info_o[9];
  assign core_npc = (N3)? { tvec_pc, 1'b0, 1'b0 } : 
                    (N195)? ret_pc : 
                    (N198)? retire_pkt_i[216:178] : 
                    (N193)? commit_pkt_o[205:167] : 1'b0;
  assign N3 = N190;
  assign commit_pkt_o[166:128] = (N4)? { cfg_npc_r[38:4], 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N200)? core_npc : 1'b0;
  assign N4 = N199;
  assign { N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, frm_dyn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mcycle_r } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, minstret_r } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N10)? sstatus_lo : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N13)? sie_lo : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N14)? { stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r[37:37], stvec_r, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, scounteren_r_ir_, 1'b0, scounteren_r_cy_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N16)? sscratch_r : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N17)? { sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r[39:39], sepc_r, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N18)? { scause_r[4:4], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, scause_r[3:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N19)? { stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r[39:39], stval_r } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N20)? sip_lo : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N21)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N23)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cfg_bus_i[20:20] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N26)? { N2053, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, 1'b0, 1'b0, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, 1'b0, 1'b0, mstatus_r_spp_, mstatus_r_mpie_, 1'b0, mstatus_r_spie_, 1'b0, mstatus_r_mie_, 1'b0, mstatus_r_sie_, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N27)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N28)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, medeleg_r[12:12], 1'b0, medeleg_r[11:10], 1'b0, 1'b0, medeleg_r[9:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N29)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mideleg_r_sei_, 1'b0, 1'b0, 1'b0, mideleg_r_sti_, 1'b0, 1'b0, 1'b0, mideleg_r_ssi_, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N30)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mie_r_meie_, 1'b0, mie_r_seie_, 1'b0, mie_r_mtie_, 1'b0, mie_r_stie_, 1'b0, mie_r_msie_, 1'b0, mie_r_ssie_, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N31)? { mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r[37:37], mtvec_r, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N32)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mcounteren_r_ir_, 1'b0, mcounteren_r_cy_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N33)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mip_r_meip_, 1'b0, mip_r_seip_, 1'b0, mip_r_mtip_, 1'b0, mip_r_stip_, 1'b0, mip_r_msip_, 1'b0, mip_r_ssip_, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N34)? mscratch_r : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N35)? { mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r[39:39], mepc_r, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N36)? { mcause_r[4:4], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mcause_r[3:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N37)? { mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r[39:39], mtval_r } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N38)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mcycle_r } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N39)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, minstret_r } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N40)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mcountinhibit_r_ir_, 1'b0, mcountinhibit_r_cy_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N41)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, decode_info_o_5_, 1'b0, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, 1'b0, 1'b0, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, 1'b0, dcsr_r_mprven_, 1'b0, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N42)? { dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r[39:39], dpc_r } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N43)? dscratch0_r : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N44)? dscratch1_r : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N382)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N5 = N204;
  assign N6 = N206;
  assign N7 = N210;
  assign N8 = N212;
  assign N9 = N217;
  assign N10 = N219;
  assign N11 = N221;
  assign N12 = N223;
  assign N13 = N225;
  assign N14 = N227;
  assign N15 = N230;
  assign N16 = N232;
  assign N17 = N234;
  assign N18 = N236;
  assign N19 = N238;
  assign N20 = N241;
  assign N21 = N247;
  assign N22 = N249;
  assign N23 = N251;
  assign N24 = N253;
  assign N25 = N260;
  assign N26 = N262;
  assign N27 = N264;
  assign N28 = N266;
  assign N29 = N268;
  assign N30 = N270;
  assign N31 = N273;
  assign N32 = N278;
  assign N33 = N283;
  assign N34 = N285;
  assign N35 = N287;
  assign N36 = N289;
  assign N37 = N295;
  assign N38 = N297;
  assign N39 = N305;
  assign N40 = N313;
  assign N41 = N316;
  assign N42 = N320;
  assign N43 = N323;
  assign N44 = N342;
  assign N447 = (N5)? 1'b0 : 
                (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N8)? 1'b0 : 
                (N9)? 1'b0 : 
                (N10)? 1'b0 : 
                (N11)? 1'b0 : 
                (N12)? 1'b0 : 
                (N13)? 1'b0 : 
                (N14)? 1'b0 : 
                (N15)? 1'b0 : 
                (N16)? 1'b0 : 
                (N17)? 1'b0 : 
                (N18)? 1'b0 : 
                (N19)? 1'b0 : 
                (N20)? 1'b0 : 
                (N21)? 1'b0 : 
                (N22)? 1'b0 : 
                (N23)? 1'b0 : 
                (N24)? 1'b0 : 
                (N25)? 1'b0 : 
                (N26)? 1'b0 : 
                (N27)? 1'b0 : 
                (N28)? 1'b0 : 
                (N29)? 1'b0 : 
                (N30)? 1'b0 : 
                (N31)? 1'b0 : 
                (N32)? 1'b0 : 
                (N33)? 1'b0 : 
                (N34)? 1'b0 : 
                (N35)? 1'b0 : 
                (N36)? 1'b0 : 
                (N37)? 1'b0 : 
                (N38)? 1'b0 : 
                (N39)? 1'b0 : 
                (N40)? 1'b0 : 
                (N41)? 1'b0 : 
                (N42)? 1'b0 : 
                (N43)? 1'b0 : 
                (N44)? 1'b0 : 
                (N382)? csr_r_v_i : 1'b0;
  assign { csr_r_data_o[63:10], csr_data_lo_9, csr_r_data_o[8:5], csr_data_lo } = (N45)? { N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383 } : 
                                                                                  (N46)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N45 = N202;
  assign N46 = csr_r_addr_i[3];
  assign csr_r_illegal_o = (N45)? N447 : 
                           (N46)? csr_r_v_i : 1'b0;
  assign { fcsr_n[7:5], N972, N971, N970, N969, N968 } = (N47)? { frm_dyn_o, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_ } : 
                                                         (N48)? { commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N49)? { commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_26_, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_ } : 
                                                         (N50)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N51)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N52)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N53)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N54)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N55)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N56)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N57)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N58)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N59)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N60)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N61)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N62)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N63)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N64)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N65)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N66)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N67)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N68)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N69)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N70)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N71)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N72)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N73)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N74)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N75)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N76)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N77)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N78)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N79)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N80)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N81)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 
                                                         (N943)? { frm_dyn_o, fcsr_r_fflags__4_, fcsr_r_fflags__3_, fcsr_r_fflags__2_, fcsr_r_fflags__1_, fcsr_r_fflags__0_ } : 1'b0;
  assign N47 = N461;
  assign N48 = N474;
  assign N49 = N487;
  assign N50 = N500;
  assign N51 = N513;
  assign N52 = N526;
  assign N53 = N539;
  assign N54 = N553;
  assign N55 = N566;
  assign N56 = N579;
  assign N57 = N593;
  assign N58 = N606;
  assign N59 = N619;
  assign N60 = N632;
  assign N61 = N645;
  assign N62 = N659;
  assign N63 = N672;
  assign N64 = N685;
  assign N65 = N698;
  assign N66 = N711;
  assign N67 = N724;
  assign N68 = N737;
  assign N69 = N750;
  assign N70 = N763;
  assign N71 = N776;
  assign N72 = N789;
  assign N73 = N802;
  assign N74 = N815;
  assign N75 = N828;
  assign N76 = N841;
  assign N77 = N855;
  assign N78 = N869;
  assign N79 = N882;
  assign N80 = N895;
  assign N81 = N908;
  assign { N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973 } = (N47)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N48)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N49)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N50)? { retire_pkt_i[120:109], commit_pkt_o_56_, commit_pkt_o_55_, commit_pkt_o_54_, commit_pkt_o_53_, commit_pkt_o_52_, commit_pkt_o_51_, commit_pkt_o_50_, commit_pkt_o_49_, commit_pkt_o_48_, commit_pkt_o_47_, commit_pkt_o_46_, commit_pkt_o_45_, commit_pkt_o_44_, commit_pkt_o_43_, commit_pkt_o_42_, commit_pkt_o_41_, commit_pkt_o_40_, commit_pkt_o_39_, commit_pkt_o_38_, commit_pkt_o_37_, commit_pkt_o_36_, commit_pkt_o_35_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_32_, commit_pkt_o_31_, commit_pkt_o_30_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_26_, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_ } : 
                                                                                                                                                                                                                                                                                                                                   (N51)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N52)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N53)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N54)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N55)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N56)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N57)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N58)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N59)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N60)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N61)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N62)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N63)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N64)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N65)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N66)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N67)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N68)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N69)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N70)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N71)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N72)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N73)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N74)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N75)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N76)? { retire_pkt_i[120:109], commit_pkt_o_56_, commit_pkt_o_55_, commit_pkt_o_54_, commit_pkt_o_53_, commit_pkt_o_52_, commit_pkt_o_51_, commit_pkt_o_50_, commit_pkt_o_49_, commit_pkt_o_48_, commit_pkt_o_47_, commit_pkt_o_46_, commit_pkt_o_45_, commit_pkt_o_44_, commit_pkt_o_43_, commit_pkt_o_42_, commit_pkt_o_41_, commit_pkt_o_40_, commit_pkt_o_39_, commit_pkt_o_38_, commit_pkt_o_37_, commit_pkt_o_36_, commit_pkt_o_35_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_32_, commit_pkt_o_31_, commit_pkt_o_30_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_26_, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_ } : 
                                                                                                                                                                                                                                                                                                                                   (N77)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N78)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N79)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N80)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N81)? minstret_r : 
                                                                                                                                                                                                                                                                                                                                   (N943)? minstret_r : 1'b0;
  assign { mstatus_n[14:10], N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021 } = (N47)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N48)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N49)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N50)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N51)? { N944, N945, N946, N947, N948, N949, N950, N951, N952, N953, N954, N955, N956, N957, N958 } : 
                                                                                                      (N52)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N53)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N54)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N55)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N56)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N57)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N58)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N59)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N60)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N61)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N62)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N63)? { commit_pkt_o_43_, commit_pkt_o_42_, commit_pkt_o_41_, commit_pkt_o_40_, commit_pkt_o_39_, commit_pkt_o_38_, commit_pkt_o_35_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_32_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_26_, commit_pkt_o_24_, commit_pkt_o_22_ } : 
                                                                                                      (N64)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N65)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N66)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N67)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N68)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N69)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N70)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N71)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N72)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N73)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N74)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N75)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N76)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N77)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N78)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N79)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N80)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N81)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 
                                                                                                      (N943)? { decode_info_o[8:6], trans_info_o[0:0], trans_info_o[1:1], mstatus_r_mprv_, mstatus_r_fs__1_, mstatus_r_fs__0_, mstatus_r_mpp__1_, mstatus_r_mpp__0_, mstatus_r_spp_, mstatus_r_mpie_, mstatus_r_spie_, mstatus_r_mie_, mstatus_r_sie_ } : 1'b0;
  assign { mie_n_meie_, mie_n_seie_, mie_n_mtie_, mie_n_stie_, mie_n_msie_, mie_n_ssie_ } = (N47)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N48)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N49)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N50)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N51)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N52)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N53)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N54)? { N959, N960, N961, N962, N963, N964 } : 
                                                                                            (N55)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N56)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N57)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N58)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N59)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N60)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N61)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N62)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N63)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N64)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N65)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N66)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N67)? { commit_pkt_o_32_, commit_pkt_o_30_, commit_pkt_o_28_, commit_pkt_o_26_, commit_pkt_o_24_, commit_pkt_o_22_ } : 
                                                                                            (N68)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N69)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N70)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N71)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N72)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N73)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N74)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N75)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N76)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N77)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N78)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N79)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N80)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N81)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 
                                                                                            (N943)? { mie_r_meie_, mie_r_seie_, mie_r_mtie_, mie_r_stie_, mie_r_msie_, mie_r_ssie_ } : 1'b0;
  assign stvec_n = (N47)? stvec_r : 
                   (N48)? stvec_r : 
                   (N49)? stvec_r : 
                   (N50)? stvec_r : 
                   (N51)? stvec_r : 
                   (N52)? stvec_r : 
                   (N53)? stvec_r : 
                   (N54)? stvec_r : 
                   (N55)? { retire_pkt_i[112:109], commit_pkt_o_56_, commit_pkt_o_55_, commit_pkt_o_54_, commit_pkt_o_53_, commit_pkt_o_52_, commit_pkt_o_51_, commit_pkt_o_50_, commit_pkt_o_49_, commit_pkt_o_48_, commit_pkt_o_47_, commit_pkt_o_46_, commit_pkt_o_45_, commit_pkt_o_44_, commit_pkt_o_43_, commit_pkt_o_42_, commit_pkt_o_41_, commit_pkt_o_40_, commit_pkt_o_39_, commit_pkt_o_38_, commit_pkt_o_37_, commit_pkt_o_36_, commit_pkt_o_35_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_32_, commit_pkt_o_31_, commit_pkt_o_30_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_26_, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_ } : 
                   (N56)? stvec_r : 
                   (N57)? stvec_r : 
                   (N58)? stvec_r : 
                   (N59)? stvec_r : 
                   (N60)? stvec_r : 
                   (N61)? stvec_r : 
                   (N62)? stvec_r : 
                   (N63)? stvec_r : 
                   (N64)? stvec_r : 
                   (N65)? stvec_r : 
                   (N66)? stvec_r : 
                   (N67)? stvec_r : 
                   (N68)? stvec_r : 
                   (N69)? stvec_r : 
                   (N70)? stvec_r : 
                   (N71)? stvec_r : 
                   (N72)? stvec_r : 
                   (N73)? stvec_r : 
                   (N74)? stvec_r : 
                   (N75)? stvec_r : 
                   (N76)? stvec_r : 
                   (N77)? stvec_r : 
                   (N78)? stvec_r : 
                   (N79)? stvec_r : 
                   (N80)? stvec_r : 
                   (N81)? stvec_r : 
                   (N943)? stvec_r : 1'b0;
  assign { scounteren_n_ir_, scounteren_n_cy_ } = (N47)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N48)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N49)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N50)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N51)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N52)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N53)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N54)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N55)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N56)? { commit_pkt_o_23_, commit_pkt_o_21_ } : 
                                                  (N57)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N58)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N59)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N60)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N61)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N62)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N63)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N64)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N65)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N66)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N67)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N68)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N69)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N70)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N71)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N72)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N73)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N74)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N75)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N76)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N77)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N78)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N79)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N80)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N81)? { scounteren_r_ir_, scounteren_r_cy_ } : 
                                                  (N943)? { scounteren_r_ir_, scounteren_r_cy_ } : 1'b0;
  assign sscratch_n = (N47)? sscratch_r : 
                      (N48)? sscratch_r : 
                      (N49)? sscratch_r : 
                      (N50)? sscratch_r : 
                      (N51)? sscratch_r : 
                      (N52)? sscratch_r : 
                      (N53)? sscratch_r : 
                      (N54)? sscratch_r : 
                      (N55)? sscratch_r : 
                      (N56)? sscratch_r : 
                      (N57)? { retire_pkt_i[136:109], commit_pkt_o_56_, commit_pkt_o_55_, commit_pkt_o_54_, commit_pkt_o_53_, commit_pkt_o_52_, commit_pkt_o_51_, commit_pkt_o_50_, commit_pkt_o_49_, commit_pkt_o_48_, commit_pkt_o_47_, commit_pkt_o_46_, commit_pkt_o_45_, commit_pkt_o_44_, commit_pkt_o_43_, commit_pkt_o_42_, commit_pkt_o_41_, commit_pkt_o_40_, commit_pkt_o_39_, commit_pkt_o_38_, commit_pkt_o_37_, commit_pkt_o_36_, commit_pkt_o_35_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_32_, commit_pkt_o_31_, commit_pkt_o_30_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_26_, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_ } : 
                      (N58)? sscratch_r : 
                      (N59)? sscratch_r : 
                      (N60)? sscratch_r : 
                      (N61)? sscratch_r : 
                      (N62)? sscratch_r : 
                      (N63)? sscratch_r : 
                      (N64)? sscratch_r : 
                      (N65)? sscratch_r : 
                      (N66)? sscratch_r : 
                      (N67)? sscratch_r : 
                      (N68)? sscratch_r : 
                      (N69)? sscratch_r : 
                      (N70)? sscratch_r : 
                      (N71)? sscratch_r : 
                      (N72)? sscratch_r : 
                      (N73)? sscratch_r : 
                      (N74)? sscratch_r : 
                      (N75)? sscratch_r : 
                      (N76)? sscratch_r : 
                      (N77)? sscratch_r : 
                      (N78)? sscratch_r : 
                      (N79)? sscratch_r : 
                      (N80)? sscratch_r : 
                      (N81)? sscratch_r : 
                      (N943)? sscratch_r : 1'b0;
  assign { N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031 } = (N47)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N48)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N49)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N50)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N51)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N52)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N53)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N54)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N55)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N56)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N57)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N58)? { retire_pkt_i[113:109], commit_pkt_o_56_, commit_pkt_o_55_, commit_pkt_o_54_, commit_pkt_o_53_, commit_pkt_o_52_, commit_pkt_o_51_, commit_pkt_o_50_, commit_pkt_o_49_, commit_pkt_o_48_, commit_pkt_o_47_, commit_pkt_o_46_, commit_pkt_o_45_, commit_pkt_o_44_, commit_pkt_o_43_, commit_pkt_o_42_, commit_pkt_o_41_, commit_pkt_o_40_, commit_pkt_o_39_, commit_pkt_o_38_, commit_pkt_o_37_, commit_pkt_o_36_, commit_pkt_o_35_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_32_, commit_pkt_o_31_, commit_pkt_o_30_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_26_, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_ } : 
                                                                                                                                                                                                                                                                                                      (N59)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N60)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N61)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N62)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N63)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N64)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N65)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N66)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N67)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N68)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N69)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N70)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N71)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N72)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N73)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N74)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N75)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N76)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N77)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N78)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N79)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N80)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N81)? sepc_r : 
                                                                                                                                                                                                                                                                                                      (N943)? sepc_r : 1'b0;
  assign { N1075, N1074, N1073, N1072, N1071 } = (N47)? scause_r : 
                                                 (N48)? scause_r : 
                                                 (N49)? scause_r : 
                                                 (N50)? scause_r : 
                                                 (N51)? scause_r : 
                                                 (N52)? scause_r : 
                                                 (N53)? scause_r : 
                                                 (N54)? scause_r : 
                                                 (N55)? scause_r : 
                                                 (N56)? scause_r : 
                                                 (N57)? scause_r : 
                                                 (N58)? scause_r : 
                                                 (N59)? { retire_pkt_i[136:136], commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_ } : 
                                                 (N60)? scause_r : 
                                                 (N61)? scause_r : 
                                                 (N62)? scause_r : 
                                                 (N63)? scause_r : 
                                                 (N64)? scause_r : 
                                                 (N65)? scause_r : 
                                                 (N66)? scause_r : 
                                                 (N67)? scause_r : 
                                                 (N68)? scause_r : 
                                                 (N69)? scause_r : 
                                                 (N70)? scause_r : 
                                                 (N71)? scause_r : 
                                                 (N72)? scause_r : 
                                                 (N73)? scause_r : 
                                                 (N74)? scause_r : 
                                                 (N75)? scause_r : 
                                                 (N76)? scause_r : 
                                                 (N77)? scause_r : 
                                                 (N78)? scause_r : 
                                                 (N79)? scause_r : 
                                                 (N80)? scause_r : 
                                                 (N81)? scause_r : 
                                                 (N943)? scause_r : 1'b0;
  assign { N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076 } = (N47)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N48)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N49)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N50)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N51)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N52)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N53)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N54)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N55)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N56)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N57)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N58)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N59)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N60)? { retire_pkt_i[112:109], commit_pkt_o_56_, commit_pkt_o_55_, commit_pkt_o_54_, commit_pkt_o_53_, commit_pkt_o_52_, commit_pkt_o_51_, commit_pkt_o_50_, commit_pkt_o_49_, commit_pkt_o_48_, commit_pkt_o_47_, commit_pkt_o_46_, commit_pkt_o_45_, commit_pkt_o_44_, commit_pkt_o_43_, commit_pkt_o_42_, commit_pkt_o_41_, commit_pkt_o_40_, commit_pkt_o_39_, commit_pkt_o_38_, commit_pkt_o_37_, commit_pkt_o_36_, commit_pkt_o_35_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_32_, commit_pkt_o_31_, commit_pkt_o_30_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_26_, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_ } : 
                                                                                                                                                                                                                                                                                                      (N61)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N62)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N63)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N64)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N65)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N66)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N67)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N68)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N69)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N70)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N71)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N72)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N73)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N74)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N75)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N76)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N77)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N78)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N79)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N80)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N81)? stval_r : 
                                                                                                                                                                                                                                                                                                      (N943)? stval_r : 1'b0;
  assign { mip_n_seip_, mip_n_stip_, mip_n_ssip_ } = (N47)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N48)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N49)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N50)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N51)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N52)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N53)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N54)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N55)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N56)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N57)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N58)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N59)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N60)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N61)? { N965, N966, N967 } : 
                                                     (N62)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N63)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N64)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N65)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N66)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N67)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N68)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N69)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N70)? { commit_pkt_o_30_, commit_pkt_o_26_, commit_pkt_o_22_ } : 
                                                     (N71)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N72)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N73)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N74)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N75)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N76)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N77)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N78)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N79)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N80)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N81)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 
                                                     (N943)? { mip_r_seip_, mip_r_stip_, mip_r_ssip_ } : 1'b0;
  assign { satp_n[28:28], satp_li_mode__2_, satp_li_mode__1_, satp_li_mode__0_, satp_n[27:0] } = (N47)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N48)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N49)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N50)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N51)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N52)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N53)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N54)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N55)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N56)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N57)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N58)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N59)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N60)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N61)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N62)? { retire_pkt_i[136:133], commit_pkt_o_48_, commit_pkt_o_47_, commit_pkt_o_46_, commit_pkt_o_45_, commit_pkt_o_44_, commit_pkt_o_43_, commit_pkt_o_42_, commit_pkt_o_41_, commit_pkt_o_40_, commit_pkt_o_39_, commit_pkt_o_38_, commit_pkt_o_37_, commit_pkt_o_36_, commit_pkt_o_35_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_32_, commit_pkt_o_31_, commit_pkt_o_30_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_26_, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_ } : 
                                                                                                 (N63)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N64)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N65)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N66)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N67)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N68)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N69)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N70)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N71)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N72)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N73)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N74)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N75)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N76)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N77)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N78)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N79)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N80)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N81)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 
                                                                                                 (N943)? { satp_r_mode_, 1'b0, 1'b0, 1'b0, trans_info_o[30:3] } : 1'b0;
  assign medeleg_n = (N47)? medeleg_r : 
                     (N48)? medeleg_r : 
                     (N49)? medeleg_r : 
                     (N50)? medeleg_r : 
                     (N51)? medeleg_r : 
                     (N52)? medeleg_r : 
                     (N53)? medeleg_r : 
                     (N54)? medeleg_r : 
                     (N55)? medeleg_r : 
                     (N56)? medeleg_r : 
                     (N57)? medeleg_r : 
                     (N58)? medeleg_r : 
                     (N59)? medeleg_r : 
                     (N60)? medeleg_r : 
                     (N61)? medeleg_r : 
                     (N62)? medeleg_r : 
                     (N63)? medeleg_r : 
                     (N64)? medeleg_r : 
                     (N65)? { commit_pkt_o_36_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_30_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_26_, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_ } : 
                     (N66)? medeleg_r : 
                     (N67)? medeleg_r : 
                     (N68)? medeleg_r : 
                     (N69)? medeleg_r : 
                     (N70)? medeleg_r : 
                     (N71)? medeleg_r : 
                     (N72)? medeleg_r : 
                     (N73)? medeleg_r : 
                     (N74)? medeleg_r : 
                     (N75)? medeleg_r : 
                     (N76)? medeleg_r : 
                     (N77)? medeleg_r : 
                     (N78)? medeleg_r : 
                     (N79)? medeleg_r : 
                     (N80)? medeleg_r : 
                     (N81)? medeleg_r : 
                     (N943)? medeleg_r : 1'b0;
  assign { mideleg_n_sei_, mideleg_n_sti_, mideleg_n_ssi_ } = (N47)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N48)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N49)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N50)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N51)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N52)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N53)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N54)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N55)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N56)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N57)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N58)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N59)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N60)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N61)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N62)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N63)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N64)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N65)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N66)? { commit_pkt_o_30_, commit_pkt_o_26_, commit_pkt_o_22_ } : 
                                                              (N67)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N68)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N69)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N70)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N71)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N72)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N73)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N74)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N75)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N76)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N77)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N78)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N79)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N80)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N81)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 
                                                              (N943)? { mideleg_r_sei_, mideleg_r_sti_, mideleg_r_ssi_ } : 1'b0;
  assign mtvec_n = (N47)? mtvec_r : 
                   (N48)? mtvec_r : 
                   (N49)? mtvec_r : 
                   (N50)? mtvec_r : 
                   (N51)? mtvec_r : 
                   (N52)? mtvec_r : 
                   (N53)? mtvec_r : 
                   (N54)? mtvec_r : 
                   (N55)? mtvec_r : 
                   (N56)? mtvec_r : 
                   (N57)? mtvec_r : 
                   (N58)? mtvec_r : 
                   (N59)? mtvec_r : 
                   (N60)? mtvec_r : 
                   (N61)? mtvec_r : 
                   (N62)? mtvec_r : 
                   (N63)? mtvec_r : 
                   (N64)? mtvec_r : 
                   (N65)? mtvec_r : 
                   (N66)? mtvec_r : 
                   (N67)? mtvec_r : 
                   (N68)? { retire_pkt_i[112:109], commit_pkt_o_56_, commit_pkt_o_55_, commit_pkt_o_54_, commit_pkt_o_53_, commit_pkt_o_52_, commit_pkt_o_51_, commit_pkt_o_50_, commit_pkt_o_49_, commit_pkt_o_48_, commit_pkt_o_47_, commit_pkt_o_46_, commit_pkt_o_45_, commit_pkt_o_44_, commit_pkt_o_43_, commit_pkt_o_42_, commit_pkt_o_41_, commit_pkt_o_40_, commit_pkt_o_39_, commit_pkt_o_38_, commit_pkt_o_37_, commit_pkt_o_36_, commit_pkt_o_35_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_32_, commit_pkt_o_31_, commit_pkt_o_30_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_26_, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_ } : 
                   (N69)? mtvec_r : 
                   (N70)? mtvec_r : 
                   (N71)? mtvec_r : 
                   (N72)? mtvec_r : 
                   (N73)? mtvec_r : 
                   (N74)? mtvec_r : 
                   (N75)? mtvec_r : 
                   (N76)? mtvec_r : 
                   (N77)? mtvec_r : 
                   (N78)? mtvec_r : 
                   (N79)? mtvec_r : 
                   (N80)? mtvec_r : 
                   (N81)? mtvec_r : 
                   (N943)? mtvec_r : 1'b0;
  assign { mcounteren_n_ir_, mcounteren_n_cy_ } = (N47)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N48)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N49)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N50)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N51)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N52)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N53)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N54)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N55)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N56)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N57)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N58)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N59)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N60)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N61)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N62)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N63)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N64)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N65)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N66)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N67)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N68)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N69)? { commit_pkt_o_23_, commit_pkt_o_21_ } : 
                                                  (N70)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N71)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N72)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N73)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N74)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N75)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N76)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N77)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N78)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N79)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N80)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N81)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 
                                                  (N943)? { mcounteren_r_ir_, mcounteren_r_cy_ } : 1'b0;
  assign mscratch_n = (N47)? mscratch_r : 
                      (N48)? mscratch_r : 
                      (N49)? mscratch_r : 
                      (N50)? mscratch_r : 
                      (N51)? mscratch_r : 
                      (N52)? mscratch_r : 
                      (N53)? mscratch_r : 
                      (N54)? mscratch_r : 
                      (N55)? mscratch_r : 
                      (N56)? mscratch_r : 
                      (N57)? mscratch_r : 
                      (N58)? mscratch_r : 
                      (N59)? mscratch_r : 
                      (N60)? mscratch_r : 
                      (N61)? mscratch_r : 
                      (N62)? mscratch_r : 
                      (N63)? mscratch_r : 
                      (N64)? mscratch_r : 
                      (N65)? mscratch_r : 
                      (N66)? mscratch_r : 
                      (N67)? mscratch_r : 
                      (N68)? mscratch_r : 
                      (N69)? mscratch_r : 
                      (N70)? mscratch_r : 
                      (N71)? { retire_pkt_i[136:109], commit_pkt_o_56_, commit_pkt_o_55_, commit_pkt_o_54_, commit_pkt_o_53_, commit_pkt_o_52_, commit_pkt_o_51_, commit_pkt_o_50_, commit_pkt_o_49_, commit_pkt_o_48_, commit_pkt_o_47_, commit_pkt_o_46_, commit_pkt_o_45_, commit_pkt_o_44_, commit_pkt_o_43_, commit_pkt_o_42_, commit_pkt_o_41_, commit_pkt_o_40_, commit_pkt_o_39_, commit_pkt_o_38_, commit_pkt_o_37_, commit_pkt_o_36_, commit_pkt_o_35_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_32_, commit_pkt_o_31_, commit_pkt_o_30_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_26_, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_ } : 
                      (N72)? mscratch_r : 
                      (N73)? mscratch_r : 
                      (N74)? mscratch_r : 
                      (N75)? mscratch_r : 
                      (N76)? mscratch_r : 
                      (N77)? mscratch_r : 
                      (N78)? mscratch_r : 
                      (N79)? mscratch_r : 
                      (N80)? mscratch_r : 
                      (N81)? mscratch_r : 
                      (N943)? mscratch_r : 1'b0;
  assign { N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116 } = (N47)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N48)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N49)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N50)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N51)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N52)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N53)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N54)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N55)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N56)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N57)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N58)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N59)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N60)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N61)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N62)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N63)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N64)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N65)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N66)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N67)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N68)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N69)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N70)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N71)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N72)? { retire_pkt_i[113:109], commit_pkt_o_56_, commit_pkt_o_55_, commit_pkt_o_54_, commit_pkt_o_53_, commit_pkt_o_52_, commit_pkt_o_51_, commit_pkt_o_50_, commit_pkt_o_49_, commit_pkt_o_48_, commit_pkt_o_47_, commit_pkt_o_46_, commit_pkt_o_45_, commit_pkt_o_44_, commit_pkt_o_43_, commit_pkt_o_42_, commit_pkt_o_41_, commit_pkt_o_40_, commit_pkt_o_39_, commit_pkt_o_38_, commit_pkt_o_37_, commit_pkt_o_36_, commit_pkt_o_35_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_32_, commit_pkt_o_31_, commit_pkt_o_30_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_26_, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_ } : 
                                                                                                                                                                                                                                                                                                      (N73)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N74)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N75)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N76)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N77)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N78)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N79)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N80)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N81)? mepc_r : 
                                                                                                                                                                                                                                                                                                      (N943)? mepc_r : 1'b0;
  assign { N1160, N1159, N1158, N1157, N1156 } = (N47)? mcause_r : 
                                                 (N48)? mcause_r : 
                                                 (N49)? mcause_r : 
                                                 (N50)? mcause_r : 
                                                 (N51)? mcause_r : 
                                                 (N52)? mcause_r : 
                                                 (N53)? mcause_r : 
                                                 (N54)? mcause_r : 
                                                 (N55)? mcause_r : 
                                                 (N56)? mcause_r : 
                                                 (N57)? mcause_r : 
                                                 (N58)? mcause_r : 
                                                 (N59)? mcause_r : 
                                                 (N60)? mcause_r : 
                                                 (N61)? mcause_r : 
                                                 (N62)? mcause_r : 
                                                 (N63)? mcause_r : 
                                                 (N64)? mcause_r : 
                                                 (N65)? mcause_r : 
                                                 (N66)? mcause_r : 
                                                 (N67)? mcause_r : 
                                                 (N68)? mcause_r : 
                                                 (N69)? mcause_r : 
                                                 (N70)? mcause_r : 
                                                 (N71)? mcause_r : 
                                                 (N72)? mcause_r : 
                                                 (N73)? { retire_pkt_i[136:136], commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_ } : 
                                                 (N74)? mcause_r : 
                                                 (N75)? mcause_r : 
                                                 (N76)? mcause_r : 
                                                 (N77)? mcause_r : 
                                                 (N78)? mcause_r : 
                                                 (N79)? mcause_r : 
                                                 (N80)? mcause_r : 
                                                 (N81)? mcause_r : 
                                                 (N943)? mcause_r : 1'b0;
  assign { N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161 } = (N47)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N48)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N49)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N50)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N51)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N52)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N53)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N54)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N55)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N56)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N57)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N58)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N59)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N60)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N61)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N62)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N63)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N64)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N65)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N66)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N67)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N68)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N69)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N70)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N71)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N72)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N73)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N74)? { retire_pkt_i[112:109], commit_pkt_o_56_, commit_pkt_o_55_, commit_pkt_o_54_, commit_pkt_o_53_, commit_pkt_o_52_, commit_pkt_o_51_, commit_pkt_o_50_, commit_pkt_o_49_, commit_pkt_o_48_, commit_pkt_o_47_, commit_pkt_o_46_, commit_pkt_o_45_, commit_pkt_o_44_, commit_pkt_o_43_, commit_pkt_o_42_, commit_pkt_o_41_, commit_pkt_o_40_, commit_pkt_o_39_, commit_pkt_o_38_, commit_pkt_o_37_, commit_pkt_o_36_, commit_pkt_o_35_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_32_, commit_pkt_o_31_, commit_pkt_o_30_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_26_, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_ } : 
                                                                                                                                                                                                                                                                                                      (N75)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N76)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N77)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N78)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N79)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N80)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N81)? mtval_r : 
                                                                                                                                                                                                                                                                                                      (N943)? mtval_r : 1'b0;
  assign { N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201 } = (N47)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N48)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N49)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N50)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N51)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N52)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N53)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N54)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N55)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N56)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N57)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N58)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N59)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N60)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N61)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N62)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N63)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N64)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N65)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N66)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N67)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N68)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N69)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N70)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N71)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N72)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N73)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N74)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N75)? { retire_pkt_i[120:109], commit_pkt_o_56_, commit_pkt_o_55_, commit_pkt_o_54_, commit_pkt_o_53_, commit_pkt_o_52_, commit_pkt_o_51_, commit_pkt_o_50_, commit_pkt_o_49_, commit_pkt_o_48_, commit_pkt_o_47_, commit_pkt_o_46_, commit_pkt_o_45_, commit_pkt_o_44_, commit_pkt_o_43_, commit_pkt_o_42_, commit_pkt_o_41_, commit_pkt_o_40_, commit_pkt_o_39_, commit_pkt_o_38_, commit_pkt_o_37_, commit_pkt_o_36_, commit_pkt_o_35_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_32_, commit_pkt_o_31_, commit_pkt_o_30_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_26_, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_ } : 
                                                                                                                                                                                                                                                                                                                                                              (N76)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N77)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N78)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N79)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N80)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N81)? mcycle_r : 
                                                                                                                                                                                                                                                                                                                                                              (N943)? mcycle_r : 1'b0;
  assign { mcountinhibit_n_ir_, mcountinhibit_n_cy_ } = (N47)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N48)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N49)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N50)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N51)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N52)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N53)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N54)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N55)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N56)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N57)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N58)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N59)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N60)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N61)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N62)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N63)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N64)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N65)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N66)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N67)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N68)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N69)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N70)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N71)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N72)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N73)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N74)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N75)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N76)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N77)? { commit_pkt_o_23_, commit_pkt_o_21_ } : 
                                                        (N78)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N79)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N80)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N81)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 
                                                        (N943)? { mcountinhibit_r_ir_, mcountinhibit_r_cy_ } : 1'b0;
  assign { dcsr_n[11:8], N1254, N1253, N1252, N1251, dcsr_n[1:0], N1250, N1249 } = (N47)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N48)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N49)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N50)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N51)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N52)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N53)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N54)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N55)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N56)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N57)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N58)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N59)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N60)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N61)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N62)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N63)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N64)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N65)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N66)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N67)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N68)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N69)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N70)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N71)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N72)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N73)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N74)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N75)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N76)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N77)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N78)? { commit_pkt_o_37_, commit_pkt_o_35_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_30_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_25_, commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_ } : 
                                                                                   (N79)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N80)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N81)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                                                                                   (N943)? { decode_info_o_5_, decode_info_o_5_, decode_info_o_5_, dcsr_r_stepie_, dcsr_r_cause__3_, dcsr_r_cause__2_, dcsr_r_cause__1_, dcsr_r_cause__0_, dcsr_r_mprven_, dcsr_r_step_, dcsr_r_prv__1_, dcsr_r_prv__0_ } : 1'b0;
  assign { N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255 } = (N47)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N48)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N49)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N50)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N51)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N52)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N53)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N54)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N55)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N56)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N57)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N58)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N59)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N60)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N61)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N62)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N63)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N64)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N65)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N66)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N67)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N68)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N69)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N70)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N71)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N72)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N73)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N74)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N75)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N76)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N77)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N78)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N79)? { retire_pkt_i[112:109], commit_pkt_o_56_, commit_pkt_o_55_, commit_pkt_o_54_, commit_pkt_o_53_, commit_pkt_o_52_, commit_pkt_o_51_, commit_pkt_o_50_, commit_pkt_o_49_, commit_pkt_o_48_, commit_pkt_o_47_, commit_pkt_o_46_, commit_pkt_o_45_, commit_pkt_o_44_, commit_pkt_o_43_, commit_pkt_o_42_, commit_pkt_o_41_, commit_pkt_o_40_, commit_pkt_o_39_, commit_pkt_o_38_, commit_pkt_o_37_, commit_pkt_o_36_, commit_pkt_o_35_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_32_, commit_pkt_o_31_, commit_pkt_o_30_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_26_, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_ } : 
                                                                                                                                                                                                                                                                                                      (N80)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N81)? dpc_r : 
                                                                                                                                                                                                                                                                                                      (N943)? dpc_r : 1'b0;
  assign dscratch0_n = (N47)? dscratch0_r : 
                       (N48)? dscratch0_r : 
                       (N49)? dscratch0_r : 
                       (N50)? dscratch0_r : 
                       (N51)? dscratch0_r : 
                       (N52)? dscratch0_r : 
                       (N53)? dscratch0_r : 
                       (N54)? dscratch0_r : 
                       (N55)? dscratch0_r : 
                       (N56)? dscratch0_r : 
                       (N57)? dscratch0_r : 
                       (N58)? dscratch0_r : 
                       (N59)? dscratch0_r : 
                       (N60)? dscratch0_r : 
                       (N61)? dscratch0_r : 
                       (N62)? dscratch0_r : 
                       (N63)? dscratch0_r : 
                       (N64)? dscratch0_r : 
                       (N65)? dscratch0_r : 
                       (N66)? dscratch0_r : 
                       (N67)? dscratch0_r : 
                       (N68)? dscratch0_r : 
                       (N69)? dscratch0_r : 
                       (N70)? dscratch0_r : 
                       (N71)? dscratch0_r : 
                       (N72)? dscratch0_r : 
                       (N73)? dscratch0_r : 
                       (N74)? dscratch0_r : 
                       (N75)? dscratch0_r : 
                       (N76)? dscratch0_r : 
                       (N77)? dscratch0_r : 
                       (N78)? dscratch0_r : 
                       (N79)? dscratch0_r : 
                       (N80)? { retire_pkt_i[136:109], commit_pkt_o_56_, commit_pkt_o_55_, commit_pkt_o_54_, commit_pkt_o_53_, commit_pkt_o_52_, commit_pkt_o_51_, commit_pkt_o_50_, commit_pkt_o_49_, commit_pkt_o_48_, commit_pkt_o_47_, commit_pkt_o_46_, commit_pkt_o_45_, commit_pkt_o_44_, commit_pkt_o_43_, commit_pkt_o_42_, commit_pkt_o_41_, commit_pkt_o_40_, commit_pkt_o_39_, commit_pkt_o_38_, commit_pkt_o_37_, commit_pkt_o_36_, commit_pkt_o_35_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_32_, commit_pkt_o_31_, commit_pkt_o_30_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_26_, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_ } : 
                       (N81)? dscratch0_r : 
                       (N943)? dscratch0_r : 1'b0;
  assign dscratch1_n = (N47)? dscratch1_r : 
                       (N48)? dscratch1_r : 
                       (N49)? dscratch1_r : 
                       (N50)? dscratch1_r : 
                       (N51)? dscratch1_r : 
                       (N52)? dscratch1_r : 
                       (N53)? dscratch1_r : 
                       (N54)? dscratch1_r : 
                       (N55)? dscratch1_r : 
                       (N56)? dscratch1_r : 
                       (N57)? dscratch1_r : 
                       (N58)? dscratch1_r : 
                       (N59)? dscratch1_r : 
                       (N60)? dscratch1_r : 
                       (N61)? dscratch1_r : 
                       (N62)? dscratch1_r : 
                       (N63)? dscratch1_r : 
                       (N64)? dscratch1_r : 
                       (N65)? dscratch1_r : 
                       (N66)? dscratch1_r : 
                       (N67)? dscratch1_r : 
                       (N68)? dscratch1_r : 
                       (N69)? dscratch1_r : 
                       (N70)? dscratch1_r : 
                       (N71)? dscratch1_r : 
                       (N72)? dscratch1_r : 
                       (N73)? dscratch1_r : 
                       (N74)? dscratch1_r : 
                       (N75)? dscratch1_r : 
                       (N76)? dscratch1_r : 
                       (N77)? dscratch1_r : 
                       (N78)? dscratch1_r : 
                       (N79)? dscratch1_r : 
                       (N80)? dscratch1_r : 
                       (N81)? { retire_pkt_i[136:109], commit_pkt_o_56_, commit_pkt_o_55_, commit_pkt_o_54_, commit_pkt_o_53_, commit_pkt_o_52_, commit_pkt_o_51_, commit_pkt_o_50_, commit_pkt_o_49_, commit_pkt_o_48_, commit_pkt_o_47_, commit_pkt_o_46_, commit_pkt_o_45_, commit_pkt_o_44_, commit_pkt_o_43_, commit_pkt_o_42_, commit_pkt_o_41_, commit_pkt_o_40_, commit_pkt_o_39_, commit_pkt_o_38_, commit_pkt_o_37_, commit_pkt_o_36_, commit_pkt_o_35_, commit_pkt_o_34_, commit_pkt_o_33_, commit_pkt_o_32_, commit_pkt_o_31_, commit_pkt_o_30_, commit_pkt_o_29_, commit_pkt_o_28_, commit_pkt_o_27_, commit_pkt_o_26_, commit_pkt_o_25_, commit_pkt_o_24_, commit_pkt_o_23_, commit_pkt_o_22_, commit_pkt_o_21_ } : 
                       (N943)? dscratch1_r : 1'b0;
  assign { N1302, N1301 } = (N82)? { 1'b1, 1'b1 } : 
                            (N1991)? { 1'b0, 1'b1 } : 
                            (N1300)? trans_info_o[32:31] : 1'b0;
  assign N82 = N1297;
  assign { N1308, N1306, N1303 } = (N82)? { N1025, N1023, N1021 } : 
                                   (N1991)? { trans_info_o[31:31], mstatus_r_sie_, 1'b0 } : 
                                   (N1300)? { N1025, N1023, N1021 } : 1'b0;
  assign { N1310, N1309, N1307, N1305 } = (N82)? { trans_info_o[32:31], mstatus_r_mie_, 1'b0 } : 
                                          (N1304)? { N1027, N1026, N1024, N1022 } : 
                                          (N0)? { N1027, N1026, N1024, N1022 } : 1'b0;
  assign { N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311 } = (N82)? { commit_pkt_o[205:205], commit_pkt_o[205:205], commit_pkt_o[205:168] } : 
                                                                                                                                                                                                                                                                                                      (N1304)? { N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116 } : 
                                                                                                                                                                                                                                                                                                      (N0)? { N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116 } : 1'b0;
  assign { N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351 } = (N82)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                      (N1304)? { N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161 } : 
                                                                                                                                                                                                                                                                                                      (N0)? { N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161 } : 1'b0;
  assign { N1395, N1394, N1393, N1392, N1391 } = (N82)? { 1'b1, m_interrupt_icode_li } : 
                                                 (N1304)? { N1160, N1159, N1158, N1157, N1156 } : 
                                                 (N0)? { N1160, N1159, N1158, N1157, N1156 } : 1'b0;
  assign N1396 = (N82)? 1'b1 : 
                 (N1991)? 1'b1 : 
                 (N1300)? 1'b0 : 1'b0;
  assign { N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397 } = (N82)? { N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031 } : 
                                                                                                                                                                                                                                                                                                      (N1991)? { commit_pkt_o[205:205], commit_pkt_o[205:205], commit_pkt_o[205:168] } : 
                                                                                                                                                                                                                                                                                                      (N1300)? { N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031 } : 1'b0;
  assign { N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437 } = (N82)? { N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076 } : 
                                                                                                                                                                                                                                                                                                      (N1991)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                      (N1300)? { N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076 } : 1'b0;
  assign { N1481, N1480, N1479, N1478, N1477 } = (N82)? { N1075, N1074, N1073, N1072, N1071 } : 
                                                 (N1991)? { 1'b1, s_interrupt_icode_li } : 
                                                 (N1300)? { N1075, N1074, N1073, N1072, N1071 } : 1'b0;
  assign { N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518 } = (N83)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, commit_pkt_o_88_, commit_pkt_o_87_, commit_pkt_o_86_, commit_pkt_o_85_, commit_pkt_o_84_, commit_pkt_o_83_, commit_pkt_o_82_, commit_pkt_o_81_, commit_pkt_o_80_, commit_pkt_o_79_, commit_pkt_o_78_, commit_pkt_o_77_, commit_pkt_o_76_, commit_pkt_o_75_, commit_pkt_o_74_, commit_pkt_o_73_, commit_pkt_o_72_, commit_pkt_o_71_, commit_pkt_o_70_, commit_pkt_o_69_, commit_pkt_o_68_, commit_pkt_o_67_, commit_pkt_o_66_, commit_pkt_o_65_, commit_pkt_o_64_, commit_pkt_o_63_, commit_pkt_o_62_, commit_pkt_o_61_, commit_pkt_o_60_, commit_pkt_o_59_, commit_pkt_o_58_, commit_pkt_o_57_ } : 
                                                                                                                                                                                                                                                                                                      (N84)? { commit_pkt_o_127_, commit_pkt_o_127_, commit_pkt_o_126_, commit_pkt_o_125_, commit_pkt_o_124_, commit_pkt_o_123_, commit_pkt_o_122_, commit_pkt_o_121_, commit_pkt_o_120_, commit_pkt_o_119_, commit_pkt_o_118_, commit_pkt_o_117_, commit_pkt_o_116_, commit_pkt_o_115_, commit_pkt_o_114_, commit_pkt_o_113_, commit_pkt_o_112_, commit_pkt_o_111_, commit_pkt_o_110_, commit_pkt_o_109_, commit_pkt_o_108_, commit_pkt_o_107_, commit_pkt_o_106_, commit_pkt_o_105_, commit_pkt_o_104_, commit_pkt_o_103_, commit_pkt_o_102_, commit_pkt_o_101_, commit_pkt_o_100_, commit_pkt_o_99_, commit_pkt_o_98_, commit_pkt_o_97_, commit_pkt_o_96_, commit_pkt_o_95_, commit_pkt_o_94_, commit_pkt_o_93_, commit_pkt_o_92_, commit_pkt_o_91_, commit_pkt_o_90_, commit_pkt_o_89_ } : 1'b0;
  assign N83 = N2062;
  assign N84 = N2061;
  assign { N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558 } = (N85)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, commit_pkt_o_88_, commit_pkt_o_87_, commit_pkt_o_86_, commit_pkt_o_85_, commit_pkt_o_84_, commit_pkt_o_83_, commit_pkt_o_82_, commit_pkt_o_81_, commit_pkt_o_80_, commit_pkt_o_79_, commit_pkt_o_78_, commit_pkt_o_77_, commit_pkt_o_76_, commit_pkt_o_75_, commit_pkt_o_74_, commit_pkt_o_73_, commit_pkt_o_72_, commit_pkt_o_71_, commit_pkt_o_70_, commit_pkt_o_69_, commit_pkt_o_68_, commit_pkt_o_67_, commit_pkt_o_66_, commit_pkt_o_65_, commit_pkt_o_64_, commit_pkt_o_63_, commit_pkt_o_62_, commit_pkt_o_61_, commit_pkt_o_60_, commit_pkt_o_59_, commit_pkt_o_58_, commit_pkt_o_57_ } : 
                                                                                                                                                                                                                                                                                                      (N86)? { commit_pkt_o_127_, commit_pkt_o_127_, commit_pkt_o_126_, commit_pkt_o_125_, commit_pkt_o_124_, commit_pkt_o_123_, commit_pkt_o_122_, commit_pkt_o_121_, commit_pkt_o_120_, commit_pkt_o_119_, commit_pkt_o_118_, commit_pkt_o_117_, commit_pkt_o_116_, commit_pkt_o_115_, commit_pkt_o_114_, commit_pkt_o_113_, commit_pkt_o_112_, commit_pkt_o_111_, commit_pkt_o_110_, commit_pkt_o_109_, commit_pkt_o_108_, commit_pkt_o_107_, commit_pkt_o_106_, commit_pkt_o_105_, commit_pkt_o_104_, commit_pkt_o_103_, commit_pkt_o_102_, commit_pkt_o_101_, commit_pkt_o_100_, commit_pkt_o_99_, commit_pkt_o_98_, commit_pkt_o_97_, commit_pkt_o_96_, commit_pkt_o_95_, commit_pkt_o_94_, commit_pkt_o_93_, commit_pkt_o_92_, commit_pkt_o_91_, commit_pkt_o_90_, commit_pkt_o_89_ } : 1'b0;
  assign N85 = N2058;
  assign N86 = N2057;
  assign { N1599, N1598 } = (N2)? trans_info_o[32:31] : 
                            (N1992)? { 1'b0, 1'b1 } : 
                            (N1517)? { 1'b1, 1'b1 } : 1'b0;
  assign { N1606, N1605, N1604, N1603, N1602, N1601, N1600 } = (N2)? { N1027, N1026, N1025, N1024, N1023, N1022, N1021 } : 
                                                               (N1992)? { N1027, N1026, trans_info_o[31:31], N1024, mstatus_r_sie_, N1022, 1'b0 } : 
                                                               (N1517)? { trans_info_o[32:31], N1025, mstatus_r_mie_, N1023, 1'b0, N1021 } : 1'b0;
  assign { N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607 } = (N2)? { N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031 } : 
                                                                                                                                                                                                                                                                                                      (N1992)? { commit_pkt_o[205:205], commit_pkt_o[205:205], commit_pkt_o[205:168] } : 
                                                                                                                                                                                                                                                                                                      (N1517)? { N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031 } : 1'b0;
  assign { N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647 } = (N2)? { N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076 } : 
                                                                                                                                                                                                                                                                                                      (N1992)? { N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518 } : 
                                                                                                                                                                                                                                                                                                      (N1517)? { N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076 } : 1'b0;
  assign { N1691, N1690, N1689, N1688, N1687 } = (N2)? { N1075, N1074, N1073, N1072, N1071 } : 
                                                 (N1992)? { 1'b0, exception_ecode_li } : 
                                                 (N1517)? { N1075, N1074, N1073, N1072, N1071 } : 1'b0;
  assign { N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692 } = (N2)? { N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116 } : 
                                                                                                                                                                                                                                                                                                      (N1992)? { N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116 } : 
                                                                                                                                                                                                                                                                                                      (N1517)? { commit_pkt_o[205:205], commit_pkt_o[205:205], commit_pkt_o[205:168] } : 1'b0;
  assign { N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732 } = (N2)? { N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161 } : 
                                                                                                                                                                                                                                                                                                      (N1992)? { N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161 } : 
                                                                                                                                                                                                                                                                                                      (N1517)? { N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558 } : 1'b0;
  assign { N1776, N1775, N1774, N1773, N1772 } = (N2)? { N1160, N1159, N1158, N1157, N1156 } : 
                                                 (N1992)? { N1160, N1159, N1158, N1157, N1156 } : 
                                                 (N1517)? { 1'b0, exception_ecode_li } : 1'b0;
  assign scause_n = (N87)? { N1481, N1480, N1479, N1478, N1477 } : 
                    (N1990)? { N1691, N1690, N1689, N1688, N1687 } : 
                    (N1296)? { N1075, N1074, N1073, N1072, N1071 } : 1'b0;
  assign N87 = retire_pkt_i[13];
  assign { N1778, N1777 } = (N87)? { N1302, N1301 } : 
                            (N1990)? { N1599, N1598 } : 
                            (N1296)? trans_info_o[32:31] : 1'b0;
  assign { N1785, N1784, N1783, N1782, N1781, N1780, N1779 } = (N87)? { N1310, N1309, N1308, N1307, N1306, N1305, N1303 } : 
                                                               (N1990)? { N1606, N1605, N1604, N1603, N1602, N1601, N1600 } : 
                                                               (N1296)? { N1027, N1026, N1025, N1024, N1023, N1022, N1021 } : 1'b0;
  assign mepc_n = (N87)? { N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311 } : 
                  (N1990)? { N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692 } : 
                  (N1296)? { N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116 } : 1'b0;
  assign mtval_n = (N87)? { N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351 } : 
                   (N1990)? { N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732 } : 
                   (N1296)? { N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161 } : 1'b0;
  assign mcause_n = (N87)? { N1395, N1394, N1393, N1392, N1391 } : 
                    (N1990)? { N1776, N1775, N1774, N1773, N1772 } : 
                    (N1296)? { N1160, N1159, N1158, N1157, N1156 } : 1'b0;
  assign interrupt_v_lo = (N87)? N1396 : 
                          (N1786)? 1'b0 : 
                          (N0)? 1'b0 : 1'b0;
  assign sepc_n = (N87)? { N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397 } : 
                  (N1990)? { N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607 } : 
                  (N1296)? { N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031 } : 1'b0;
  assign stval_n = (N87)? { N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437 } : 
                   (N1990)? { N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647 } : 
                   (N1296)? { N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076 } : 1'b0;
  assign commit_pkt_o[17] = (N87)? 1'b0 : 
                            (N1990)? 1'b1 : 
                            (N1296)? 1'b0 : 1'b0;
  assign enter_debug = (N2)? retire_pkt_i[7] : 
                       (N1993)? 1'b1 : 
                       (N1996)? 1'b1 : 
                       (N1999)? 1'b1 : 
                       (N1792)? 1'b0 : 1'b0;
  assign dpc_n = (N2)? { N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255 } : 
                 (N1993)? { commit_pkt_o[205:205], commit_pkt_o[205:167] } : 
                 (N1996)? { commit_pkt_o[205:205], commit_pkt_o[205:167] } : 
                 (N1999)? { core_npc[38:38], core_npc } : 
                 (N1792)? { N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255 } : 1'b0;
  assign dcsr_n[7:2] = (N2)? { N1254, N1253, N1252, N1251, N1250, N1249 } : 
                       (N1993)? { 1'b0, 1'b0, 1'b1, 1'b1, trans_info_o[32:31] } : 
                       (N1996)? { 1'b0, 1'b0, 1'b0, 1'b1, trans_info_o[32:31] } : 
                       (N1999)? { 1'b0, 1'b1, 1'b0, 1'b0, trans_info_o[32:31] } : 
                       (N1792)? { N1254, N1253, N1252, N1251, N1250, N1249 } : 1'b0;
  assign { N1795, N1794 } = (N88)? { dcsr_r_prv__1_, dcsr_r_prv__0_ } : 
                            (N1793)? { N1778, N1777 } : 1'b0;
  assign N88 = exit_debug;
  assign N1799 = (N89)? 1'b0 : 
                 (N1798)? N1030 : 1'b0;
  assign N89 = N1797;
  assign { N1801, N1800 } = (N90)? { mstatus_r_mpp__1_, mstatus_r_mpp__0_ } : 
                            (N1796)? { N1795, N1794 } : 1'b0;
  assign N90 = retire_pkt_i[5];
  assign { N1802, mstatus_n[6:5], mstatus_n[3:3], mstatus_n[1:1] } = (N90)? { N1799, 1'b0, 1'b0, 1'b1, mstatus_r_mpie_ } : 
                                                                     (N1796)? { N1030, N1785, N1784, N1782, N1780 } : 1'b0;
  assign commit_pkt_o[20:19] = (N1)? { 1'b0, mstatus_r_spp_ } : 
                               (N184)? { N1801, N1800 } : 1'b0;
  assign { mstatus_n[9:9], mstatus_n[4:4], mstatus_n[2:2], mstatus_n[0:0] } = (N1)? { 1'b0, 1'b0, 1'b1, mstatus_r_spie_ } : 
                                                                              (N184)? { N1802, N1783, N1781, N1779 } : 1'b0;
  assign fcsr_n[4:0] = (N91)? { N1829, N1830, N1831, N1832, N1833 } : 
                       (N92)? { N972, N971, N970, N969, N968 } : 1'b0;
  assign N91 = N1828;
  assign N92 = N2173;
  assign mcycle_n = (N93)? { N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865 } : 
                    (N1864)? { N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201 } : 1'b0;
  assign N93 = N1863;
  assign minstret_n = (N94)? { N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940 } : 
                      (N1939)? { N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973 } : 1'b0;
  assign N94 = N1938;
  assign { N2045, N2044, N2043, N2042, N2041, N2040 } = (N95)? { N2033, csr_data_lo } : 
                                                        (N96)? { N2034, csr_data_lo } : 
                                                        (N97)? { csr_data_lo_9, N2035, N2036, N2037, N2038, N2039 } : 
                                                        (N2032)? { csr_data_lo_9, csr_data_lo } : 1'b0;
  assign N95 = N2012;
  assign N96 = N2018;
  assign N97 = N2029;
  assign { csr_r_data_o[9:9], csr_r_data_o[4:0] } = (N98)? { N2045, N2044, N2043, N2042, N2041, N2040 } : 
                                                    (N2006)? { csr_data_lo_9, csr_data_lo } : 1'b0;
  assign N98 = N2005;
  assign decode_info_o[10] = decode_info_o[9] | N2071;
  assign sstatus_lo[63] = N2053 & 1'b1;
  assign sstatus_lo[62] = 1'b0 & 1'b0;
  assign sstatus_lo[61] = 1'b0 & 1'b0;
  assign sstatus_lo[60] = 1'b0 & 1'b0;
  assign sstatus_lo[59] = 1'b0 & 1'b0;
  assign sstatus_lo[58] = 1'b0 & 1'b0;
  assign sstatus_lo[57] = 1'b0 & 1'b0;
  assign sstatus_lo[56] = 1'b0 & 1'b0;
  assign sstatus_lo[55] = 1'b0 & 1'b0;
  assign sstatus_lo[54] = 1'b0 & 1'b0;
  assign sstatus_lo[53] = 1'b0 & 1'b0;
  assign sstatus_lo[52] = 1'b0 & 1'b0;
  assign sstatus_lo[51] = 1'b0 & 1'b0;
  assign sstatus_lo[50] = 1'b0 & 1'b0;
  assign sstatus_lo[49] = 1'b0 & 1'b0;
  assign sstatus_lo[48] = 1'b0 & 1'b0;
  assign sstatus_lo[47] = 1'b0 & 1'b0;
  assign sstatus_lo[46] = 1'b0 & 1'b0;
  assign sstatus_lo[45] = 1'b0 & 1'b0;
  assign sstatus_lo[44] = 1'b0 & 1'b0;
  assign sstatus_lo[43] = 1'b0 & 1'b0;
  assign sstatus_lo[42] = 1'b0 & 1'b0;
  assign sstatus_lo[41] = 1'b0 & 1'b0;
  assign sstatus_lo[40] = 1'b0 & 1'b0;
  assign sstatus_lo[39] = 1'b0 & 1'b0;
  assign sstatus_lo[38] = 1'b0 & 1'b0;
  assign sstatus_lo[37] = 1'b0 & 1'b0;
  assign sstatus_lo[36] = 1'b0 & 1'b0;
  assign sstatus_lo[35] = 1'b1 & 1'b0;
  assign sstatus_lo[34] = 1'b0 & 1'b0;
  assign sstatus_lo[33] = 1'b1 & 1'b1;
  assign sstatus_lo[32] = 1'b0 & 1'b1;
  assign sstatus_lo[31] = 1'b0 & 1'b0;
  assign sstatus_lo[30] = 1'b0 & 1'b0;
  assign sstatus_lo[29] = 1'b0 & 1'b0;
  assign sstatus_lo[28] = 1'b0 & 1'b0;
  assign sstatus_lo[27] = 1'b0 & 1'b0;
  assign sstatus_lo[26] = 1'b0 & 1'b0;
  assign sstatus_lo[25] = 1'b0 & 1'b0;
  assign sstatus_lo[24] = 1'b0 & 1'b0;
  assign sstatus_lo[23] = 1'b0 & 1'b0;
  assign sstatus_lo[22] = decode_info_o[8] & 1'b0;
  assign sstatus_lo[21] = decode_info_o[7] & 1'b0;
  assign sstatus_lo[20] = decode_info_o[6] & 1'b0;
  assign sstatus_lo[19] = trans_info_o[0] & 1'b1;
  assign sstatus_lo[18] = trans_info_o[1] & 1'b1;
  assign sstatus_lo[17] = mstatus_r_mprv_ & 1'b0;
  assign sstatus_lo[16] = 1'b0 & 1'b0;
  assign sstatus_lo[15] = 1'b0 & 1'b0;
  assign sstatus_lo[14] = mstatus_r_fs__1_ & 1'b1;
  assign sstatus_lo[13] = mstatus_r_fs__0_ & 1'b1;
  assign sstatus_lo[12] = mstatus_r_mpp__1_ & 1'b0;
  assign sstatus_lo[11] = mstatus_r_mpp__0_ & 1'b0;
  assign sstatus_lo[10] = 1'b0 & 1'b0;
  assign sstatus_lo[9] = 1'b0 & 1'b0;
  assign sstatus_lo[8] = mstatus_r_spp_ & 1'b1;
  assign sstatus_lo[7] = mstatus_r_mpie_ & 1'b0;
  assign sstatus_lo[6] = 1'b0 & 1'b0;
  assign sstatus_lo[5] = mstatus_r_spie_ & 1'b1;
  assign sstatus_lo[4] = 1'b0 & 1'b0;
  assign sstatus_lo[3] = mstatus_r_mie_ & 1'b0;
  assign sstatus_lo[2] = 1'b0 & 1'b0;
  assign sstatus_lo[1] = mstatus_r_sie_ & 1'b1;
  assign sstatus_lo[0] = 1'b0 & 1'b0;
  assign sie_lo[63] = 1'b0 & 1'b0;
  assign sie_lo[62] = 1'b0 & 1'b0;
  assign sie_lo[61] = 1'b0 & 1'b0;
  assign sie_lo[60] = 1'b0 & 1'b0;
  assign sie_lo[59] = 1'b0 & 1'b0;
  assign sie_lo[58] = 1'b0 & 1'b0;
  assign sie_lo[57] = 1'b0 & 1'b0;
  assign sie_lo[56] = 1'b0 & 1'b0;
  assign sie_lo[55] = 1'b0 & 1'b0;
  assign sie_lo[54] = 1'b0 & 1'b0;
  assign sie_lo[53] = 1'b0 & 1'b0;
  assign sie_lo[52] = 1'b0 & 1'b0;
  assign sie_lo[51] = 1'b0 & 1'b0;
  assign sie_lo[50] = 1'b0 & 1'b0;
  assign sie_lo[49] = 1'b0 & 1'b0;
  assign sie_lo[48] = 1'b0 & 1'b0;
  assign sie_lo[47] = 1'b0 & 1'b0;
  assign sie_lo[46] = 1'b0 & 1'b0;
  assign sie_lo[45] = 1'b0 & 1'b0;
  assign sie_lo[44] = 1'b0 & 1'b0;
  assign sie_lo[43] = 1'b0 & 1'b0;
  assign sie_lo[42] = 1'b0 & 1'b0;
  assign sie_lo[41] = 1'b0 & 1'b0;
  assign sie_lo[40] = 1'b0 & 1'b0;
  assign sie_lo[39] = 1'b0 & 1'b0;
  assign sie_lo[38] = 1'b0 & 1'b0;
  assign sie_lo[37] = 1'b0 & 1'b0;
  assign sie_lo[36] = 1'b0 & 1'b0;
  assign sie_lo[35] = 1'b0 & 1'b0;
  assign sie_lo[34] = 1'b0 & 1'b0;
  assign sie_lo[33] = 1'b0 & 1'b0;
  assign sie_lo[32] = 1'b0 & 1'b0;
  assign sie_lo[31] = 1'b0 & 1'b0;
  assign sie_lo[30] = 1'b0 & 1'b0;
  assign sie_lo[29] = 1'b0 & 1'b0;
  assign sie_lo[28] = 1'b0 & 1'b0;
  assign sie_lo[27] = 1'b0 & 1'b0;
  assign sie_lo[26] = 1'b0 & 1'b0;
  assign sie_lo[25] = 1'b0 & 1'b0;
  assign sie_lo[24] = 1'b0 & 1'b0;
  assign sie_lo[23] = 1'b0 & 1'b0;
  assign sie_lo[22] = 1'b0 & 1'b0;
  assign sie_lo[21] = 1'b0 & 1'b0;
  assign sie_lo[20] = 1'b0 & 1'b0;
  assign sie_lo[19] = 1'b0 & 1'b0;
  assign sie_lo[18] = 1'b0 & 1'b0;
  assign sie_lo[17] = 1'b0 & 1'b0;
  assign sie_lo[16] = 1'b0 & 1'b0;
  assign sie_lo[15] = 1'b0 & 1'b0;
  assign sie_lo[14] = 1'b0 & 1'b0;
  assign sie_lo[13] = 1'b0 & 1'b0;
  assign sie_lo[12] = 1'b0 & 1'b0;
  assign sie_lo[11] = mie_r_meie_ & 1'b0;
  assign sie_lo[10] = 1'b0 & 1'b0;
  assign sie_lo[9] = mie_r_seie_ & mideleg_r_sei_;
  assign sie_lo[8] = 1'b0 & 1'b0;
  assign sie_lo[7] = mie_r_mtie_ & 1'b0;
  assign sie_lo[6] = 1'b0 & 1'b0;
  assign sie_lo[5] = mie_r_stie_ & mideleg_r_sti_;
  assign sie_lo[4] = 1'b0 & 1'b0;
  assign sie_lo[3] = mie_r_msie_ & 1'b0;
  assign sie_lo[2] = 1'b0 & 1'b0;
  assign sie_lo[1] = mie_r_ssie_ & mideleg_r_ssi_;
  assign sie_lo[0] = 1'b0 & 1'b0;
  assign sip_lo[63] = 1'b0 & 1'b0;
  assign sip_lo[62] = 1'b0 & 1'b0;
  assign sip_lo[61] = 1'b0 & 1'b0;
  assign sip_lo[60] = 1'b0 & 1'b0;
  assign sip_lo[59] = 1'b0 & 1'b0;
  assign sip_lo[58] = 1'b0 & 1'b0;
  assign sip_lo[57] = 1'b0 & 1'b0;
  assign sip_lo[56] = 1'b0 & 1'b0;
  assign sip_lo[55] = 1'b0 & 1'b0;
  assign sip_lo[54] = 1'b0 & 1'b0;
  assign sip_lo[53] = 1'b0 & 1'b0;
  assign sip_lo[52] = 1'b0 & 1'b0;
  assign sip_lo[51] = 1'b0 & 1'b0;
  assign sip_lo[50] = 1'b0 & 1'b0;
  assign sip_lo[49] = 1'b0 & 1'b0;
  assign sip_lo[48] = 1'b0 & 1'b0;
  assign sip_lo[47] = 1'b0 & 1'b0;
  assign sip_lo[46] = 1'b0 & 1'b0;
  assign sip_lo[45] = 1'b0 & 1'b0;
  assign sip_lo[44] = 1'b0 & 1'b0;
  assign sip_lo[43] = 1'b0 & 1'b0;
  assign sip_lo[42] = 1'b0 & 1'b0;
  assign sip_lo[41] = 1'b0 & 1'b0;
  assign sip_lo[40] = 1'b0 & 1'b0;
  assign sip_lo[39] = 1'b0 & 1'b0;
  assign sip_lo[38] = 1'b0 & 1'b0;
  assign sip_lo[37] = 1'b0 & 1'b0;
  assign sip_lo[36] = 1'b0 & 1'b0;
  assign sip_lo[35] = 1'b0 & 1'b0;
  assign sip_lo[34] = 1'b0 & 1'b0;
  assign sip_lo[33] = 1'b0 & 1'b0;
  assign sip_lo[32] = 1'b0 & 1'b0;
  assign sip_lo[31] = 1'b0 & 1'b0;
  assign sip_lo[30] = 1'b0 & 1'b0;
  assign sip_lo[29] = 1'b0 & 1'b0;
  assign sip_lo[28] = 1'b0 & 1'b0;
  assign sip_lo[27] = 1'b0 & 1'b0;
  assign sip_lo[26] = 1'b0 & 1'b0;
  assign sip_lo[25] = 1'b0 & 1'b0;
  assign sip_lo[24] = 1'b0 & 1'b0;
  assign sip_lo[23] = 1'b0 & 1'b0;
  assign sip_lo[22] = 1'b0 & 1'b0;
  assign sip_lo[21] = 1'b0 & 1'b0;
  assign sip_lo[20] = 1'b0 & 1'b0;
  assign sip_lo[19] = 1'b0 & 1'b0;
  assign sip_lo[18] = 1'b0 & 1'b0;
  assign sip_lo[17] = 1'b0 & 1'b0;
  assign sip_lo[16] = 1'b0 & 1'b0;
  assign sip_lo[15] = 1'b0 & 1'b0;
  assign sip_lo[14] = 1'b0 & 1'b0;
  assign sip_lo[13] = 1'b0 & 1'b0;
  assign sip_lo[12] = 1'b0 & 1'b0;
  assign sip_lo[11] = mip_r_meip_ & 1'b0;
  assign sip_lo[10] = 1'b0 & 1'b0;
  assign sip_lo[9] = mip_r_seip_ & mideleg_r_sei_;
  assign sip_lo[8] = 1'b0 & 1'b0;
  assign sip_lo[7] = mip_r_mtip_ & 1'b0;
  assign sip_lo[6] = 1'b0 & 1'b0;
  assign sip_lo[5] = mip_r_stip_ & mideleg_r_sti_;
  assign sip_lo[4] = 1'b0 & 1'b0;
  assign sip_lo[3] = mip_r_msip_ & 1'b0;
  assign sip_lo[2] = 1'b0 & 1'b0;
  assign sip_lo[1] = mip_r_ssip_ & mideleg_r_ssi_;
  assign sip_lo[0] = 1'b0 & 1'b0;
  assign dgie = ~decode_info_o[9];
  assign mgie = N2075 | decode_info_o[12];
  assign N2075 = N2074 | decode_info_o[11];
  assign N2074 = N2072 & N2073;
  assign N2072 = ~decode_info_o[9];
  assign N2073 = mstatus_r_mie_ & decode_info_o[10];
  assign sgie = N2077 | decode_info_o[12];
  assign N2077 = N2072 & N2076;
  assign N2076 = mstatus_r_sie_ & decode_info_o[11];
  assign interrupt_icode_dec_li_7 = mie_r_mtie_ & mip_r_mtip_;
  assign interrupt_icode_dec_li_3 = mie_r_msie_ & mip_r_msip_;
  assign interrupt_icode_dec_li[11] = mie_r_meie_ & mip_r_meip_;
  assign interrupt_icode_dec_li_5 = mie_r_stie_ & mip_r_stip_;
  assign interrupt_icode_dec_li_1 = mie_r_ssie_ & mip_r_ssip_;
  assign interrupt_icode_dec_li_9 = mie_r_seie_ & N2078;
  assign N2078 = mip_r_seip_ | s_external_irq_i;
  assign irq_waiting_o = N2092 | 1'b0;
  assign N2092 = N2091 | interrupt_icode_dec_li_1;
  assign N2091 = N2090 | 1'b0;
  assign N2090 = N2089 | interrupt_icode_dec_li_3;
  assign N2089 = N2088 | 1'b0;
  assign N2088 = N2087 | interrupt_icode_dec_li_5;
  assign N2087 = N2086 | 1'b0;
  assign N2086 = N2085 | interrupt_icode_dec_li_7;
  assign N2085 = N2084 | 1'b0;
  assign N2084 = N2083 | interrupt_icode_dec_li_9;
  assign N2083 = N2082 | 1'b0;
  assign N2082 = N2081 | interrupt_icode_dec_li[11];
  assign N2081 = N2080 | 1'b0;
  assign N2080 = N2079 | 1'b0;
  assign N2079 = 1'b0 | 1'b0;
  assign _0_net__15_ = 1'b0 & N2093;
  assign N2093 = ~1'b0;
  assign _0_net__14_ = 1'b0 & N2094;
  assign N2094 = ~1'b0;
  assign _0_net__13_ = 1'b0 & N2095;
  assign N2095 = ~1'b0;
  assign _0_net__12_ = 1'b0 & N2096;
  assign N2096 = ~1'b0;
  assign _0_net__11_ = interrupt_icode_dec_li[11] & N2097;
  assign N2097 = ~1'b0;
  assign _0_net__10_ = 1'b0 & N2098;
  assign N2098 = ~1'b0;
  assign _0_net__9_ = interrupt_icode_dec_li_9 & N2099;
  assign N2099 = ~mideleg_r_sei_;
  assign _0_net__8_ = 1'b0 & N2100;
  assign N2100 = ~1'b0;
  assign _0_net__7_ = interrupt_icode_dec_li_7 & N2101;
  assign N2101 = ~1'b0;
  assign _0_net__6_ = 1'b0 & N2102;
  assign N2102 = ~1'b0;
  assign _0_net__5_ = interrupt_icode_dec_li_5 & N2103;
  assign N2103 = ~mideleg_r_sti_;
  assign _0_net__4_ = 1'b0 & N2104;
  assign N2104 = ~1'b0;
  assign _0_net__3_ = interrupt_icode_dec_li_3 & N2105;
  assign N2105 = ~1'b0;
  assign _0_net__2_ = 1'b0 & N2106;
  assign N2106 = ~1'b0;
  assign _0_net__1_ = interrupt_icode_dec_li_1 & N2107;
  assign N2107 = ~mideleg_r_ssi_;
  assign _0_net__0_ = 1'b0 & N2108;
  assign N2108 = ~1'b0;
  assign _1_net__15_ = 1'b0 & 1'b0;
  assign _1_net__14_ = 1'b0 & 1'b0;
  assign _1_net__13_ = 1'b0 & 1'b0;
  assign _1_net__12_ = 1'b0 & 1'b0;
  assign _1_net__11_ = interrupt_icode_dec_li[11] & 1'b0;
  assign _1_net__10_ = 1'b0 & 1'b0;
  assign _1_net__9_ = interrupt_icode_dec_li_9 & mideleg_r_sei_;
  assign _1_net__8_ = 1'b0 & 1'b0;
  assign _1_net__7_ = interrupt_icode_dec_li_7 & 1'b0;
  assign _1_net__6_ = 1'b0 & 1'b0;
  assign _1_net__5_ = interrupt_icode_dec_li_5 & mideleg_r_sti_;
  assign _1_net__4_ = 1'b0 & 1'b0;
  assign _1_net__3_ = interrupt_icode_dec_li_3 & 1'b0;
  assign _1_net__2_ = 1'b0 & 1'b0;
  assign _1_net__1_ = interrupt_icode_dec_li_1 & mideleg_r_ssi_;
  assign _1_net__0_ = 1'b0 & 1'b0;
  assign N182 = retire_pkt_i[5] | retire_pkt_i[4];
  assign N183 = ~N182;
  assign N184 = ~retire_pkt_i[4];
  assign N185 = retire_pkt_i[5] & N184;
  assign N186 = N2065 | decode_info_o[9];
  assign N187 = ~N186;
  assign N188 = ~decode_info_o[9];
  assign N189 = N2065 & N188;
  assign N190 = commit_pkt_o[17] | interrupt_v_lo;
  assign N191 = commit_pkt_o[14] | N190;
  assign N192 = commit_pkt_o_211_ | N191;
  assign N193 = ~N192;
  assign N194 = ~N190;
  assign N195 = commit_pkt_o[14] & N194;
  assign N196 = ~commit_pkt_o[14];
  assign N197 = N194 & N196;
  assign N198 = commit_pkt_o_211_ & N197;
  assign N199 = enter_debug | cfg_bus_i[60];
  assign N200 = ~N199;
  assign commit_pkt_o[18] = N201 & N2052;
  assign N202 = ~csr_r_addr_i[3];
  assign N204 = ~N203;
  assign N206 = ~N205;
  assign N210 = ~N209;
  assign N212 = ~N211;
  assign N217 = ~N216;
  assign N219 = ~N218;
  assign N221 = ~N220;
  assign N223 = ~N222;
  assign N225 = ~N224;
  assign N227 = ~N226;
  assign N230 = ~N229;
  assign N232 = ~N231;
  assign N234 = ~N233;
  assign N236 = ~N235;
  assign N238 = ~N237;
  assign N241 = ~N240;
  assign N247 = ~N246;
  assign N249 = ~N248;
  assign N251 = ~N250;
  assign N253 = ~N252;
  assign N260 = ~N259;
  assign N262 = ~N261;
  assign N264 = ~N263;
  assign N266 = ~N265;
  assign N268 = ~N267;
  assign N270 = ~N269;
  assign N273 = ~N272;
  assign N278 = ~N277;
  assign N279 = ~csr_r_addr_i[2];
  assign N283 = ~N282;
  assign N285 = ~N284;
  assign N287 = ~N286;
  assign N289 = ~N288;
  assign N290 = ~csr_r_addr_i[6];
  assign N295 = ~N294;
  assign N297 = ~N296;
  assign N298 = ~csr_r_addr_i[11];
  assign N305 = ~N304;
  assign N313 = ~N312;
  assign N316 = ~N315;
  assign N320 = ~N319;
  assign N323 = ~N322;
  assign N324 = ~csr_r_addr_i[10];
  assign N325 = ~csr_r_addr_i[9];
  assign N326 = ~csr_r_addr_i[8];
  assign N327 = ~csr_r_addr_i[7];
  assign N328 = ~csr_r_addr_i[5];
  assign N329 = ~csr_r_addr_i[4];
  assign N330 = ~csr_r_addr_i[1];
  assign N331 = ~csr_r_addr_i[0];
  assign N342 = ~N341;
  assign N343 = N206 | N204;
  assign N344 = N210 | N343;
  assign N345 = N212 | N344;
  assign N346 = N217 | N345;
  assign N347 = N219 | N346;
  assign N348 = N221 | N347;
  assign N349 = N223 | N348;
  assign N350 = N225 | N349;
  assign N351 = N227 | N350;
  assign N352 = N230 | N351;
  assign N353 = N232 | N352;
  assign N354 = N234 | N353;
  assign N355 = N236 | N354;
  assign N356 = N238 | N355;
  assign N357 = N241 | N356;
  assign N358 = N247 | N357;
  assign N359 = N249 | N358;
  assign N360 = N251 | N359;
  assign N361 = N253 | N360;
  assign N362 = N260 | N361;
  assign N363 = N262 | N362;
  assign N364 = N264 | N363;
  assign N365 = N266 | N364;
  assign N366 = N268 | N365;
  assign N367 = N270 | N366;
  assign N368 = N273 | N367;
  assign N369 = N278 | N368;
  assign N370 = N283 | N369;
  assign N371 = N285 | N370;
  assign N372 = N287 | N371;
  assign N373 = N289 | N372;
  assign N374 = N295 | N373;
  assign N375 = N297 | N374;
  assign N376 = N305 | N375;
  assign N377 = N313 | N376;
  assign N378 = N316 | N377;
  assign N379 = N320 | N378;
  assign N380 = N323 | N379;
  assign N381 = N342 | N380;
  assign N382 = ~N381;
  assign N448 = ~commit_pkt_o_11_;
  assign N461 = ~N460;
  assign N474 = ~N473;
  assign N487 = ~N486;
  assign N500 = ~N499;
  assign N513 = ~N512;
  assign N526 = ~N525;
  assign N539 = ~N538;
  assign N540 = ~commit_pkt_o_79_;
  assign N553 = ~N552;
  assign N566 = ~N565;
  assign N579 = ~N578;
  assign N580 = ~commit_pkt_o_83_;
  assign N593 = ~N592;
  assign N606 = ~N605;
  assign N619 = ~N618;
  assign N632 = ~N631;
  assign N645 = ~N644;
  assign N646 = ~commit_pkt_o_84_;
  assign N659 = ~N658;
  assign N672 = ~N671;
  assign N685 = ~N684;
  assign N698 = ~N697;
  assign N711 = ~N710;
  assign N724 = ~N723;
  assign N737 = ~N736;
  assign N750 = ~N749;
  assign N763 = ~N762;
  assign N776 = ~N775;
  assign N789 = ~N788;
  assign N802 = ~N801;
  assign N815 = ~N814;
  assign N828 = ~N827;
  assign N841 = ~N840;
  assign N842 = ~commit_pkt_o_82_;
  assign N855 = ~N854;
  assign N856 = ~commit_pkt_o_81_;
  assign N869 = ~N868;
  assign N882 = ~N881;
  assign N895 = ~N894;
  assign N908 = ~N907;
  assign N909 = N474 | N461;
  assign N910 = N487 | N909;
  assign N911 = N500 | N910;
  assign N912 = N513 | N911;
  assign N913 = N526 | N912;
  assign N914 = N539 | N913;
  assign N915 = N553 | N914;
  assign N916 = N566 | N915;
  assign N917 = N579 | N916;
  assign N918 = N593 | N917;
  assign N919 = N606 | N918;
  assign N920 = N619 | N919;
  assign N921 = N632 | N920;
  assign N922 = N645 | N921;
  assign N923 = N659 | N922;
  assign N924 = N672 | N923;
  assign N925 = N685 | N924;
  assign N926 = N698 | N925;
  assign N927 = N711 | N926;
  assign N928 = N724 | N927;
  assign N929 = N737 | N928;
  assign N930 = N750 | N929;
  assign N931 = N763 | N930;
  assign N932 = N776 | N931;
  assign N933 = N789 | N932;
  assign N934 = N802 | N933;
  assign N935 = N815 | N934;
  assign N936 = N828 | N935;
  assign N937 = N841 | N936;
  assign N938 = N855 | N937;
  assign N939 = N869 | N938;
  assign N940 = N882 | N939;
  assign N941 = N895 | N940;
  assign N942 = N908 | N941;
  assign N943 = ~N942;
  assign N944 = N2110 | N2111;
  assign N2110 = decode_info_o[8] & N2109;
  assign N2109 = ~1'b0;
  assign N2111 = commit_pkt_o_43_ & 1'b0;
  assign N945 = N2113 | N2114;
  assign N2113 = decode_info_o[7] & N2112;
  assign N2112 = ~1'b0;
  assign N2114 = commit_pkt_o_42_ & 1'b0;
  assign N946 = N2116 | N2117;
  assign N2116 = decode_info_o[6] & N2115;
  assign N2115 = ~1'b0;
  assign N2117 = commit_pkt_o_41_ & 1'b0;
  assign N947 = N2119 | N2120;
  assign N2119 = trans_info_o[0] & N2118;
  assign N2118 = ~1'b1;
  assign N2120 = commit_pkt_o_40_ & 1'b1;
  assign N948 = N2121 | N2122;
  assign N2121 = trans_info_o[1] & N2118;
  assign N2122 = commit_pkt_o_39_ & 1'b1;
  assign N949 = N2124 | N2125;
  assign N2124 = mstatus_r_mprv_ & N2123;
  assign N2123 = ~1'b0;
  assign N2125 = commit_pkt_o_38_ & 1'b0;
  assign N950 = N2126 | N2127;
  assign N2126 = mstatus_r_fs__1_ & N2118;
  assign N2127 = commit_pkt_o_35_ & 1'b1;
  assign N951 = N2128 | N2129;
  assign N2128 = mstatus_r_fs__0_ & N2118;
  assign N2129 = commit_pkt_o_34_ & 1'b1;
  assign N952 = N2131 | N2132;
  assign N2131 = mstatus_r_mpp__1_ & N2130;
  assign N2130 = ~1'b0;
  assign N2132 = commit_pkt_o_33_ & 1'b0;
  assign N953 = N2134 | N2135;
  assign N2134 = mstatus_r_mpp__0_ & N2133;
  assign N2133 = ~1'b0;
  assign N2135 = commit_pkt_o_32_ & 1'b0;
  assign N954 = N2136 | N2137;
  assign N2136 = mstatus_r_spp_ & N2118;
  assign N2137 = commit_pkt_o_29_ & 1'b1;
  assign N955 = N2139 | N2140;
  assign N2139 = mstatus_r_mpie_ & N2138;
  assign N2138 = ~1'b0;
  assign N2140 = commit_pkt_o_28_ & 1'b0;
  assign N956 = N2141 | N2142;
  assign N2141 = mstatus_r_spie_ & N2118;
  assign N2142 = commit_pkt_o_26_ & 1'b1;
  assign N957 = N2144 | N2145;
  assign N2144 = mstatus_r_mie_ & N2143;
  assign N2143 = ~1'b0;
  assign N2145 = commit_pkt_o_24_ & 1'b0;
  assign N958 = N2146 | N2147;
  assign N2146 = mstatus_r_sie_ & N2118;
  assign N2147 = commit_pkt_o_22_ & 1'b1;
  assign N959 = N2149 | N2150;
  assign N2149 = mie_r_meie_ & N2148;
  assign N2148 = ~1'b0;
  assign N2150 = commit_pkt_o_32_ & 1'b0;
  assign N960 = N2151 | N2152;
  assign N2151 = mie_r_seie_ & N2099;
  assign N2152 = commit_pkt_o_30_ & mideleg_r_sei_;
  assign N961 = N2154 | N2155;
  assign N2154 = mie_r_mtie_ & N2153;
  assign N2153 = ~1'b0;
  assign N2155 = commit_pkt_o_28_ & 1'b0;
  assign N962 = N2156 | N2157;
  assign N2156 = mie_r_stie_ & N2103;
  assign N2157 = commit_pkt_o_26_ & mideleg_r_sti_;
  assign N963 = N2159 | N2160;
  assign N2159 = mie_r_msie_ & N2158;
  assign N2158 = ~1'b0;
  assign N2160 = commit_pkt_o_24_ & 1'b0;
  assign N964 = N2161 | N2162;
  assign N2161 = mie_r_ssie_ & N2107;
  assign N2162 = commit_pkt_o_22_ & mideleg_r_ssi_;
  assign N965 = N2164 | N2165;
  assign N2164 = mip_r_seip_ & N2163;
  assign N2163 = ~1'b0;
  assign N2165 = commit_pkt_o_30_ & 1'b0;
  assign N966 = N2167 | N2168;
  assign N2167 = mip_r_stip_ & N2166;
  assign N2166 = ~1'b0;
  assign N2168 = commit_pkt_o_26_ & 1'b0;
  assign N967 = N2169 | N2170;
  assign N2169 = mip_r_ssip_ & N2107;
  assign N2170 = commit_pkt_o_22_ & mideleg_r_ssi_;
  assign N1295 = exception_ecode_v_li | retire_pkt_i[13];
  assign N1296 = ~N1295;
  assign N1297 = m_interrupt_icode_v_li & mgie;
  assign N1298 = s_interrupt_icode_v_li & sgie;
  assign N1299 = N1298 | N1297;
  assign N1300 = ~N1299;
  assign N1304 = ~N1297;
  assign N1482 = ~exception_ecode_li[0];
  assign N1483 = ~exception_ecode_li[1];
  assign N1484 = N1482 & N1483;
  assign N1485 = N1482 & exception_ecode_li[1];
  assign N1486 = exception_ecode_li[0] & N1483;
  assign N1487 = exception_ecode_li[0] & exception_ecode_li[1];
  assign N1488 = ~exception_ecode_li[2];
  assign N1489 = N1484 & N1488;
  assign N1490 = N1484 & exception_ecode_li[2];
  assign N1491 = N1486 & N1488;
  assign N1492 = N1486 & exception_ecode_li[2];
  assign N1493 = N1485 & N1488;
  assign N1494 = N1485 & exception_ecode_li[2];
  assign N1495 = N1487 & N1488;
  assign N1496 = N1487 & exception_ecode_li[2];
  assign N1497 = ~exception_ecode_li[3];
  assign N1498 = N1489 & N1497;
  assign N1499 = N1489 & exception_ecode_li[3];
  assign N1500 = N1491 & N1497;
  assign N1501 = N1491 & exception_ecode_li[3];
  assign N1502 = N1493 & N1497;
  assign N1503 = N1493 & exception_ecode_li[3];
  assign N1504 = N1495 & N1497;
  assign N1505 = N1495 & exception_ecode_li[3];
  assign N1506 = N1490 & N1497;
  assign N1507 = N1490 & exception_ecode_li[3];
  assign N1508 = N1492 & N1497;
  assign N1509 = N1492 & exception_ecode_li[3];
  assign N1510 = N1494 & N1497;
  assign N1511 = N1494 & exception_ecode_li[3];
  assign N1512 = N1496 & N1497;
  assign N1513 = N1496 & exception_ecode_li[3];
  assign N1515 = N1514 & N2171;
  assign N2171 = ~decode_info_o[10];
  assign N1516 = N1515 | decode_info_o[9];
  assign N1517 = ~N1516;
  assign N1786 = ~retire_pkt_i[13];
  assign N1787 = N2172 & dgie;
  assign N2172 = retire_pkt_i[13] & debug_irq_i;
  assign N1788 = retire_pkt_i[218] & dcsr_r_step_;
  assign N1789 = N1787 | decode_info_o[9];
  assign N1790 = retire_pkt_i[7] | N1789;
  assign N1791 = N1788 | N1790;
  assign N1792 = ~N1791;
  assign exit_debug = retire_pkt_i[6];
  assign N1793 = ~exit_debug;
  assign N1796 = ~retire_pkt_i[5];
  assign N1798 = ~N1797;
  assign N1828 = ~N2173;
  assign N2173 = commit_pkt_o_11_ & N1827;
  assign N1829 = N972 | fflags_acc_i_nv_;
  assign N1830 = N971 | fflags_acc_i_dz_;
  assign N1831 = N970 | fflags_acc_i_of_;
  assign N1832 = N969 | fflags_acc_i_uf_;
  assign N1833 = N968 | fflags_acc_i_nx_;
  assign N1863 = N2175 & N2176;
  assign N2175 = ~N2174;
  assign N2174 = commit_pkt_o_11_ & N1862;
  assign N2176 = ~mcountinhibit_r_cy_;
  assign N1864 = ~N1863;
  assign N1938 = N2178 & N2179;
  assign N2178 = ~N2177;
  assign N2177 = commit_pkt_o_11_ & N1937;
  assign N2179 = ~mcountinhibit_r_ir_;
  assign N1939 = ~N1938;
  assign N1988 = N1029 | N2180;
  assign N2180 = commit_pkt_o_11_ & csr_fany_li;
  assign N1989 = N1028 | N2181;
  assign N2181 = commit_pkt_o_11_ & csr_fany_li;
  assign mstatus_n[8] = N1988 | N2182;
  assign N2182 = commit_pkt_o_211_ & instr_fany_li;
  assign mstatus_n[7] = N1989 | N2183;
  assign N2183 = commit_pkt_o_211_ & instr_fany_li;
  assign N1990 = exception_ecode_v_li & N1786;
  assign N1991 = N1298 & N1304;
  assign N1992 = N1515 & N188;
  assign N1993 = N1787 & N188;
  assign N1994 = ~N1787;
  assign N1995 = N188 & N1994;
  assign N1996 = retire_pkt_i[7] & N1995;
  assign N1997 = ~retire_pkt_i[7];
  assign N1998 = N1995 & N1997;
  assign N1999 = N1788 & N1998;
  assign irq_pending_o = N2185 & N2190;
  assign N2185 = N2184 | dcsr_r_stepie_;
  assign N2184 = ~dcsr_r_step_;
  assign N2190 = N2188 | N2189;
  assign N2188 = N2186 | N2187;
  assign N2186 = debug_irq_i & dgie;
  assign N2187 = m_interrupt_icode_v_li & mgie;
  assign N2189 = s_interrupt_icode_v_li & sgie;
  assign N2000 = ~commit_pkt_o_80_;
  assign N2006 = ~N2005;
  assign N2012 = ~N2011;
  assign N2018 = ~N2017;
  assign N2029 = N2191 | N2192;
  assign N2191 = ~N2023;
  assign N2192 = ~N2028;
  assign N2030 = N2018 | N2012;
  assign N2031 = N2029 | N2030;
  assign N2032 = ~N2031;
  assign N2033 = csr_data_lo_9 | N2193;
  assign N2193 = s_external_irq_i & 1'b0;
  assign N2034 = csr_data_lo_9 | s_external_irq_i;
  assign N2035 = csr_data_lo[4] | fflags_acc_i_nv_;
  assign N2036 = csr_data_lo[3] | fflags_acc_i_dz_;
  assign N2037 = csr_data_lo[2] | fflags_acc_i_of_;
  assign N2038 = csr_data_lo[1] | fflags_acc_i_uf_;
  assign N2039 = csr_data_lo[0] | fflags_acc_i_nx_;
  assign commit_pkt_o[213] = N2225 | retire_pkt_i[11];
  assign N2225 = N2224 | retire_pkt_i[12];
  assign N2224 = N2223 | retire_pkt_i[13];
  assign N2223 = N2222 | commit_pkt_o_2_;
  assign N2222 = N2221 | commit_pkt_o_3_;
  assign N2221 = N2220 | commit_pkt_o_7_;
  assign N2220 = N2219 | commit_pkt_o_6_;
  assign N2219 = N2218 | commit_pkt_o_4_;
  assign N2218 = N2217 | commit_pkt_o_8_;
  assign N2217 = N2216 | commit_pkt_o_9_;
  assign N2216 = N2215 | commit_pkt_o_15_;
  assign N2215 = N2214 | retire_pkt_i[22];
  assign N2214 = N2213 | retire_pkt_i[23];
  assign N2213 = N2212 | retire_pkt_i[24];
  assign N2212 = N2211 | retire_pkt_i[25];
  assign N2211 = N2210 | retire_pkt_i[26];
  assign N2210 = N2209 | retire_pkt_i[27];
  assign N2209 = N2208 | retire_pkt_i[28];
  assign N2208 = N2207 | retire_pkt_i[29];
  assign N2207 = N2206 | retire_pkt_i[30];
  assign N2206 = N2205 | retire_pkt_i[31];
  assign N2205 = N2204 | retire_pkt_i[32];
  assign N2204 = N2203 | retire_pkt_i[33];
  assign N2203 = N2202 | retire_pkt_i[34];
  assign N2202 = N2201 | retire_pkt_i[35];
  assign N2201 = N2200 | commit_pkt_o_11_;
  assign N2200 = N2199 | commit_pkt_o_10_;
  assign N2199 = N2198 | retire_pkt_i[4];
  assign N2198 = N2197 | retire_pkt_i[5];
  assign N2197 = N2196 | retire_pkt_i[6];
  assign N2196 = N2195 | retire_pkt_i[7];
  assign N2195 = N2194 | commit_pkt_o_12_;
  assign N2194 = commit_pkt_o_5_ | commit_pkt_o_13_;
  assign commit_pkt_o[212] = retire_pkt_i[218] & N2250;
  assign N2250 = ~N2249;
  assign N2249 = N2248 | retire_pkt_i[11];
  assign N2248 = N2247 | retire_pkt_i[12];
  assign N2247 = N2246 | retire_pkt_i[13];
  assign N2246 = N2245 | commit_pkt_o_2_;
  assign N2245 = N2244 | commit_pkt_o_3_;
  assign N2244 = N2243 | commit_pkt_o_7_;
  assign N2243 = N2242 | commit_pkt_o_6_;
  assign N2242 = N2241 | commit_pkt_o_4_;
  assign N2241 = N2240 | commit_pkt_o_8_;
  assign N2240 = N2239 | commit_pkt_o_9_;
  assign N2239 = N2238 | commit_pkt_o_15_;
  assign N2238 = N2237 | retire_pkt_i[22];
  assign N2237 = N2236 | retire_pkt_i[23];
  assign N2236 = N2235 | retire_pkt_i[24];
  assign N2235 = N2234 | retire_pkt_i[25];
  assign N2234 = N2233 | retire_pkt_i[26];
  assign N2233 = N2232 | retire_pkt_i[27];
  assign N2232 = N2231 | retire_pkt_i[28];
  assign N2231 = N2230 | retire_pkt_i[29];
  assign N2230 = N2229 | retire_pkt_i[30];
  assign N2229 = N2228 | retire_pkt_i[31];
  assign N2228 = N2227 | retire_pkt_i[32];
  assign N2227 = N2226 | retire_pkt_i[33];
  assign N2226 = retire_pkt_i[35] | retire_pkt_i[34];
  assign commit_pkt_o[16] = interrupt_v_lo | enter_debug;
  assign commit_pkt_o[14] = N2251 | retire_pkt_i[4];
  assign N2251 = retire_pkt_i[6] | retire_pkt_i[5];
  assign trans_info_o[2] = translation_en_r | N2255;
  assign N2255 = N2254 & satp_r_mode_;
  assign N2254 = N2253 & N2046;
  assign N2253 = N2252 & mstatus_r_mprv_;
  assign N2252 = N2072 | dcsr_r_mprven_;
  assign decode_info_o[1] = N2257 | N2258;
  assign N2257 = decode_info_o[10] | N2256;
  assign N2256 = decode_info_o[11] & mcounteren_r_cy_;
  assign N2258 = decode_info_o[12] & scounteren_r_cy_;
  assign decode_info_o[0] = N2260 | N2261;
  assign N2260 = decode_info_o[10] | N2259;
  assign N2259 = decode_info_o[10] & mcounteren_r_ir_;
  assign N2261 = decode_info_o[12] & mcounteren_r_ir_;

endmodule



module bp_be_pipe_sys_00
(
  clk_i,
  reset_i,
  cfg_bus_i,
  reservation_i,
  flush_i,
  retire_v_i,
  retire_queue_v_i,
  retire_data_i,
  retire_exception_i,
  retire_special_i,
  data_o,
  v_o,
  illegal_instr_o,
  iwb_pkt_i,
  fwb_pkt_i,
  commit_pkt_o,
  debug_irq_i,
  timer_irq_i,
  software_irq_i,
  m_external_irq_i,
  s_external_irq_i,
  irq_pending_o,
  irq_waiting_o,
  decode_info_o,
  trans_info_o,
  frm_dyn_o
);

  input [60:0] cfg_bus_i;
  input [520:0] reservation_i;
  input [65:0] retire_data_i;
  input [24:0] retire_exception_i;
  input [8:0] retire_special_i;
  output [65:0] data_o;
  input [78:0] iwb_pkt_i;
  input [78:0] fwb_pkt_i;
  output [213:0] commit_pkt_o;
  output [12:0] decode_info_o;
  output [32:0] trans_info_o;
  output [2:0] frm_dyn_o;
  input clk_i;
  input reset_i;
  input flush_i;
  input retire_v_i;
  input retire_queue_v_i;
  input debug_irq_i;
  input timer_irq_i;
  input software_irq_i;
  input m_external_irq_i;
  input s_external_irq_i;
  output v_o;
  output illegal_instr_o;
  output irq_pending_o;
  output irq_waiting_o;
  wire [65:0] data_o;
  wire [213:0] commit_pkt_o;
  wire [12:0] decode_info_o;
  wire [32:0] trans_info_o;
  wire [2:0] frm_dyn_o,retire_ncount_r,retire_count_r;
  wire v_o,illegal_instr_o,irq_pending_o,irq_waiting_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,
  N10,N11,N12,N13,N14,N15,retire_pkt_instret_,
  retire_pkt_exception__store_page_fault_,retire_pkt_exception__load_page_fault_,
  retire_pkt_exception__instr_page_fault_,retire_pkt_exception__ecall_m_,retire_pkt_exception__ecall_s_,
  retire_pkt_exception__ecall_u_,retire_pkt_exception__store_access_fault_,
  retire_pkt_exception__store_misaligned_,retire_pkt_exception__load_access_fault_,
  retire_pkt_exception__load_misaligned_,retire_pkt_exception__ebreak_,
  retire_pkt_exception__illegal_instr_,retire_pkt_exception__instr_access_fault_,
  retire_pkt_exception__instr_misaligned_,retire_pkt_exception__resume_,retire_pkt_exception__itlb_miss_,
  retire_pkt_exception__icache_miss_,retire_pkt_exception__dcache_replay_,
  retire_pkt_exception__dtlb_load_miss_,retire_pkt_exception__dtlb_store_miss_,
  retire_pkt_exception__itlb_fill_,retire_pkt_exception__dtlb_fill_,retire_pkt_exception___interrupt_,
  retire_pkt_exception__cmd_full_,retire_pkt_exception__mispredict_,
  retire_pkt_special__dcache_miss_,retire_pkt_special__fencei_,retire_pkt_special__sfence_vma_,
  retire_pkt_special__dbreak_,retire_pkt_special__dret_,retire_pkt_special__mret_,
  retire_pkt_special__sret_,retire_pkt_special__wfi_,retire_pkt_special__csrw_,
  retire_pkt_iscore_,retire_pkt_fscore_,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,
  N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,
  N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,
  N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,retire_niscore_r,
  retire_iscore_r,N81,retire_nfscore_r,retire_fscore_r,N82,retire_nspec_w_r,retire_spec_w_r,
  N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,iscore_li,
  fscore_li,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,
  N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,
  N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,
  N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,
  N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,
  N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
  N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
  N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,
  N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,
  N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
  N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,
  N610,N611,N612,N613,N614,N615,N616,N617,N618,N619;
  wire [4:0] fflags_acc_li;
  wire [38:0] retire_npc_r;
  wire [63:0] retire_nvaddr_r,retire_vaddr_r,retire_data_li;
  wire [1:0] retire_nsize_r,retire_size_r;
  wire [31:0] retire_ninstr_r,retire_instr_r;
  reg retire_npc_r_38_sv2v_reg,retire_npc_r_37_sv2v_reg,retire_npc_r_36_sv2v_reg,
  retire_npc_r_35_sv2v_reg,retire_npc_r_34_sv2v_reg,retire_npc_r_33_sv2v_reg,
  retire_npc_r_32_sv2v_reg,retire_npc_r_31_sv2v_reg,retire_npc_r_30_sv2v_reg,
  retire_npc_r_29_sv2v_reg,retire_npc_r_28_sv2v_reg,retire_npc_r_27_sv2v_reg,
  retire_npc_r_26_sv2v_reg,retire_npc_r_25_sv2v_reg,retire_npc_r_24_sv2v_reg,retire_npc_r_23_sv2v_reg,
  retire_npc_r_22_sv2v_reg,retire_npc_r_21_sv2v_reg,retire_npc_r_20_sv2v_reg,
  retire_npc_r_19_sv2v_reg,retire_npc_r_18_sv2v_reg,retire_npc_r_17_sv2v_reg,
  retire_npc_r_16_sv2v_reg,retire_npc_r_15_sv2v_reg,retire_npc_r_14_sv2v_reg,
  retire_npc_r_13_sv2v_reg,retire_npc_r_12_sv2v_reg,retire_npc_r_11_sv2v_reg,
  retire_npc_r_10_sv2v_reg,retire_npc_r_9_sv2v_reg,retire_npc_r_8_sv2v_reg,retire_npc_r_7_sv2v_reg,
  retire_npc_r_6_sv2v_reg,retire_npc_r_5_sv2v_reg,retire_npc_r_4_sv2v_reg,
  retire_npc_r_3_sv2v_reg,retire_npc_r_2_sv2v_reg,retire_npc_r_1_sv2v_reg,
  retire_npc_r_0_sv2v_reg,retire_nvaddr_r_63_sv2v_reg,retire_nvaddr_r_62_sv2v_reg,
  retire_nvaddr_r_61_sv2v_reg,retire_nvaddr_r_60_sv2v_reg,retire_nvaddr_r_59_sv2v_reg,
  retire_nvaddr_r_58_sv2v_reg,retire_nvaddr_r_57_sv2v_reg,retire_nvaddr_r_56_sv2v_reg,
  retire_nvaddr_r_55_sv2v_reg,retire_nvaddr_r_54_sv2v_reg,retire_nvaddr_r_53_sv2v_reg,
  retire_nvaddr_r_52_sv2v_reg,retire_nvaddr_r_51_sv2v_reg,retire_nvaddr_r_50_sv2v_reg,
  retire_nvaddr_r_49_sv2v_reg,retire_nvaddr_r_48_sv2v_reg,
  retire_nvaddr_r_47_sv2v_reg,retire_nvaddr_r_46_sv2v_reg,retire_nvaddr_r_45_sv2v_reg,
  retire_nvaddr_r_44_sv2v_reg,retire_nvaddr_r_43_sv2v_reg,retire_nvaddr_r_42_sv2v_reg,
  retire_nvaddr_r_41_sv2v_reg,retire_nvaddr_r_40_sv2v_reg,retire_nvaddr_r_39_sv2v_reg,
  retire_nvaddr_r_38_sv2v_reg,retire_nvaddr_r_37_sv2v_reg,retire_nvaddr_r_36_sv2v_reg,
  retire_nvaddr_r_35_sv2v_reg,retire_nvaddr_r_34_sv2v_reg,retire_nvaddr_r_33_sv2v_reg,
  retire_nvaddr_r_32_sv2v_reg,retire_nvaddr_r_31_sv2v_reg,retire_nvaddr_r_30_sv2v_reg,
  retire_nvaddr_r_29_sv2v_reg,retire_nvaddr_r_28_sv2v_reg,
  retire_nvaddr_r_27_sv2v_reg,retire_nvaddr_r_26_sv2v_reg,retire_nvaddr_r_25_sv2v_reg,
  retire_nvaddr_r_24_sv2v_reg,retire_nvaddr_r_23_sv2v_reg,retire_nvaddr_r_22_sv2v_reg,
  retire_nvaddr_r_21_sv2v_reg,retire_nvaddr_r_20_sv2v_reg,retire_nvaddr_r_19_sv2v_reg,
  retire_nvaddr_r_18_sv2v_reg,retire_nvaddr_r_17_sv2v_reg,retire_nvaddr_r_16_sv2v_reg,
  retire_nvaddr_r_15_sv2v_reg,retire_nvaddr_r_14_sv2v_reg,retire_nvaddr_r_13_sv2v_reg,
  retire_nvaddr_r_12_sv2v_reg,retire_nvaddr_r_11_sv2v_reg,retire_nvaddr_r_10_sv2v_reg,
  retire_nvaddr_r_9_sv2v_reg,retire_nvaddr_r_8_sv2v_reg,retire_nvaddr_r_7_sv2v_reg,
  retire_nvaddr_r_6_sv2v_reg,retire_nvaddr_r_5_sv2v_reg,retire_nvaddr_r_4_sv2v_reg,
  retire_nvaddr_r_3_sv2v_reg,retire_nvaddr_r_2_sv2v_reg,retire_nvaddr_r_1_sv2v_reg,
  retire_nvaddr_r_0_sv2v_reg,retire_vaddr_r_63_sv2v_reg,
  retire_vaddr_r_62_sv2v_reg,retire_vaddr_r_61_sv2v_reg,retire_vaddr_r_60_sv2v_reg,
  retire_vaddr_r_59_sv2v_reg,retire_vaddr_r_58_sv2v_reg,retire_vaddr_r_57_sv2v_reg,
  retire_vaddr_r_56_sv2v_reg,retire_vaddr_r_55_sv2v_reg,retire_vaddr_r_54_sv2v_reg,
  retire_vaddr_r_53_sv2v_reg,retire_vaddr_r_52_sv2v_reg,retire_vaddr_r_51_sv2v_reg,
  retire_vaddr_r_50_sv2v_reg,retire_vaddr_r_49_sv2v_reg,retire_vaddr_r_48_sv2v_reg,
  retire_vaddr_r_47_sv2v_reg,retire_vaddr_r_46_sv2v_reg,retire_vaddr_r_45_sv2v_reg,
  retire_vaddr_r_44_sv2v_reg,retire_vaddr_r_43_sv2v_reg,retire_vaddr_r_42_sv2v_reg,
  retire_vaddr_r_41_sv2v_reg,retire_vaddr_r_40_sv2v_reg,retire_vaddr_r_39_sv2v_reg,
  retire_vaddr_r_38_sv2v_reg,retire_vaddr_r_37_sv2v_reg,retire_vaddr_r_36_sv2v_reg,
  retire_vaddr_r_35_sv2v_reg,retire_vaddr_r_34_sv2v_reg,retire_vaddr_r_33_sv2v_reg,
  retire_vaddr_r_32_sv2v_reg,retire_vaddr_r_31_sv2v_reg,retire_vaddr_r_30_sv2v_reg,
  retire_vaddr_r_29_sv2v_reg,retire_vaddr_r_28_sv2v_reg,retire_vaddr_r_27_sv2v_reg,
  retire_vaddr_r_26_sv2v_reg,retire_vaddr_r_25_sv2v_reg,retire_vaddr_r_24_sv2v_reg,
  retire_vaddr_r_23_sv2v_reg,retire_vaddr_r_22_sv2v_reg,retire_vaddr_r_21_sv2v_reg,
  retire_vaddr_r_20_sv2v_reg,retire_vaddr_r_19_sv2v_reg,retire_vaddr_r_18_sv2v_reg,
  retire_vaddr_r_17_sv2v_reg,retire_vaddr_r_16_sv2v_reg,retire_vaddr_r_15_sv2v_reg,
  retire_vaddr_r_14_sv2v_reg,retire_vaddr_r_13_sv2v_reg,retire_vaddr_r_12_sv2v_reg,
  retire_vaddr_r_11_sv2v_reg,retire_vaddr_r_10_sv2v_reg,retire_vaddr_r_9_sv2v_reg,
  retire_vaddr_r_8_sv2v_reg,retire_vaddr_r_7_sv2v_reg,retire_vaddr_r_6_sv2v_reg,
  retire_vaddr_r_5_sv2v_reg,retire_vaddr_r_4_sv2v_reg,retire_vaddr_r_3_sv2v_reg,
  retire_vaddr_r_2_sv2v_reg,retire_vaddr_r_1_sv2v_reg,retire_vaddr_r_0_sv2v_reg,
  retire_nsize_r_1_sv2v_reg,retire_nsize_r_0_sv2v_reg,retire_size_r_1_sv2v_reg,
  retire_size_r_0_sv2v_reg,retire_ncount_r_2_sv2v_reg,retire_ncount_r_1_sv2v_reg,
  retire_ncount_r_0_sv2v_reg,retire_count_r_2_sv2v_reg,retire_count_r_1_sv2v_reg,
  retire_count_r_0_sv2v_reg,retire_ninstr_r_31_sv2v_reg,retire_ninstr_r_30_sv2v_reg,
  retire_ninstr_r_29_sv2v_reg,retire_ninstr_r_28_sv2v_reg,retire_ninstr_r_27_sv2v_reg,
  retire_ninstr_r_26_sv2v_reg,retire_ninstr_r_25_sv2v_reg,retire_ninstr_r_24_sv2v_reg,
  retire_ninstr_r_23_sv2v_reg,retire_ninstr_r_22_sv2v_reg,retire_ninstr_r_21_sv2v_reg,
  retire_ninstr_r_20_sv2v_reg,retire_ninstr_r_19_sv2v_reg,retire_ninstr_r_18_sv2v_reg,
  retire_ninstr_r_17_sv2v_reg,retire_ninstr_r_16_sv2v_reg,
  retire_ninstr_r_15_sv2v_reg,retire_ninstr_r_14_sv2v_reg,retire_ninstr_r_13_sv2v_reg,
  retire_ninstr_r_12_sv2v_reg,retire_ninstr_r_11_sv2v_reg,retire_ninstr_r_10_sv2v_reg,
  retire_ninstr_r_9_sv2v_reg,retire_ninstr_r_8_sv2v_reg,retire_ninstr_r_7_sv2v_reg,
  retire_ninstr_r_6_sv2v_reg,retire_ninstr_r_5_sv2v_reg,retire_ninstr_r_4_sv2v_reg,
  retire_ninstr_r_3_sv2v_reg,retire_ninstr_r_2_sv2v_reg,retire_ninstr_r_1_sv2v_reg,
  retire_ninstr_r_0_sv2v_reg,retire_instr_r_31_sv2v_reg,retire_instr_r_30_sv2v_reg,
  retire_instr_r_29_sv2v_reg,retire_instr_r_28_sv2v_reg,retire_instr_r_27_sv2v_reg,
  retire_instr_r_26_sv2v_reg,retire_instr_r_25_sv2v_reg,retire_instr_r_24_sv2v_reg,
  retire_instr_r_23_sv2v_reg,retire_instr_r_22_sv2v_reg,retire_instr_r_21_sv2v_reg,
  retire_instr_r_20_sv2v_reg,retire_instr_r_19_sv2v_reg,retire_instr_r_18_sv2v_reg,
  retire_instr_r_17_sv2v_reg,retire_instr_r_16_sv2v_reg,retire_instr_r_15_sv2v_reg,
  retire_instr_r_14_sv2v_reg,retire_instr_r_13_sv2v_reg,retire_instr_r_12_sv2v_reg,
  retire_instr_r_11_sv2v_reg,retire_instr_r_10_sv2v_reg,retire_instr_r_9_sv2v_reg,
  retire_instr_r_8_sv2v_reg,retire_instr_r_7_sv2v_reg,retire_instr_r_6_sv2v_reg,
  retire_instr_r_5_sv2v_reg,retire_instr_r_4_sv2v_reg,retire_instr_r_3_sv2v_reg,
  retire_instr_r_2_sv2v_reg,retire_instr_r_1_sv2v_reg,retire_instr_r_0_sv2v_reg,
  retire_niscore_r_sv2v_reg,retire_iscore_r_sv2v_reg,retire_nfscore_r_sv2v_reg,
  retire_fscore_r_sv2v_reg,retire_nspec_w_r_sv2v_reg,retire_spec_w_r_sv2v_reg;
  assign retire_npc_r[38] = retire_npc_r_38_sv2v_reg;
  assign retire_npc_r[37] = retire_npc_r_37_sv2v_reg;
  assign retire_npc_r[36] = retire_npc_r_36_sv2v_reg;
  assign retire_npc_r[35] = retire_npc_r_35_sv2v_reg;
  assign retire_npc_r[34] = retire_npc_r_34_sv2v_reg;
  assign retire_npc_r[33] = retire_npc_r_33_sv2v_reg;
  assign retire_npc_r[32] = retire_npc_r_32_sv2v_reg;
  assign retire_npc_r[31] = retire_npc_r_31_sv2v_reg;
  assign retire_npc_r[30] = retire_npc_r_30_sv2v_reg;
  assign retire_npc_r[29] = retire_npc_r_29_sv2v_reg;
  assign retire_npc_r[28] = retire_npc_r_28_sv2v_reg;
  assign retire_npc_r[27] = retire_npc_r_27_sv2v_reg;
  assign retire_npc_r[26] = retire_npc_r_26_sv2v_reg;
  assign retire_npc_r[25] = retire_npc_r_25_sv2v_reg;
  assign retire_npc_r[24] = retire_npc_r_24_sv2v_reg;
  assign retire_npc_r[23] = retire_npc_r_23_sv2v_reg;
  assign retire_npc_r[22] = retire_npc_r_22_sv2v_reg;
  assign retire_npc_r[21] = retire_npc_r_21_sv2v_reg;
  assign retire_npc_r[20] = retire_npc_r_20_sv2v_reg;
  assign retire_npc_r[19] = retire_npc_r_19_sv2v_reg;
  assign retire_npc_r[18] = retire_npc_r_18_sv2v_reg;
  assign retire_npc_r[17] = retire_npc_r_17_sv2v_reg;
  assign retire_npc_r[16] = retire_npc_r_16_sv2v_reg;
  assign retire_npc_r[15] = retire_npc_r_15_sv2v_reg;
  assign retire_npc_r[14] = retire_npc_r_14_sv2v_reg;
  assign retire_npc_r[13] = retire_npc_r_13_sv2v_reg;
  assign retire_npc_r[12] = retire_npc_r_12_sv2v_reg;
  assign retire_npc_r[11] = retire_npc_r_11_sv2v_reg;
  assign retire_npc_r[10] = retire_npc_r_10_sv2v_reg;
  assign retire_npc_r[9] = retire_npc_r_9_sv2v_reg;
  assign retire_npc_r[8] = retire_npc_r_8_sv2v_reg;
  assign retire_npc_r[7] = retire_npc_r_7_sv2v_reg;
  assign retire_npc_r[6] = retire_npc_r_6_sv2v_reg;
  assign retire_npc_r[5] = retire_npc_r_5_sv2v_reg;
  assign retire_npc_r[4] = retire_npc_r_4_sv2v_reg;
  assign retire_npc_r[3] = retire_npc_r_3_sv2v_reg;
  assign retire_npc_r[2] = retire_npc_r_2_sv2v_reg;
  assign retire_npc_r[1] = retire_npc_r_1_sv2v_reg;
  assign retire_npc_r[0] = retire_npc_r_0_sv2v_reg;
  assign retire_nvaddr_r[63] = retire_nvaddr_r_63_sv2v_reg;
  assign retire_nvaddr_r[62] = retire_nvaddr_r_62_sv2v_reg;
  assign retire_nvaddr_r[61] = retire_nvaddr_r_61_sv2v_reg;
  assign retire_nvaddr_r[60] = retire_nvaddr_r_60_sv2v_reg;
  assign retire_nvaddr_r[59] = retire_nvaddr_r_59_sv2v_reg;
  assign retire_nvaddr_r[58] = retire_nvaddr_r_58_sv2v_reg;
  assign retire_nvaddr_r[57] = retire_nvaddr_r_57_sv2v_reg;
  assign retire_nvaddr_r[56] = retire_nvaddr_r_56_sv2v_reg;
  assign retire_nvaddr_r[55] = retire_nvaddr_r_55_sv2v_reg;
  assign retire_nvaddr_r[54] = retire_nvaddr_r_54_sv2v_reg;
  assign retire_nvaddr_r[53] = retire_nvaddr_r_53_sv2v_reg;
  assign retire_nvaddr_r[52] = retire_nvaddr_r_52_sv2v_reg;
  assign retire_nvaddr_r[51] = retire_nvaddr_r_51_sv2v_reg;
  assign retire_nvaddr_r[50] = retire_nvaddr_r_50_sv2v_reg;
  assign retire_nvaddr_r[49] = retire_nvaddr_r_49_sv2v_reg;
  assign retire_nvaddr_r[48] = retire_nvaddr_r_48_sv2v_reg;
  assign retire_nvaddr_r[47] = retire_nvaddr_r_47_sv2v_reg;
  assign retire_nvaddr_r[46] = retire_nvaddr_r_46_sv2v_reg;
  assign retire_nvaddr_r[45] = retire_nvaddr_r_45_sv2v_reg;
  assign retire_nvaddr_r[44] = retire_nvaddr_r_44_sv2v_reg;
  assign retire_nvaddr_r[43] = retire_nvaddr_r_43_sv2v_reg;
  assign retire_nvaddr_r[42] = retire_nvaddr_r_42_sv2v_reg;
  assign retire_nvaddr_r[41] = retire_nvaddr_r_41_sv2v_reg;
  assign retire_nvaddr_r[40] = retire_nvaddr_r_40_sv2v_reg;
  assign retire_nvaddr_r[39] = retire_nvaddr_r_39_sv2v_reg;
  assign retire_nvaddr_r[38] = retire_nvaddr_r_38_sv2v_reg;
  assign retire_nvaddr_r[37] = retire_nvaddr_r_37_sv2v_reg;
  assign retire_nvaddr_r[36] = retire_nvaddr_r_36_sv2v_reg;
  assign retire_nvaddr_r[35] = retire_nvaddr_r_35_sv2v_reg;
  assign retire_nvaddr_r[34] = retire_nvaddr_r_34_sv2v_reg;
  assign retire_nvaddr_r[33] = retire_nvaddr_r_33_sv2v_reg;
  assign retire_nvaddr_r[32] = retire_nvaddr_r_32_sv2v_reg;
  assign retire_nvaddr_r[31] = retire_nvaddr_r_31_sv2v_reg;
  assign retire_nvaddr_r[30] = retire_nvaddr_r_30_sv2v_reg;
  assign retire_nvaddr_r[29] = retire_nvaddr_r_29_sv2v_reg;
  assign retire_nvaddr_r[28] = retire_nvaddr_r_28_sv2v_reg;
  assign retire_nvaddr_r[27] = retire_nvaddr_r_27_sv2v_reg;
  assign retire_nvaddr_r[26] = retire_nvaddr_r_26_sv2v_reg;
  assign retire_nvaddr_r[25] = retire_nvaddr_r_25_sv2v_reg;
  assign retire_nvaddr_r[24] = retire_nvaddr_r_24_sv2v_reg;
  assign retire_nvaddr_r[23] = retire_nvaddr_r_23_sv2v_reg;
  assign retire_nvaddr_r[22] = retire_nvaddr_r_22_sv2v_reg;
  assign retire_nvaddr_r[21] = retire_nvaddr_r_21_sv2v_reg;
  assign retire_nvaddr_r[20] = retire_nvaddr_r_20_sv2v_reg;
  assign retire_nvaddr_r[19] = retire_nvaddr_r_19_sv2v_reg;
  assign retire_nvaddr_r[18] = retire_nvaddr_r_18_sv2v_reg;
  assign retire_nvaddr_r[17] = retire_nvaddr_r_17_sv2v_reg;
  assign retire_nvaddr_r[16] = retire_nvaddr_r_16_sv2v_reg;
  assign retire_nvaddr_r[15] = retire_nvaddr_r_15_sv2v_reg;
  assign retire_nvaddr_r[14] = retire_nvaddr_r_14_sv2v_reg;
  assign retire_nvaddr_r[13] = retire_nvaddr_r_13_sv2v_reg;
  assign retire_nvaddr_r[12] = retire_nvaddr_r_12_sv2v_reg;
  assign retire_nvaddr_r[11] = retire_nvaddr_r_11_sv2v_reg;
  assign retire_nvaddr_r[10] = retire_nvaddr_r_10_sv2v_reg;
  assign retire_nvaddr_r[9] = retire_nvaddr_r_9_sv2v_reg;
  assign retire_nvaddr_r[8] = retire_nvaddr_r_8_sv2v_reg;
  assign retire_nvaddr_r[7] = retire_nvaddr_r_7_sv2v_reg;
  assign retire_nvaddr_r[6] = retire_nvaddr_r_6_sv2v_reg;
  assign retire_nvaddr_r[5] = retire_nvaddr_r_5_sv2v_reg;
  assign retire_nvaddr_r[4] = retire_nvaddr_r_4_sv2v_reg;
  assign retire_nvaddr_r[3] = retire_nvaddr_r_3_sv2v_reg;
  assign retire_nvaddr_r[2] = retire_nvaddr_r_2_sv2v_reg;
  assign retire_nvaddr_r[1] = retire_nvaddr_r_1_sv2v_reg;
  assign retire_nvaddr_r[0] = retire_nvaddr_r_0_sv2v_reg;
  assign retire_vaddr_r[63] = retire_vaddr_r_63_sv2v_reg;
  assign retire_vaddr_r[62] = retire_vaddr_r_62_sv2v_reg;
  assign retire_vaddr_r[61] = retire_vaddr_r_61_sv2v_reg;
  assign retire_vaddr_r[60] = retire_vaddr_r_60_sv2v_reg;
  assign retire_vaddr_r[59] = retire_vaddr_r_59_sv2v_reg;
  assign retire_vaddr_r[58] = retire_vaddr_r_58_sv2v_reg;
  assign retire_vaddr_r[57] = retire_vaddr_r_57_sv2v_reg;
  assign retire_vaddr_r[56] = retire_vaddr_r_56_sv2v_reg;
  assign retire_vaddr_r[55] = retire_vaddr_r_55_sv2v_reg;
  assign retire_vaddr_r[54] = retire_vaddr_r_54_sv2v_reg;
  assign retire_vaddr_r[53] = retire_vaddr_r_53_sv2v_reg;
  assign retire_vaddr_r[52] = retire_vaddr_r_52_sv2v_reg;
  assign retire_vaddr_r[51] = retire_vaddr_r_51_sv2v_reg;
  assign retire_vaddr_r[50] = retire_vaddr_r_50_sv2v_reg;
  assign retire_vaddr_r[49] = retire_vaddr_r_49_sv2v_reg;
  assign retire_vaddr_r[48] = retire_vaddr_r_48_sv2v_reg;
  assign retire_vaddr_r[47] = retire_vaddr_r_47_sv2v_reg;
  assign retire_vaddr_r[46] = retire_vaddr_r_46_sv2v_reg;
  assign retire_vaddr_r[45] = retire_vaddr_r_45_sv2v_reg;
  assign retire_vaddr_r[44] = retire_vaddr_r_44_sv2v_reg;
  assign retire_vaddr_r[43] = retire_vaddr_r_43_sv2v_reg;
  assign retire_vaddr_r[42] = retire_vaddr_r_42_sv2v_reg;
  assign retire_vaddr_r[41] = retire_vaddr_r_41_sv2v_reg;
  assign retire_vaddr_r[40] = retire_vaddr_r_40_sv2v_reg;
  assign retire_vaddr_r[39] = retire_vaddr_r_39_sv2v_reg;
  assign retire_vaddr_r[38] = retire_vaddr_r_38_sv2v_reg;
  assign retire_vaddr_r[37] = retire_vaddr_r_37_sv2v_reg;
  assign retire_vaddr_r[36] = retire_vaddr_r_36_sv2v_reg;
  assign retire_vaddr_r[35] = retire_vaddr_r_35_sv2v_reg;
  assign retire_vaddr_r[34] = retire_vaddr_r_34_sv2v_reg;
  assign retire_vaddr_r[33] = retire_vaddr_r_33_sv2v_reg;
  assign retire_vaddr_r[32] = retire_vaddr_r_32_sv2v_reg;
  assign retire_vaddr_r[31] = retire_vaddr_r_31_sv2v_reg;
  assign retire_vaddr_r[30] = retire_vaddr_r_30_sv2v_reg;
  assign retire_vaddr_r[29] = retire_vaddr_r_29_sv2v_reg;
  assign retire_vaddr_r[28] = retire_vaddr_r_28_sv2v_reg;
  assign retire_vaddr_r[27] = retire_vaddr_r_27_sv2v_reg;
  assign retire_vaddr_r[26] = retire_vaddr_r_26_sv2v_reg;
  assign retire_vaddr_r[25] = retire_vaddr_r_25_sv2v_reg;
  assign retire_vaddr_r[24] = retire_vaddr_r_24_sv2v_reg;
  assign retire_vaddr_r[23] = retire_vaddr_r_23_sv2v_reg;
  assign retire_vaddr_r[22] = retire_vaddr_r_22_sv2v_reg;
  assign retire_vaddr_r[21] = retire_vaddr_r_21_sv2v_reg;
  assign retire_vaddr_r[20] = retire_vaddr_r_20_sv2v_reg;
  assign retire_vaddr_r[19] = retire_vaddr_r_19_sv2v_reg;
  assign retire_vaddr_r[18] = retire_vaddr_r_18_sv2v_reg;
  assign retire_vaddr_r[17] = retire_vaddr_r_17_sv2v_reg;
  assign retire_vaddr_r[16] = retire_vaddr_r_16_sv2v_reg;
  assign retire_vaddr_r[15] = retire_vaddr_r_15_sv2v_reg;
  assign retire_vaddr_r[14] = retire_vaddr_r_14_sv2v_reg;
  assign retire_vaddr_r[13] = retire_vaddr_r_13_sv2v_reg;
  assign retire_vaddr_r[12] = retire_vaddr_r_12_sv2v_reg;
  assign retire_vaddr_r[11] = retire_vaddr_r_11_sv2v_reg;
  assign retire_vaddr_r[10] = retire_vaddr_r_10_sv2v_reg;
  assign retire_vaddr_r[9] = retire_vaddr_r_9_sv2v_reg;
  assign retire_vaddr_r[8] = retire_vaddr_r_8_sv2v_reg;
  assign retire_vaddr_r[7] = retire_vaddr_r_7_sv2v_reg;
  assign retire_vaddr_r[6] = retire_vaddr_r_6_sv2v_reg;
  assign retire_vaddr_r[5] = retire_vaddr_r_5_sv2v_reg;
  assign retire_vaddr_r[4] = retire_vaddr_r_4_sv2v_reg;
  assign retire_vaddr_r[3] = retire_vaddr_r_3_sv2v_reg;
  assign retire_vaddr_r[2] = retire_vaddr_r_2_sv2v_reg;
  assign retire_vaddr_r[1] = retire_vaddr_r_1_sv2v_reg;
  assign retire_vaddr_r[0] = retire_vaddr_r_0_sv2v_reg;
  assign retire_nsize_r[1] = retire_nsize_r_1_sv2v_reg;
  assign retire_nsize_r[0] = retire_nsize_r_0_sv2v_reg;
  assign retire_size_r[1] = retire_size_r_1_sv2v_reg;
  assign retire_size_r[0] = retire_size_r_0_sv2v_reg;
  assign retire_ncount_r[2] = retire_ncount_r_2_sv2v_reg;
  assign retire_ncount_r[1] = retire_ncount_r_1_sv2v_reg;
  assign retire_ncount_r[0] = retire_ncount_r_0_sv2v_reg;
  assign retire_count_r[2] = retire_count_r_2_sv2v_reg;
  assign retire_count_r[1] = retire_count_r_1_sv2v_reg;
  assign retire_count_r[0] = retire_count_r_0_sv2v_reg;
  assign retire_ninstr_r[31] = retire_ninstr_r_31_sv2v_reg;
  assign retire_ninstr_r[30] = retire_ninstr_r_30_sv2v_reg;
  assign retire_ninstr_r[29] = retire_ninstr_r_29_sv2v_reg;
  assign retire_ninstr_r[28] = retire_ninstr_r_28_sv2v_reg;
  assign retire_ninstr_r[27] = retire_ninstr_r_27_sv2v_reg;
  assign retire_ninstr_r[26] = retire_ninstr_r_26_sv2v_reg;
  assign retire_ninstr_r[25] = retire_ninstr_r_25_sv2v_reg;
  assign retire_ninstr_r[24] = retire_ninstr_r_24_sv2v_reg;
  assign retire_ninstr_r[23] = retire_ninstr_r_23_sv2v_reg;
  assign retire_ninstr_r[22] = retire_ninstr_r_22_sv2v_reg;
  assign retire_ninstr_r[21] = retire_ninstr_r_21_sv2v_reg;
  assign retire_ninstr_r[20] = retire_ninstr_r_20_sv2v_reg;
  assign retire_ninstr_r[19] = retire_ninstr_r_19_sv2v_reg;
  assign retire_ninstr_r[18] = retire_ninstr_r_18_sv2v_reg;
  assign retire_ninstr_r[17] = retire_ninstr_r_17_sv2v_reg;
  assign retire_ninstr_r[16] = retire_ninstr_r_16_sv2v_reg;
  assign retire_ninstr_r[15] = retire_ninstr_r_15_sv2v_reg;
  assign retire_ninstr_r[14] = retire_ninstr_r_14_sv2v_reg;
  assign retire_ninstr_r[13] = retire_ninstr_r_13_sv2v_reg;
  assign retire_ninstr_r[12] = retire_ninstr_r_12_sv2v_reg;
  assign retire_ninstr_r[11] = retire_ninstr_r_11_sv2v_reg;
  assign retire_ninstr_r[10] = retire_ninstr_r_10_sv2v_reg;
  assign retire_ninstr_r[9] = retire_ninstr_r_9_sv2v_reg;
  assign retire_ninstr_r[8] = retire_ninstr_r_8_sv2v_reg;
  assign retire_ninstr_r[7] = retire_ninstr_r_7_sv2v_reg;
  assign retire_ninstr_r[6] = retire_ninstr_r_6_sv2v_reg;
  assign retire_ninstr_r[5] = retire_ninstr_r_5_sv2v_reg;
  assign retire_ninstr_r[4] = retire_ninstr_r_4_sv2v_reg;
  assign retire_ninstr_r[3] = retire_ninstr_r_3_sv2v_reg;
  assign retire_ninstr_r[2] = retire_ninstr_r_2_sv2v_reg;
  assign retire_ninstr_r[1] = retire_ninstr_r_1_sv2v_reg;
  assign retire_ninstr_r[0] = retire_ninstr_r_0_sv2v_reg;
  assign retire_instr_r[31] = retire_instr_r_31_sv2v_reg;
  assign retire_instr_r[30] = retire_instr_r_30_sv2v_reg;
  assign retire_instr_r[29] = retire_instr_r_29_sv2v_reg;
  assign retire_instr_r[28] = retire_instr_r_28_sv2v_reg;
  assign retire_instr_r[27] = retire_instr_r_27_sv2v_reg;
  assign retire_instr_r[26] = retire_instr_r_26_sv2v_reg;
  assign retire_instr_r[25] = retire_instr_r_25_sv2v_reg;
  assign retire_instr_r[24] = retire_instr_r_24_sv2v_reg;
  assign retire_instr_r[23] = retire_instr_r_23_sv2v_reg;
  assign retire_instr_r[22] = retire_instr_r_22_sv2v_reg;
  assign retire_instr_r[21] = retire_instr_r_21_sv2v_reg;
  assign retire_instr_r[20] = retire_instr_r_20_sv2v_reg;
  assign retire_instr_r[19] = retire_instr_r_19_sv2v_reg;
  assign retire_instr_r[18] = retire_instr_r_18_sv2v_reg;
  assign retire_instr_r[17] = retire_instr_r_17_sv2v_reg;
  assign retire_instr_r[16] = retire_instr_r_16_sv2v_reg;
  assign retire_instr_r[15] = retire_instr_r_15_sv2v_reg;
  assign retire_instr_r[14] = retire_instr_r_14_sv2v_reg;
  assign retire_instr_r[13] = retire_instr_r_13_sv2v_reg;
  assign retire_instr_r[12] = retire_instr_r_12_sv2v_reg;
  assign retire_instr_r[11] = retire_instr_r_11_sv2v_reg;
  assign retire_instr_r[10] = retire_instr_r_10_sv2v_reg;
  assign retire_instr_r[9] = retire_instr_r_9_sv2v_reg;
  assign retire_instr_r[8] = retire_instr_r_8_sv2v_reg;
  assign retire_instr_r[7] = retire_instr_r_7_sv2v_reg;
  assign retire_instr_r[6] = retire_instr_r_6_sv2v_reg;
  assign retire_instr_r[5] = retire_instr_r_5_sv2v_reg;
  assign retire_instr_r[4] = retire_instr_r_4_sv2v_reg;
  assign retire_instr_r[3] = retire_instr_r_3_sv2v_reg;
  assign retire_instr_r[2] = retire_instr_r_2_sv2v_reg;
  assign retire_instr_r[1] = retire_instr_r_1_sv2v_reg;
  assign retire_instr_r[0] = retire_instr_r_0_sv2v_reg;
  assign retire_niscore_r = retire_niscore_r_sv2v_reg;
  assign retire_iscore_r = retire_iscore_r_sv2v_reg;
  assign retire_nfscore_r = retire_nfscore_r_sv2v_reg;
  assign retire_fscore_r = retire_fscore_r_sv2v_reg;
  assign retire_nspec_w_r = retire_nspec_w_r_sv2v_reg;
  assign retire_spec_w_r = retire_spec_w_r_sv2v_reg;
  assign data_o[64] = 1'b0;
  assign data_o[65] = 1'b0;

  bp_be_csr_00
  csr
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .cfg_bus_i(cfg_bus_i),
    .csr_r_v_i(v_o),
    .csr_r_addr_i(reservation_i[480:469]),
    .csr_r_data_o(data_o[63:0]),
    .csr_r_illegal_o(illegal_instr_o),
    .retire_pkt_i({ retire_v_i, retire_queue_v_i, retire_pkt_instret_, retire_npc_r, retire_vaddr_r[38:0], 1'b0, 1'b0, retire_data_li, retire_instr_r, retire_count_r, retire_size_r, retire_pkt_exception__store_page_fault_, retire_pkt_exception__load_page_fault_, retire_pkt_exception__instr_page_fault_, retire_pkt_exception__ecall_m_, retire_pkt_exception__ecall_s_, retire_pkt_exception__ecall_u_, retire_pkt_exception__store_access_fault_, retire_pkt_exception__store_misaligned_, retire_pkt_exception__load_access_fault_, retire_pkt_exception__load_misaligned_, retire_pkt_exception__ebreak_, retire_pkt_exception__illegal_instr_, retire_pkt_exception__instr_access_fault_, retire_pkt_exception__instr_misaligned_, retire_pkt_exception__resume_, retire_pkt_exception__itlb_miss_, retire_pkt_exception__icache_miss_, retire_pkt_exception__dcache_replay_, retire_pkt_exception__dtlb_load_miss_, retire_pkt_exception__dtlb_store_miss_, retire_pkt_exception__itlb_fill_, retire_pkt_exception__dtlb_fill_, retire_pkt_exception___interrupt_, retire_pkt_exception__cmd_full_, retire_pkt_exception__mispredict_, retire_pkt_special__dcache_miss_, retire_pkt_special__fencei_, retire_pkt_special__sfence_vma_, retire_pkt_special__dbreak_, retire_pkt_special__dret_, retire_pkt_special__mret_, retire_pkt_special__sret_, retire_pkt_special__wfi_, retire_pkt_special__csrw_, retire_pkt_iscore_, retire_pkt_fscore_ }),
    .frf_w_v_i(fwb_pkt_i[77]),
    .debug_irq_i(debug_irq_i),
    .timer_irq_i(timer_irq_i),
    .software_irq_i(software_irq_i),
    .m_external_irq_i(m_external_irq_i),
    .s_external_irq_i(s_external_irq_i),
    .irq_pending_o(irq_pending_o),
    .irq_waiting_o(irq_waiting_o),
    .commit_pkt_o(commit_pkt_o),
    .decode_info_o(decode_info_o),
    .trans_info_o(trans_info_o),
    .frm_dyn_o(frm_dyn_o),
    .fflags_acc_i_nv_(fflags_acc_li[4]),
    .fflags_acc_i_dz_(fflags_acc_li[3]),
    .fflags_acc_i_of_(fflags_acc_li[2]),
    .fflags_acc_i_uf_(fflags_acc_li[1]),
    .fflags_acc_i_nx_(fflags_acc_li[0])
  );

  assign N85 = retire_queue_v_i & retire_instr_r[6];
  assign N86 = retire_instr_r[5] & retire_instr_r[4];
  assign N87 = N83 & N84;
  assign N88 = retire_instr_r[1] & retire_instr_r[0];
  assign N89 = N85 & N86;
  assign N90 = N87 & N88;
  assign N91 = N89 & N90;
  assign N94 = retire_instr_r[14] & retire_instr_r[13];
  assign N95 = N94 & N93;
  assign N96 = retire_instr_r[14] & retire_instr_r[13];
  assign N97 = N96 & retire_instr_r[12];
  assign N99 = retire_instr_r[14] & N98;
  assign N100 = N99 & retire_instr_r[12];
  assign N103 = N101 & retire_instr_r[13];
  assign N104 = N103 & N102;
  assign N106 = N105 & retire_instr_r[13];
  assign N107 = N106 & retire_instr_r[12];
  assign N110 = N108 & N109;
  assign N111 = N110 & retire_instr_r[12];
  assign N114 = N112 & N113;
  assign { N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16 } = reservation_i[388:325] + reservation_i[258:195];
  assign { N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371 } = (N0)? { N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N1)? { N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, retire_instr_r[19:15] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N3)? { N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N4)? { N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N5)? retire_vaddr_r : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N6)? retire_data_i[63:0] : 1'b0;
  assign N0 = N95;
  assign N1 = N97;
  assign N2 = N100;
  assign N3 = N104;
  assign N4 = N107;
  assign N5 = N111;
  assign N6 = N114;
  assign retire_data_li = (N7)? { N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371 } : 
                          (N92)? retire_data_i[63:0] : 1'b0;
  assign N7 = N91;
  assign { retire_pkt_exception__store_page_fault_, retire_pkt_exception__load_page_fault_, retire_pkt_exception__instr_page_fault_, retire_pkt_exception__ecall_m_, retire_pkt_exception__ecall_s_, retire_pkt_exception__ecall_u_, retire_pkt_exception__store_access_fault_, retire_pkt_exception__store_misaligned_, retire_pkt_exception__load_access_fault_, retire_pkt_exception__load_misaligned_, retire_pkt_exception__ebreak_, retire_pkt_exception__illegal_instr_, retire_pkt_exception__instr_access_fault_, retire_pkt_exception__instr_misaligned_, retire_pkt_exception__resume_, retire_pkt_exception__itlb_miss_, retire_pkt_exception__icache_miss_, retire_pkt_exception__dcache_replay_, retire_pkt_exception__dtlb_load_miss_, retire_pkt_exception__dtlb_store_miss_, retire_pkt_exception__itlb_fill_, retire_pkt_exception__dtlb_fill_, retire_pkt_exception___interrupt_, retire_pkt_exception__cmd_full_, retire_pkt_exception__mispredict_ } = (N8)? retire_exception_i : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = N436;
  assign N9 = N435;
  assign { retire_pkt_special__dcache_miss_, retire_pkt_special__fencei_, retire_pkt_special__sfence_vma_, retire_pkt_special__dbreak_, retire_pkt_special__dret_, retire_pkt_special__mret_, retire_pkt_special__sret_, retire_pkt_special__wfi_, retire_pkt_special__csrw_ } = (N10)? retire_special_i : 
                                                                                                                                                                                                                                                                                 (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = N438;
  assign N11 = N437;
  assign retire_pkt_iscore_ = (N12)? iscore_li : 
                              (N13)? 1'b0 : 1'b0;
  assign N12 = N440;
  assign N13 = N439;
  assign retire_pkt_fscore_ = (N14)? fscore_li : 
                              (N15)? 1'b0 : 1'b0;
  assign N14 = N442;
  assign N15 = N441;
  assign v_o = reservation_i[424] | reservation_i[425];
  assign fflags_acc_li[4] = iwb_pkt_i[4] | fwb_pkt_i[4];
  assign fflags_acc_li[3] = iwb_pkt_i[3] | fwb_pkt_i[3];
  assign fflags_acc_li[2] = iwb_pkt_i[2] | fwb_pkt_i[2];
  assign fflags_acc_li[1] = iwb_pkt_i[1] | fwb_pkt_i[1];
  assign fflags_acc_li[0] = iwb_pkt_i[0] | fwb_pkt_i[0];
  assign N80 = reservation_i[422] & reservation_i[435];
  assign N81 = reservation_i[422] & reservation_i[434];
  assign N82 = reservation_i[422] & reservation_i[421];
  assign N83 = ~retire_instr_r[3];
  assign N84 = ~retire_instr_r[2];
  assign N92 = ~N91;
  assign N93 = ~retire_instr_r[12];
  assign N98 = ~retire_instr_r[13];
  assign N101 = ~retire_instr_r[14];
  assign N102 = ~retire_instr_r[12];
  assign N105 = ~retire_instr_r[14];
  assign N108 = ~retire_instr_r[14];
  assign N109 = ~retire_instr_r[13];
  assign N112 = ~retire_instr_r[13];
  assign N113 = ~retire_instr_r[12];
  assign N115 = 1'b0 | retire_data_i[63];
  assign N116 = 1'b0 | retire_data_i[62];
  assign N117 = 1'b0 | retire_data_i[61];
  assign N118 = 1'b0 | retire_data_i[60];
  assign N119 = 1'b0 | retire_data_i[59];
  assign N120 = 1'b0 | retire_data_i[58];
  assign N121 = 1'b0 | retire_data_i[57];
  assign N122 = 1'b0 | retire_data_i[56];
  assign N123 = 1'b0 | retire_data_i[55];
  assign N124 = 1'b0 | retire_data_i[54];
  assign N125 = 1'b0 | retire_data_i[53];
  assign N126 = 1'b0 | retire_data_i[52];
  assign N127 = 1'b0 | retire_data_i[51];
  assign N128 = 1'b0 | retire_data_i[50];
  assign N129 = 1'b0 | retire_data_i[49];
  assign N130 = 1'b0 | retire_data_i[48];
  assign N131 = 1'b0 | retire_data_i[47];
  assign N132 = 1'b0 | retire_data_i[46];
  assign N133 = 1'b0 | retire_data_i[45];
  assign N134 = 1'b0 | retire_data_i[44];
  assign N135 = 1'b0 | retire_data_i[43];
  assign N136 = 1'b0 | retire_data_i[42];
  assign N137 = 1'b0 | retire_data_i[41];
  assign N138 = 1'b0 | retire_data_i[40];
  assign N139 = 1'b0 | retire_data_i[39];
  assign N140 = 1'b0 | retire_data_i[38];
  assign N141 = 1'b0 | retire_data_i[37];
  assign N142 = 1'b0 | retire_data_i[36];
  assign N143 = 1'b0 | retire_data_i[35];
  assign N144 = 1'b0 | retire_data_i[34];
  assign N145 = 1'b0 | retire_data_i[33];
  assign N146 = 1'b0 | retire_data_i[32];
  assign N147 = 1'b0 | retire_data_i[31];
  assign N148 = 1'b0 | retire_data_i[30];
  assign N149 = 1'b0 | retire_data_i[29];
  assign N150 = 1'b0 | retire_data_i[28];
  assign N151 = 1'b0 | retire_data_i[27];
  assign N152 = 1'b0 | retire_data_i[26];
  assign N153 = 1'b0 | retire_data_i[25];
  assign N154 = 1'b0 | retire_data_i[24];
  assign N155 = 1'b0 | retire_data_i[23];
  assign N156 = 1'b0 | retire_data_i[22];
  assign N157 = 1'b0 | retire_data_i[21];
  assign N158 = 1'b0 | retire_data_i[20];
  assign N159 = 1'b0 | retire_data_i[19];
  assign N160 = 1'b0 | retire_data_i[18];
  assign N161 = 1'b0 | retire_data_i[17];
  assign N162 = 1'b0 | retire_data_i[16];
  assign N163 = 1'b0 | retire_data_i[15];
  assign N164 = 1'b0 | retire_data_i[14];
  assign N165 = 1'b0 | retire_data_i[13];
  assign N166 = 1'b0 | retire_data_i[12];
  assign N167 = 1'b0 | retire_data_i[11];
  assign N168 = 1'b0 | retire_data_i[10];
  assign N169 = 1'b0 | retire_data_i[9];
  assign N170 = 1'b0 | retire_data_i[8];
  assign N171 = 1'b0 | retire_data_i[7];
  assign N172 = 1'b0 | retire_data_i[6];
  assign N173 = 1'b0 | retire_data_i[5];
  assign N174 = retire_instr_r[19] | retire_data_i[4];
  assign N175 = retire_instr_r[18] | retire_data_i[3];
  assign N176 = retire_instr_r[17] | retire_data_i[2];
  assign N177 = retire_instr_r[16] | retire_data_i[1];
  assign N178 = retire_instr_r[15] | retire_data_i[0];
  assign N179 = N443 & retire_data_i[63];
  assign N443 = ~1'b0;
  assign N180 = N444 & retire_data_i[62];
  assign N444 = ~1'b0;
  assign N181 = N445 & retire_data_i[61];
  assign N445 = ~1'b0;
  assign N182 = N446 & retire_data_i[60];
  assign N446 = ~1'b0;
  assign N183 = N447 & retire_data_i[59];
  assign N447 = ~1'b0;
  assign N184 = N448 & retire_data_i[58];
  assign N448 = ~1'b0;
  assign N185 = N449 & retire_data_i[57];
  assign N449 = ~1'b0;
  assign N186 = N450 & retire_data_i[56];
  assign N450 = ~1'b0;
  assign N187 = N451 & retire_data_i[55];
  assign N451 = ~1'b0;
  assign N188 = N452 & retire_data_i[54];
  assign N452 = ~1'b0;
  assign N189 = N453 & retire_data_i[53];
  assign N453 = ~1'b0;
  assign N190 = N454 & retire_data_i[52];
  assign N454 = ~1'b0;
  assign N191 = N455 & retire_data_i[51];
  assign N455 = ~1'b0;
  assign N192 = N456 & retire_data_i[50];
  assign N456 = ~1'b0;
  assign N193 = N457 & retire_data_i[49];
  assign N457 = ~1'b0;
  assign N194 = N458 & retire_data_i[48];
  assign N458 = ~1'b0;
  assign N195 = N459 & retire_data_i[47];
  assign N459 = ~1'b0;
  assign N196 = N460 & retire_data_i[46];
  assign N460 = ~1'b0;
  assign N197 = N461 & retire_data_i[45];
  assign N461 = ~1'b0;
  assign N198 = N462 & retire_data_i[44];
  assign N462 = ~1'b0;
  assign N199 = N463 & retire_data_i[43];
  assign N463 = ~1'b0;
  assign N200 = N464 & retire_data_i[42];
  assign N464 = ~1'b0;
  assign N201 = N465 & retire_data_i[41];
  assign N465 = ~1'b0;
  assign N202 = N466 & retire_data_i[40];
  assign N466 = ~1'b0;
  assign N203 = N467 & retire_data_i[39];
  assign N467 = ~1'b0;
  assign N204 = N468 & retire_data_i[38];
  assign N468 = ~1'b0;
  assign N205 = N469 & retire_data_i[37];
  assign N469 = ~1'b0;
  assign N206 = N470 & retire_data_i[36];
  assign N470 = ~1'b0;
  assign N207 = N471 & retire_data_i[35];
  assign N471 = ~1'b0;
  assign N208 = N472 & retire_data_i[34];
  assign N472 = ~1'b0;
  assign N209 = N473 & retire_data_i[33];
  assign N473 = ~1'b0;
  assign N210 = N474 & retire_data_i[32];
  assign N474 = ~1'b0;
  assign N211 = N475 & retire_data_i[31];
  assign N475 = ~1'b0;
  assign N212 = N476 & retire_data_i[30];
  assign N476 = ~1'b0;
  assign N213 = N477 & retire_data_i[29];
  assign N477 = ~1'b0;
  assign N214 = N478 & retire_data_i[28];
  assign N478 = ~1'b0;
  assign N215 = N479 & retire_data_i[27];
  assign N479 = ~1'b0;
  assign N216 = N480 & retire_data_i[26];
  assign N480 = ~1'b0;
  assign N217 = N481 & retire_data_i[25];
  assign N481 = ~1'b0;
  assign N218 = N482 & retire_data_i[24];
  assign N482 = ~1'b0;
  assign N219 = N483 & retire_data_i[23];
  assign N483 = ~1'b0;
  assign N220 = N484 & retire_data_i[22];
  assign N484 = ~1'b0;
  assign N221 = N485 & retire_data_i[21];
  assign N485 = ~1'b0;
  assign N222 = N486 & retire_data_i[20];
  assign N486 = ~1'b0;
  assign N223 = N487 & retire_data_i[19];
  assign N487 = ~1'b0;
  assign N224 = N488 & retire_data_i[18];
  assign N488 = ~1'b0;
  assign N225 = N489 & retire_data_i[17];
  assign N489 = ~1'b0;
  assign N226 = N490 & retire_data_i[16];
  assign N490 = ~1'b0;
  assign N227 = N491 & retire_data_i[15];
  assign N491 = ~1'b0;
  assign N228 = N492 & retire_data_i[14];
  assign N492 = ~1'b0;
  assign N229 = N493 & retire_data_i[13];
  assign N493 = ~1'b0;
  assign N230 = N494 & retire_data_i[12];
  assign N494 = ~1'b0;
  assign N231 = N495 & retire_data_i[11];
  assign N495 = ~1'b0;
  assign N232 = N496 & retire_data_i[10];
  assign N496 = ~1'b0;
  assign N233 = N497 & retire_data_i[9];
  assign N497 = ~1'b0;
  assign N234 = N498 & retire_data_i[8];
  assign N498 = ~1'b0;
  assign N235 = N499 & retire_data_i[7];
  assign N499 = ~1'b0;
  assign N236 = N500 & retire_data_i[6];
  assign N500 = ~1'b0;
  assign N237 = N501 & retire_data_i[5];
  assign N501 = ~1'b0;
  assign N238 = N502 & retire_data_i[4];
  assign N502 = ~retire_instr_r[19];
  assign N239 = N503 & retire_data_i[3];
  assign N503 = ~retire_instr_r[18];
  assign N240 = N504 & retire_data_i[2];
  assign N504 = ~retire_instr_r[17];
  assign N241 = N505 & retire_data_i[1];
  assign N505 = ~retire_instr_r[16];
  assign N242 = N506 & retire_data_i[0];
  assign N506 = ~retire_instr_r[15];
  assign N243 = retire_vaddr_r[63] | retire_data_i[63];
  assign N244 = retire_vaddr_r[62] | retire_data_i[62];
  assign N245 = retire_vaddr_r[61] | retire_data_i[61];
  assign N246 = retire_vaddr_r[60] | retire_data_i[60];
  assign N247 = retire_vaddr_r[59] | retire_data_i[59];
  assign N248 = retire_vaddr_r[58] | retire_data_i[58];
  assign N249 = retire_vaddr_r[57] | retire_data_i[57];
  assign N250 = retire_vaddr_r[56] | retire_data_i[56];
  assign N251 = retire_vaddr_r[55] | retire_data_i[55];
  assign N252 = retire_vaddr_r[54] | retire_data_i[54];
  assign N253 = retire_vaddr_r[53] | retire_data_i[53];
  assign N254 = retire_vaddr_r[52] | retire_data_i[52];
  assign N255 = retire_vaddr_r[51] | retire_data_i[51];
  assign N256 = retire_vaddr_r[50] | retire_data_i[50];
  assign N257 = retire_vaddr_r[49] | retire_data_i[49];
  assign N258 = retire_vaddr_r[48] | retire_data_i[48];
  assign N259 = retire_vaddr_r[47] | retire_data_i[47];
  assign N260 = retire_vaddr_r[46] | retire_data_i[46];
  assign N261 = retire_vaddr_r[45] | retire_data_i[45];
  assign N262 = retire_vaddr_r[44] | retire_data_i[44];
  assign N263 = retire_vaddr_r[43] | retire_data_i[43];
  assign N264 = retire_vaddr_r[42] | retire_data_i[42];
  assign N265 = retire_vaddr_r[41] | retire_data_i[41];
  assign N266 = retire_vaddr_r[40] | retire_data_i[40];
  assign N267 = retire_vaddr_r[39] | retire_data_i[39];
  assign N268 = retire_vaddr_r[38] | retire_data_i[38];
  assign N269 = retire_vaddr_r[37] | retire_data_i[37];
  assign N270 = retire_vaddr_r[36] | retire_data_i[36];
  assign N271 = retire_vaddr_r[35] | retire_data_i[35];
  assign N272 = retire_vaddr_r[34] | retire_data_i[34];
  assign N273 = retire_vaddr_r[33] | retire_data_i[33];
  assign N274 = retire_vaddr_r[32] | retire_data_i[32];
  assign N275 = retire_vaddr_r[31] | retire_data_i[31];
  assign N276 = retire_vaddr_r[30] | retire_data_i[30];
  assign N277 = retire_vaddr_r[29] | retire_data_i[29];
  assign N278 = retire_vaddr_r[28] | retire_data_i[28];
  assign N279 = retire_vaddr_r[27] | retire_data_i[27];
  assign N280 = retire_vaddr_r[26] | retire_data_i[26];
  assign N281 = retire_vaddr_r[25] | retire_data_i[25];
  assign N282 = retire_vaddr_r[24] | retire_data_i[24];
  assign N283 = retire_vaddr_r[23] | retire_data_i[23];
  assign N284 = retire_vaddr_r[22] | retire_data_i[22];
  assign N285 = retire_vaddr_r[21] | retire_data_i[21];
  assign N286 = retire_vaddr_r[20] | retire_data_i[20];
  assign N287 = retire_vaddr_r[19] | retire_data_i[19];
  assign N288 = retire_vaddr_r[18] | retire_data_i[18];
  assign N289 = retire_vaddr_r[17] | retire_data_i[17];
  assign N290 = retire_vaddr_r[16] | retire_data_i[16];
  assign N291 = retire_vaddr_r[15] | retire_data_i[15];
  assign N292 = retire_vaddr_r[14] | retire_data_i[14];
  assign N293 = retire_vaddr_r[13] | retire_data_i[13];
  assign N294 = retire_vaddr_r[12] | retire_data_i[12];
  assign N295 = retire_vaddr_r[11] | retire_data_i[11];
  assign N296 = retire_vaddr_r[10] | retire_data_i[10];
  assign N297 = retire_vaddr_r[9] | retire_data_i[9];
  assign N298 = retire_vaddr_r[8] | retire_data_i[8];
  assign N299 = retire_vaddr_r[7] | retire_data_i[7];
  assign N300 = retire_vaddr_r[6] | retire_data_i[6];
  assign N301 = retire_vaddr_r[5] | retire_data_i[5];
  assign N302 = retire_vaddr_r[4] | retire_data_i[4];
  assign N303 = retire_vaddr_r[3] | retire_data_i[3];
  assign N304 = retire_vaddr_r[2] | retire_data_i[2];
  assign N305 = retire_vaddr_r[1] | retire_data_i[1];
  assign N306 = retire_vaddr_r[0] | retire_data_i[0];
  assign N307 = N507 & retire_data_i[63];
  assign N507 = ~retire_vaddr_r[63];
  assign N308 = N508 & retire_data_i[62];
  assign N508 = ~retire_vaddr_r[62];
  assign N309 = N509 & retire_data_i[61];
  assign N509 = ~retire_vaddr_r[61];
  assign N310 = N510 & retire_data_i[60];
  assign N510 = ~retire_vaddr_r[60];
  assign N311 = N511 & retire_data_i[59];
  assign N511 = ~retire_vaddr_r[59];
  assign N312 = N512 & retire_data_i[58];
  assign N512 = ~retire_vaddr_r[58];
  assign N313 = N513 & retire_data_i[57];
  assign N513 = ~retire_vaddr_r[57];
  assign N314 = N514 & retire_data_i[56];
  assign N514 = ~retire_vaddr_r[56];
  assign N315 = N515 & retire_data_i[55];
  assign N515 = ~retire_vaddr_r[55];
  assign N316 = N516 & retire_data_i[54];
  assign N516 = ~retire_vaddr_r[54];
  assign N317 = N517 & retire_data_i[53];
  assign N517 = ~retire_vaddr_r[53];
  assign N318 = N518 & retire_data_i[52];
  assign N518 = ~retire_vaddr_r[52];
  assign N319 = N519 & retire_data_i[51];
  assign N519 = ~retire_vaddr_r[51];
  assign N320 = N520 & retire_data_i[50];
  assign N520 = ~retire_vaddr_r[50];
  assign N321 = N521 & retire_data_i[49];
  assign N521 = ~retire_vaddr_r[49];
  assign N322 = N522 & retire_data_i[48];
  assign N522 = ~retire_vaddr_r[48];
  assign N323 = N523 & retire_data_i[47];
  assign N523 = ~retire_vaddr_r[47];
  assign N324 = N524 & retire_data_i[46];
  assign N524 = ~retire_vaddr_r[46];
  assign N325 = N525 & retire_data_i[45];
  assign N525 = ~retire_vaddr_r[45];
  assign N326 = N526 & retire_data_i[44];
  assign N526 = ~retire_vaddr_r[44];
  assign N327 = N527 & retire_data_i[43];
  assign N527 = ~retire_vaddr_r[43];
  assign N328 = N528 & retire_data_i[42];
  assign N528 = ~retire_vaddr_r[42];
  assign N329 = N529 & retire_data_i[41];
  assign N529 = ~retire_vaddr_r[41];
  assign N330 = N530 & retire_data_i[40];
  assign N530 = ~retire_vaddr_r[40];
  assign N331 = N531 & retire_data_i[39];
  assign N531 = ~retire_vaddr_r[39];
  assign N332 = N532 & retire_data_i[38];
  assign N532 = ~retire_vaddr_r[38];
  assign N333 = N533 & retire_data_i[37];
  assign N533 = ~retire_vaddr_r[37];
  assign N334 = N534 & retire_data_i[36];
  assign N534 = ~retire_vaddr_r[36];
  assign N335 = N535 & retire_data_i[35];
  assign N535 = ~retire_vaddr_r[35];
  assign N336 = N536 & retire_data_i[34];
  assign N536 = ~retire_vaddr_r[34];
  assign N337 = N537 & retire_data_i[33];
  assign N537 = ~retire_vaddr_r[33];
  assign N338 = N538 & retire_data_i[32];
  assign N538 = ~retire_vaddr_r[32];
  assign N339 = N539 & retire_data_i[31];
  assign N539 = ~retire_vaddr_r[31];
  assign N340 = N540 & retire_data_i[30];
  assign N540 = ~retire_vaddr_r[30];
  assign N341 = N541 & retire_data_i[29];
  assign N541 = ~retire_vaddr_r[29];
  assign N342 = N542 & retire_data_i[28];
  assign N542 = ~retire_vaddr_r[28];
  assign N343 = N543 & retire_data_i[27];
  assign N543 = ~retire_vaddr_r[27];
  assign N344 = N544 & retire_data_i[26];
  assign N544 = ~retire_vaddr_r[26];
  assign N345 = N545 & retire_data_i[25];
  assign N545 = ~retire_vaddr_r[25];
  assign N346 = N546 & retire_data_i[24];
  assign N546 = ~retire_vaddr_r[24];
  assign N347 = N547 & retire_data_i[23];
  assign N547 = ~retire_vaddr_r[23];
  assign N348 = N548 & retire_data_i[22];
  assign N548 = ~retire_vaddr_r[22];
  assign N349 = N549 & retire_data_i[21];
  assign N549 = ~retire_vaddr_r[21];
  assign N350 = N550 & retire_data_i[20];
  assign N550 = ~retire_vaddr_r[20];
  assign N351 = N551 & retire_data_i[19];
  assign N551 = ~retire_vaddr_r[19];
  assign N352 = N552 & retire_data_i[18];
  assign N552 = ~retire_vaddr_r[18];
  assign N353 = N553 & retire_data_i[17];
  assign N553 = ~retire_vaddr_r[17];
  assign N354 = N554 & retire_data_i[16];
  assign N554 = ~retire_vaddr_r[16];
  assign N355 = N555 & retire_data_i[15];
  assign N555 = ~retire_vaddr_r[15];
  assign N356 = N556 & retire_data_i[14];
  assign N556 = ~retire_vaddr_r[14];
  assign N357 = N557 & retire_data_i[13];
  assign N557 = ~retire_vaddr_r[13];
  assign N358 = N558 & retire_data_i[12];
  assign N558 = ~retire_vaddr_r[12];
  assign N359 = N559 & retire_data_i[11];
  assign N559 = ~retire_vaddr_r[11];
  assign N360 = N560 & retire_data_i[10];
  assign N560 = ~retire_vaddr_r[10];
  assign N361 = N561 & retire_data_i[9];
  assign N561 = ~retire_vaddr_r[9];
  assign N362 = N562 & retire_data_i[8];
  assign N562 = ~retire_vaddr_r[8];
  assign N363 = N563 & retire_data_i[7];
  assign N563 = ~retire_vaddr_r[7];
  assign N364 = N564 & retire_data_i[6];
  assign N564 = ~retire_vaddr_r[6];
  assign N365 = N565 & retire_data_i[5];
  assign N565 = ~retire_vaddr_r[5];
  assign N366 = N566 & retire_data_i[4];
  assign N566 = ~retire_vaddr_r[4];
  assign N367 = N567 & retire_data_i[3];
  assign N567 = ~retire_vaddr_r[3];
  assign N368 = N568 & retire_data_i[2];
  assign N568 = ~retire_vaddr_r[2];
  assign N369 = N569 & retire_data_i[1];
  assign N569 = ~retire_vaddr_r[1];
  assign N370 = N570 & retire_data_i[0];
  assign N570 = ~retire_vaddr_r[0];
  assign retire_pkt_instret_ = N571 & N596;
  assign N571 = retire_v_i & retire_queue_v_i;
  assign N596 = ~N595;
  assign N595 = N594 | retire_exception_i[0];
  assign N594 = N593 | retire_exception_i[1];
  assign N593 = N592 | retire_exception_i[2];
  assign N592 = N591 | retire_exception_i[3];
  assign N591 = N590 | retire_exception_i[4];
  assign N590 = N589 | retire_exception_i[5];
  assign N589 = N588 | retire_exception_i[6];
  assign N588 = N587 | retire_exception_i[7];
  assign N587 = N586 | retire_exception_i[8];
  assign N586 = N585 | retire_exception_i[9];
  assign N585 = N584 | retire_exception_i[10];
  assign N584 = N583 | retire_exception_i[11];
  assign N583 = N582 | retire_exception_i[12];
  assign N582 = N581 | retire_exception_i[13];
  assign N581 = N580 | retire_exception_i[14];
  assign N580 = N579 | retire_exception_i[15];
  assign N579 = N578 | retire_exception_i[16];
  assign N578 = N577 | retire_exception_i[17];
  assign N577 = N576 | retire_exception_i[18];
  assign N576 = N575 | retire_exception_i[19];
  assign N575 = N574 | retire_exception_i[20];
  assign N574 = N573 | retire_exception_i[21];
  assign N573 = N572 | retire_exception_i[22];
  assign N572 = retire_exception_i[24] | retire_exception_i[23];
  assign iscore_li = N598 | N608;
  assign N598 = N597 & retire_iscore_r;
  assign N597 = ~retire_spec_w_r;
  assign N608 = N599 & N607;
  assign N599 = retire_spec_w_r & retire_iscore_r;
  assign N607 = N606 | retire_special_i[0];
  assign N606 = N605 | retire_special_i[1];
  assign N605 = N604 | retire_special_i[2];
  assign N604 = N603 | retire_special_i[3];
  assign N603 = N602 | retire_special_i[4];
  assign N602 = N601 | retire_special_i[5];
  assign N601 = N600 | retire_special_i[6];
  assign N600 = retire_special_i[8] | retire_special_i[7];
  assign fscore_li = N609 | N619;
  assign N609 = N597 & retire_fscore_r;
  assign N619 = N610 & N618;
  assign N610 = retire_spec_w_r & retire_fscore_r;
  assign N618 = N617 | retire_special_i[0];
  assign N617 = N616 | retire_special_i[1];
  assign N616 = N615 | retire_special_i[2];
  assign N615 = N614 | retire_special_i[3];
  assign N614 = N613 | retire_special_i[4];
  assign N613 = N612 | retire_special_i[5];
  assign N612 = N611 | retire_special_i[6];
  assign N611 = retire_special_i[8] | retire_special_i[7];
  assign N435 = ~retire_v_i;
  assign N436 = retire_v_i;
  assign N437 = ~retire_pkt_instret_;
  assign N438 = retire_pkt_instret_;
  assign N439 = ~retire_pkt_instret_;
  assign N440 = retire_pkt_instret_;
  assign N441 = ~retire_pkt_instret_;
  assign N442 = retire_pkt_instret_;

  always @(posedge clk_i) begin
    if(1'b1) begin
      retire_npc_r_38_sv2v_reg <= reservation_i[519];
      retire_npc_r_37_sv2v_reg <= reservation_i[518];
      retire_npc_r_36_sv2v_reg <= reservation_i[517];
      retire_npc_r_35_sv2v_reg <= reservation_i[516];
      retire_npc_r_34_sv2v_reg <= reservation_i[515];
      retire_npc_r_33_sv2v_reg <= reservation_i[514];
      retire_npc_r_32_sv2v_reg <= reservation_i[513];
      retire_npc_r_31_sv2v_reg <= reservation_i[512];
      retire_npc_r_30_sv2v_reg <= reservation_i[511];
      retire_npc_r_29_sv2v_reg <= reservation_i[510];
      retire_npc_r_28_sv2v_reg <= reservation_i[509];
      retire_npc_r_27_sv2v_reg <= reservation_i[508];
      retire_npc_r_26_sv2v_reg <= reservation_i[507];
      retire_npc_r_25_sv2v_reg <= reservation_i[506];
      retire_npc_r_24_sv2v_reg <= reservation_i[505];
      retire_npc_r_23_sv2v_reg <= reservation_i[504];
      retire_npc_r_22_sv2v_reg <= reservation_i[503];
      retire_npc_r_21_sv2v_reg <= reservation_i[502];
      retire_npc_r_20_sv2v_reg <= reservation_i[501];
      retire_npc_r_19_sv2v_reg <= reservation_i[500];
      retire_npc_r_18_sv2v_reg <= reservation_i[499];
      retire_npc_r_17_sv2v_reg <= reservation_i[498];
      retire_npc_r_16_sv2v_reg <= reservation_i[497];
      retire_npc_r_15_sv2v_reg <= reservation_i[496];
      retire_npc_r_14_sv2v_reg <= reservation_i[495];
      retire_npc_r_13_sv2v_reg <= reservation_i[494];
      retire_npc_r_12_sv2v_reg <= reservation_i[493];
      retire_npc_r_11_sv2v_reg <= reservation_i[492];
      retire_npc_r_10_sv2v_reg <= reservation_i[491];
      retire_npc_r_9_sv2v_reg <= reservation_i[490];
      retire_npc_r_8_sv2v_reg <= reservation_i[489];
      retire_npc_r_7_sv2v_reg <= reservation_i[488];
      retire_npc_r_6_sv2v_reg <= reservation_i[487];
      retire_npc_r_5_sv2v_reg <= reservation_i[486];
      retire_npc_r_4_sv2v_reg <= reservation_i[485];
      retire_npc_r_3_sv2v_reg <= reservation_i[484];
      retire_npc_r_2_sv2v_reg <= reservation_i[483];
      retire_npc_r_1_sv2v_reg <= reservation_i[482];
      retire_npc_r_0_sv2v_reg <= reservation_i[481];
      retire_nvaddr_r_63_sv2v_reg <= N79;
      retire_nvaddr_r_62_sv2v_reg <= N78;
      retire_nvaddr_r_61_sv2v_reg <= N77;
      retire_nvaddr_r_60_sv2v_reg <= N76;
      retire_nvaddr_r_59_sv2v_reg <= N75;
      retire_nvaddr_r_58_sv2v_reg <= N74;
      retire_nvaddr_r_57_sv2v_reg <= N73;
      retire_nvaddr_r_56_sv2v_reg <= N72;
      retire_nvaddr_r_55_sv2v_reg <= N71;
      retire_nvaddr_r_54_sv2v_reg <= N70;
      retire_nvaddr_r_53_sv2v_reg <= N69;
      retire_nvaddr_r_52_sv2v_reg <= N68;
      retire_nvaddr_r_51_sv2v_reg <= N67;
      retire_nvaddr_r_50_sv2v_reg <= N66;
      retire_nvaddr_r_49_sv2v_reg <= N65;
      retire_nvaddr_r_48_sv2v_reg <= N64;
      retire_nvaddr_r_47_sv2v_reg <= N63;
      retire_nvaddr_r_46_sv2v_reg <= N62;
      retire_nvaddr_r_45_sv2v_reg <= N61;
      retire_nvaddr_r_44_sv2v_reg <= N60;
      retire_nvaddr_r_43_sv2v_reg <= N59;
      retire_nvaddr_r_42_sv2v_reg <= N58;
      retire_nvaddr_r_41_sv2v_reg <= N57;
      retire_nvaddr_r_40_sv2v_reg <= N56;
      retire_nvaddr_r_39_sv2v_reg <= N55;
      retire_nvaddr_r_38_sv2v_reg <= N54;
      retire_nvaddr_r_37_sv2v_reg <= N53;
      retire_nvaddr_r_36_sv2v_reg <= N52;
      retire_nvaddr_r_35_sv2v_reg <= N51;
      retire_nvaddr_r_34_sv2v_reg <= N50;
      retire_nvaddr_r_33_sv2v_reg <= N49;
      retire_nvaddr_r_32_sv2v_reg <= N48;
      retire_nvaddr_r_31_sv2v_reg <= N47;
      retire_nvaddr_r_30_sv2v_reg <= N46;
      retire_nvaddr_r_29_sv2v_reg <= N45;
      retire_nvaddr_r_28_sv2v_reg <= N44;
      retire_nvaddr_r_27_sv2v_reg <= N43;
      retire_nvaddr_r_26_sv2v_reg <= N42;
      retire_nvaddr_r_25_sv2v_reg <= N41;
      retire_nvaddr_r_24_sv2v_reg <= N40;
      retire_nvaddr_r_23_sv2v_reg <= N39;
      retire_nvaddr_r_22_sv2v_reg <= N38;
      retire_nvaddr_r_21_sv2v_reg <= N37;
      retire_nvaddr_r_20_sv2v_reg <= N36;
      retire_nvaddr_r_19_sv2v_reg <= N35;
      retire_nvaddr_r_18_sv2v_reg <= N34;
      retire_nvaddr_r_17_sv2v_reg <= N33;
      retire_nvaddr_r_16_sv2v_reg <= N32;
      retire_nvaddr_r_15_sv2v_reg <= N31;
      retire_nvaddr_r_14_sv2v_reg <= N30;
      retire_nvaddr_r_13_sv2v_reg <= N29;
      retire_nvaddr_r_12_sv2v_reg <= N28;
      retire_nvaddr_r_11_sv2v_reg <= N27;
      retire_nvaddr_r_10_sv2v_reg <= N26;
      retire_nvaddr_r_9_sv2v_reg <= N25;
      retire_nvaddr_r_8_sv2v_reg <= N24;
      retire_nvaddr_r_7_sv2v_reg <= N23;
      retire_nvaddr_r_6_sv2v_reg <= N22;
      retire_nvaddr_r_5_sv2v_reg <= N21;
      retire_nvaddr_r_4_sv2v_reg <= N20;
      retire_nvaddr_r_3_sv2v_reg <= N19;
      retire_nvaddr_r_2_sv2v_reg <= N18;
      retire_nvaddr_r_1_sv2v_reg <= N17;
      retire_nvaddr_r_0_sv2v_reg <= N16;
      retire_vaddr_r_63_sv2v_reg <= retire_nvaddr_r[63];
      retire_vaddr_r_62_sv2v_reg <= retire_nvaddr_r[62];
      retire_vaddr_r_61_sv2v_reg <= retire_nvaddr_r[61];
      retire_vaddr_r_60_sv2v_reg <= retire_nvaddr_r[60];
      retire_vaddr_r_59_sv2v_reg <= retire_nvaddr_r[59];
      retire_vaddr_r_58_sv2v_reg <= retire_nvaddr_r[58];
      retire_vaddr_r_57_sv2v_reg <= retire_nvaddr_r[57];
      retire_vaddr_r_56_sv2v_reg <= retire_nvaddr_r[56];
      retire_vaddr_r_55_sv2v_reg <= retire_nvaddr_r[55];
      retire_vaddr_r_54_sv2v_reg <= retire_nvaddr_r[54];
      retire_vaddr_r_53_sv2v_reg <= retire_nvaddr_r[53];
      retire_vaddr_r_52_sv2v_reg <= retire_nvaddr_r[52];
      retire_vaddr_r_51_sv2v_reg <= retire_nvaddr_r[51];
      retire_vaddr_r_50_sv2v_reg <= retire_nvaddr_r[50];
      retire_vaddr_r_49_sv2v_reg <= retire_nvaddr_r[49];
      retire_vaddr_r_48_sv2v_reg <= retire_nvaddr_r[48];
      retire_vaddr_r_47_sv2v_reg <= retire_nvaddr_r[47];
      retire_vaddr_r_46_sv2v_reg <= retire_nvaddr_r[46];
      retire_vaddr_r_45_sv2v_reg <= retire_nvaddr_r[45];
      retire_vaddr_r_44_sv2v_reg <= retire_nvaddr_r[44];
      retire_vaddr_r_43_sv2v_reg <= retire_nvaddr_r[43];
      retire_vaddr_r_42_sv2v_reg <= retire_nvaddr_r[42];
      retire_vaddr_r_41_sv2v_reg <= retire_nvaddr_r[41];
      retire_vaddr_r_40_sv2v_reg <= retire_nvaddr_r[40];
      retire_vaddr_r_39_sv2v_reg <= retire_nvaddr_r[39];
      retire_vaddr_r_38_sv2v_reg <= retire_nvaddr_r[38];
      retire_vaddr_r_37_sv2v_reg <= retire_nvaddr_r[37];
      retire_vaddr_r_36_sv2v_reg <= retire_nvaddr_r[36];
      retire_vaddr_r_35_sv2v_reg <= retire_nvaddr_r[35];
      retire_vaddr_r_34_sv2v_reg <= retire_nvaddr_r[34];
      retire_vaddr_r_33_sv2v_reg <= retire_nvaddr_r[33];
      retire_vaddr_r_32_sv2v_reg <= retire_nvaddr_r[32];
      retire_vaddr_r_31_sv2v_reg <= retire_nvaddr_r[31];
      retire_vaddr_r_30_sv2v_reg <= retire_nvaddr_r[30];
      retire_vaddr_r_29_sv2v_reg <= retire_nvaddr_r[29];
      retire_vaddr_r_28_sv2v_reg <= retire_nvaddr_r[28];
      retire_vaddr_r_27_sv2v_reg <= retire_nvaddr_r[27];
      retire_vaddr_r_26_sv2v_reg <= retire_nvaddr_r[26];
      retire_vaddr_r_25_sv2v_reg <= retire_nvaddr_r[25];
      retire_vaddr_r_24_sv2v_reg <= retire_nvaddr_r[24];
      retire_vaddr_r_23_sv2v_reg <= retire_nvaddr_r[23];
      retire_vaddr_r_22_sv2v_reg <= retire_nvaddr_r[22];
      retire_vaddr_r_21_sv2v_reg <= retire_nvaddr_r[21];
      retire_vaddr_r_20_sv2v_reg <= retire_nvaddr_r[20];
      retire_vaddr_r_19_sv2v_reg <= retire_nvaddr_r[19];
      retire_vaddr_r_18_sv2v_reg <= retire_nvaddr_r[18];
      retire_vaddr_r_17_sv2v_reg <= retire_nvaddr_r[17];
      retire_vaddr_r_16_sv2v_reg <= retire_nvaddr_r[16];
      retire_vaddr_r_15_sv2v_reg <= retire_nvaddr_r[15];
      retire_vaddr_r_14_sv2v_reg <= retire_nvaddr_r[14];
      retire_vaddr_r_13_sv2v_reg <= retire_nvaddr_r[13];
      retire_vaddr_r_12_sv2v_reg <= retire_nvaddr_r[12];
      retire_vaddr_r_11_sv2v_reg <= retire_nvaddr_r[11];
      retire_vaddr_r_10_sv2v_reg <= retire_nvaddr_r[10];
      retire_vaddr_r_9_sv2v_reg <= retire_nvaddr_r[9];
      retire_vaddr_r_8_sv2v_reg <= retire_nvaddr_r[8];
      retire_vaddr_r_7_sv2v_reg <= retire_nvaddr_r[7];
      retire_vaddr_r_6_sv2v_reg <= retire_nvaddr_r[6];
      retire_vaddr_r_5_sv2v_reg <= retire_nvaddr_r[5];
      retire_vaddr_r_4_sv2v_reg <= retire_nvaddr_r[4];
      retire_vaddr_r_3_sv2v_reg <= retire_nvaddr_r[3];
      retire_vaddr_r_2_sv2v_reg <= retire_nvaddr_r[2];
      retire_vaddr_r_1_sv2v_reg <= retire_nvaddr_r[1];
      retire_vaddr_r_0_sv2v_reg <= retire_nvaddr_r[0];
      retire_nsize_r_1_sv2v_reg <= reservation_i[391];
      retire_nsize_r_0_sv2v_reg <= reservation_i[390];
      retire_size_r_1_sv2v_reg <= retire_nsize_r[1];
      retire_size_r_0_sv2v_reg <= retire_nsize_r[0];
      retire_ncount_r_2_sv2v_reg <= reservation_i[394];
      retire_ncount_r_1_sv2v_reg <= reservation_i[393];
      retire_ncount_r_0_sv2v_reg <= reservation_i[392];
      retire_count_r_2_sv2v_reg <= retire_ncount_r[2];
      retire_count_r_1_sv2v_reg <= retire_ncount_r[1];
      retire_count_r_0_sv2v_reg <= retire_ncount_r[0];
      retire_ninstr_r_31_sv2v_reg <= reservation_i[480];
      retire_ninstr_r_30_sv2v_reg <= reservation_i[479];
      retire_ninstr_r_29_sv2v_reg <= reservation_i[478];
      retire_ninstr_r_28_sv2v_reg <= reservation_i[477];
      retire_ninstr_r_27_sv2v_reg <= reservation_i[476];
      retire_ninstr_r_26_sv2v_reg <= reservation_i[475];
      retire_ninstr_r_25_sv2v_reg <= reservation_i[474];
      retire_ninstr_r_24_sv2v_reg <= reservation_i[473];
      retire_ninstr_r_23_sv2v_reg <= reservation_i[472];
      retire_ninstr_r_22_sv2v_reg <= reservation_i[471];
      retire_ninstr_r_21_sv2v_reg <= reservation_i[470];
      retire_ninstr_r_20_sv2v_reg <= reservation_i[469];
      retire_ninstr_r_19_sv2v_reg <= reservation_i[468];
      retire_ninstr_r_18_sv2v_reg <= reservation_i[467];
      retire_ninstr_r_17_sv2v_reg <= reservation_i[466];
      retire_ninstr_r_16_sv2v_reg <= reservation_i[465];
      retire_ninstr_r_15_sv2v_reg <= reservation_i[464];
      retire_ninstr_r_14_sv2v_reg <= reservation_i[463];
      retire_ninstr_r_13_sv2v_reg <= reservation_i[462];
      retire_ninstr_r_12_sv2v_reg <= reservation_i[461];
      retire_ninstr_r_11_sv2v_reg <= reservation_i[460];
      retire_ninstr_r_10_sv2v_reg <= reservation_i[459];
      retire_ninstr_r_9_sv2v_reg <= reservation_i[458];
      retire_ninstr_r_8_sv2v_reg <= reservation_i[457];
      retire_ninstr_r_7_sv2v_reg <= reservation_i[456];
      retire_ninstr_r_6_sv2v_reg <= reservation_i[455];
      retire_ninstr_r_5_sv2v_reg <= reservation_i[454];
      retire_ninstr_r_4_sv2v_reg <= reservation_i[453];
      retire_ninstr_r_3_sv2v_reg <= reservation_i[452];
      retire_ninstr_r_2_sv2v_reg <= reservation_i[451];
      retire_ninstr_r_1_sv2v_reg <= reservation_i[450];
      retire_ninstr_r_0_sv2v_reg <= reservation_i[449];
      retire_instr_r_31_sv2v_reg <= retire_ninstr_r[31];
      retire_instr_r_30_sv2v_reg <= retire_ninstr_r[30];
      retire_instr_r_29_sv2v_reg <= retire_ninstr_r[29];
      retire_instr_r_28_sv2v_reg <= retire_ninstr_r[28];
      retire_instr_r_27_sv2v_reg <= retire_ninstr_r[27];
      retire_instr_r_26_sv2v_reg <= retire_ninstr_r[26];
      retire_instr_r_25_sv2v_reg <= retire_ninstr_r[25];
      retire_instr_r_24_sv2v_reg <= retire_ninstr_r[24];
      retire_instr_r_23_sv2v_reg <= retire_ninstr_r[23];
      retire_instr_r_22_sv2v_reg <= retire_ninstr_r[22];
      retire_instr_r_21_sv2v_reg <= retire_ninstr_r[21];
      retire_instr_r_20_sv2v_reg <= retire_ninstr_r[20];
      retire_instr_r_19_sv2v_reg <= retire_ninstr_r[19];
      retire_instr_r_18_sv2v_reg <= retire_ninstr_r[18];
      retire_instr_r_17_sv2v_reg <= retire_ninstr_r[17];
      retire_instr_r_16_sv2v_reg <= retire_ninstr_r[16];
      retire_instr_r_15_sv2v_reg <= retire_ninstr_r[15];
      retire_instr_r_14_sv2v_reg <= retire_ninstr_r[14];
      retire_instr_r_13_sv2v_reg <= retire_ninstr_r[13];
      retire_instr_r_12_sv2v_reg <= retire_ninstr_r[12];
      retire_instr_r_11_sv2v_reg <= retire_ninstr_r[11];
      retire_instr_r_10_sv2v_reg <= retire_ninstr_r[10];
      retire_instr_r_9_sv2v_reg <= retire_ninstr_r[9];
      retire_instr_r_8_sv2v_reg <= retire_ninstr_r[8];
      retire_instr_r_7_sv2v_reg <= retire_ninstr_r[7];
      retire_instr_r_6_sv2v_reg <= retire_ninstr_r[6];
      retire_instr_r_5_sv2v_reg <= retire_ninstr_r[5];
      retire_instr_r_4_sv2v_reg <= retire_ninstr_r[4];
      retire_instr_r_3_sv2v_reg <= retire_ninstr_r[3];
      retire_instr_r_2_sv2v_reg <= retire_ninstr_r[2];
      retire_instr_r_1_sv2v_reg <= retire_ninstr_r[1];
      retire_instr_r_0_sv2v_reg <= retire_ninstr_r[0];
      retire_niscore_r_sv2v_reg <= N80;
      retire_iscore_r_sv2v_reg <= retire_niscore_r;
      retire_nfscore_r_sv2v_reg <= N81;
      retire_fscore_r_sv2v_reg <= retire_nfscore_r;
      retire_nspec_w_r_sv2v_reg <= N82;
      retire_spec_w_r_sv2v_reg <= retire_nspec_w_r;
    end 
  end


endmodule



module bsg_popcount_width_p4
(
  i,
  o
);

  input [3:0] i;
  output [2:0] o;
  wire [2:0] o;
  wire N0,N1;
  wire [1:0] \four.s0 ,\four.c0 ;
  assign \four.s0 [1] = i[3] ^ i[2];
  assign \four.s0 [0] = i[1] ^ i[0];
  assign \four.c0 [1] = i[3] & i[2];
  assign \four.c0 [0] = i[1] & i[0];
  assign o[0] = \four.s0 [1] ^ \four.s0 [0];
  assign o[1] = N0 | N1;
  assign N0 = \four.c0 [1] ^ \four.c0 [0];
  assign N1 = \four.s0 [1] & \four.s0 [0];
  assign o[2] = \four.c0 [1] & \four.c0 [0];

endmodule



module bsg_popcount_width_p8
(
  i,
  o
);

  input [7:0] i;
  output [3:0] o;
  wire [3:0] o;
  wire [2:0] \recurse.lo ,\recurse.hi ;

  bsg_popcount_width_p4
  \recurse.left 
  (
    .i(i[3:0]),
    .o(\recurse.lo )
  );


  bsg_popcount_width_p4
  \recurse.right 
  (
    .i(i[7:4]),
    .o(\recurse.hi )
  );

  assign o = \recurse.lo  + \recurse.hi ;

endmodule



module bsg_popcount_width_p16
(
  i,
  o
);

  input [15:0] i;
  output [4:0] o;
  wire [4:0] o;
  wire [3:0] \recurse.lo ,\recurse.hi ;

  bsg_popcount_width_p8
  \recurse.left 
  (
    .i(i[7:0]),
    .o(\recurse.lo )
  );


  bsg_popcount_width_p8
  \recurse.right 
  (
    .i(i[15:8]),
    .o(\recurse.hi )
  );

  assign o = \recurse.lo  + \recurse.hi ;

endmodule



module bsg_popcount_width_p32
(
  i,
  o
);

  input [31:0] i;
  output [5:0] o;
  wire [5:0] o;
  wire [4:0] \recurse.lo ,\recurse.hi ;

  bsg_popcount_width_p16
  \recurse.left 
  (
    .i(i[15:0]),
    .o(\recurse.lo )
  );


  bsg_popcount_width_p16
  \recurse.right 
  (
    .i(i[31:16]),
    .o(\recurse.hi )
  );

  assign o = \recurse.lo  + \recurse.hi ;

endmodule



module bsg_popcount_width_p64
(
  i,
  o
);

  input [63:0] i;
  output [6:0] o;
  wire [6:0] o;
  wire [5:0] \recurse.lo ,\recurse.hi ;

  bsg_popcount_width_p32
  \recurse.left 
  (
    .i(i[31:0]),
    .o(\recurse.lo )
  );


  bsg_popcount_width_p32
  \recurse.right 
  (
    .i(i[63:32]),
    .o(\recurse.hi )
  );

  assign o = \recurse.lo  + \recurse.hi ;

endmodule



module bsg_scan_width_p33_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [32:0] i;
  output [32:0] o;
  wire [32:0] o;
  wire t_5__32_,t_5__31_,t_5__30_,t_5__29_,t_5__28_,t_5__27_,t_5__26_,t_5__25_,
  t_5__24_,t_5__23_,t_5__22_,t_5__21_,t_5__20_,t_5__19_,t_5__18_,t_5__17_,t_5__16_,
  t_5__15_,t_5__14_,t_5__13_,t_5__12_,t_5__11_,t_5__10_,t_5__9_,t_5__8_,t_5__7_,t_5__6_,
  t_5__5_,t_5__4_,t_5__3_,t_5__2_,t_5__1_,t_5__0_,t_4__32_,t_4__31_,t_4__30_,
  t_4__29_,t_4__28_,t_4__27_,t_4__26_,t_4__25_,t_4__24_,t_4__23_,t_4__22_,t_4__21_,
  t_4__20_,t_4__19_,t_4__18_,t_4__17_,t_4__16_,t_4__15_,t_4__14_,t_4__13_,t_4__12_,
  t_4__11_,t_4__10_,t_4__9_,t_4__8_,t_4__7_,t_4__6_,t_4__5_,t_4__4_,t_4__3_,t_4__2_,
  t_4__1_,t_4__0_,t_3__32_,t_3__31_,t_3__30_,t_3__29_,t_3__28_,t_3__27_,t_3__26_,
  t_3__25_,t_3__24_,t_3__23_,t_3__22_,t_3__21_,t_3__20_,t_3__19_,t_3__18_,t_3__17_,
  t_3__16_,t_3__15_,t_3__14_,t_3__13_,t_3__12_,t_3__11_,t_3__10_,t_3__9_,t_3__8_,
  t_3__7_,t_3__6_,t_3__5_,t_3__4_,t_3__3_,t_3__2_,t_3__1_,t_3__0_,t_2__32_,t_2__31_,
  t_2__30_,t_2__29_,t_2__28_,t_2__27_,t_2__26_,t_2__25_,t_2__24_,t_2__23_,t_2__22_,
  t_2__21_,t_2__20_,t_2__19_,t_2__18_,t_2__17_,t_2__16_,t_2__15_,t_2__14_,
  t_2__13_,t_2__12_,t_2__11_,t_2__10_,t_2__9_,t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,
  t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__32_,t_1__31_,t_1__30_,t_1__29_,t_1__28_,
  t_1__27_,t_1__26_,t_1__25_,t_1__24_,t_1__23_,t_1__22_,t_1__21_,t_1__20_,t_1__19_,
  t_1__18_,t_1__17_,t_1__16_,t_1__15_,t_1__14_,t_1__13_,t_1__12_,t_1__11_,t_1__10_,
  t_1__9_,t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__32_ = i[0] | 1'b0;
  assign t_1__31_ = i[1] | i[0];
  assign t_1__30_ = i[2] | i[1];
  assign t_1__29_ = i[3] | i[2];
  assign t_1__28_ = i[4] | i[3];
  assign t_1__27_ = i[5] | i[4];
  assign t_1__26_ = i[6] | i[5];
  assign t_1__25_ = i[7] | i[6];
  assign t_1__24_ = i[8] | i[7];
  assign t_1__23_ = i[9] | i[8];
  assign t_1__22_ = i[10] | i[9];
  assign t_1__21_ = i[11] | i[10];
  assign t_1__20_ = i[12] | i[11];
  assign t_1__19_ = i[13] | i[12];
  assign t_1__18_ = i[14] | i[13];
  assign t_1__17_ = i[15] | i[14];
  assign t_1__16_ = i[16] | i[15];
  assign t_1__15_ = i[17] | i[16];
  assign t_1__14_ = i[18] | i[17];
  assign t_1__13_ = i[19] | i[18];
  assign t_1__12_ = i[20] | i[19];
  assign t_1__11_ = i[21] | i[20];
  assign t_1__10_ = i[22] | i[21];
  assign t_1__9_ = i[23] | i[22];
  assign t_1__8_ = i[24] | i[23];
  assign t_1__7_ = i[25] | i[24];
  assign t_1__6_ = i[26] | i[25];
  assign t_1__5_ = i[27] | i[26];
  assign t_1__4_ = i[28] | i[27];
  assign t_1__3_ = i[29] | i[28];
  assign t_1__2_ = i[30] | i[29];
  assign t_1__1_ = i[31] | i[30];
  assign t_1__0_ = i[32] | i[31];
  assign t_2__32_ = t_1__32_ | 1'b0;
  assign t_2__31_ = t_1__31_ | 1'b0;
  assign t_2__30_ = t_1__30_ | t_1__32_;
  assign t_2__29_ = t_1__29_ | t_1__31_;
  assign t_2__28_ = t_1__28_ | t_1__30_;
  assign t_2__27_ = t_1__27_ | t_1__29_;
  assign t_2__26_ = t_1__26_ | t_1__28_;
  assign t_2__25_ = t_1__25_ | t_1__27_;
  assign t_2__24_ = t_1__24_ | t_1__26_;
  assign t_2__23_ = t_1__23_ | t_1__25_;
  assign t_2__22_ = t_1__22_ | t_1__24_;
  assign t_2__21_ = t_1__21_ | t_1__23_;
  assign t_2__20_ = t_1__20_ | t_1__22_;
  assign t_2__19_ = t_1__19_ | t_1__21_;
  assign t_2__18_ = t_1__18_ | t_1__20_;
  assign t_2__17_ = t_1__17_ | t_1__19_;
  assign t_2__16_ = t_1__16_ | t_1__18_;
  assign t_2__15_ = t_1__15_ | t_1__17_;
  assign t_2__14_ = t_1__14_ | t_1__16_;
  assign t_2__13_ = t_1__13_ | t_1__15_;
  assign t_2__12_ = t_1__12_ | t_1__14_;
  assign t_2__11_ = t_1__11_ | t_1__13_;
  assign t_2__10_ = t_1__10_ | t_1__12_;
  assign t_2__9_ = t_1__9_ | t_1__11_;
  assign t_2__8_ = t_1__8_ | t_1__10_;
  assign t_2__7_ = t_1__7_ | t_1__9_;
  assign t_2__6_ = t_1__6_ | t_1__8_;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign t_3__32_ = t_2__32_ | 1'b0;
  assign t_3__31_ = t_2__31_ | 1'b0;
  assign t_3__30_ = t_2__30_ | 1'b0;
  assign t_3__29_ = t_2__29_ | 1'b0;
  assign t_3__28_ = t_2__28_ | t_2__32_;
  assign t_3__27_ = t_2__27_ | t_2__31_;
  assign t_3__26_ = t_2__26_ | t_2__30_;
  assign t_3__25_ = t_2__25_ | t_2__29_;
  assign t_3__24_ = t_2__24_ | t_2__28_;
  assign t_3__23_ = t_2__23_ | t_2__27_;
  assign t_3__22_ = t_2__22_ | t_2__26_;
  assign t_3__21_ = t_2__21_ | t_2__25_;
  assign t_3__20_ = t_2__20_ | t_2__24_;
  assign t_3__19_ = t_2__19_ | t_2__23_;
  assign t_3__18_ = t_2__18_ | t_2__22_;
  assign t_3__17_ = t_2__17_ | t_2__21_;
  assign t_3__16_ = t_2__16_ | t_2__20_;
  assign t_3__15_ = t_2__15_ | t_2__19_;
  assign t_3__14_ = t_2__14_ | t_2__18_;
  assign t_3__13_ = t_2__13_ | t_2__17_;
  assign t_3__12_ = t_2__12_ | t_2__16_;
  assign t_3__11_ = t_2__11_ | t_2__15_;
  assign t_3__10_ = t_2__10_ | t_2__14_;
  assign t_3__9_ = t_2__9_ | t_2__13_;
  assign t_3__8_ = t_2__8_ | t_2__12_;
  assign t_3__7_ = t_2__7_ | t_2__11_;
  assign t_3__6_ = t_2__6_ | t_2__10_;
  assign t_3__5_ = t_2__5_ | t_2__9_;
  assign t_3__4_ = t_2__4_ | t_2__8_;
  assign t_3__3_ = t_2__3_ | t_2__7_;
  assign t_3__2_ = t_2__2_ | t_2__6_;
  assign t_3__1_ = t_2__1_ | t_2__5_;
  assign t_3__0_ = t_2__0_ | t_2__4_;
  assign t_4__32_ = t_3__32_ | 1'b0;
  assign t_4__31_ = t_3__31_ | 1'b0;
  assign t_4__30_ = t_3__30_ | 1'b0;
  assign t_4__29_ = t_3__29_ | 1'b0;
  assign t_4__28_ = t_3__28_ | 1'b0;
  assign t_4__27_ = t_3__27_ | 1'b0;
  assign t_4__26_ = t_3__26_ | 1'b0;
  assign t_4__25_ = t_3__25_ | 1'b0;
  assign t_4__24_ = t_3__24_ | t_3__32_;
  assign t_4__23_ = t_3__23_ | t_3__31_;
  assign t_4__22_ = t_3__22_ | t_3__30_;
  assign t_4__21_ = t_3__21_ | t_3__29_;
  assign t_4__20_ = t_3__20_ | t_3__28_;
  assign t_4__19_ = t_3__19_ | t_3__27_;
  assign t_4__18_ = t_3__18_ | t_3__26_;
  assign t_4__17_ = t_3__17_ | t_3__25_;
  assign t_4__16_ = t_3__16_ | t_3__24_;
  assign t_4__15_ = t_3__15_ | t_3__23_;
  assign t_4__14_ = t_3__14_ | t_3__22_;
  assign t_4__13_ = t_3__13_ | t_3__21_;
  assign t_4__12_ = t_3__12_ | t_3__20_;
  assign t_4__11_ = t_3__11_ | t_3__19_;
  assign t_4__10_ = t_3__10_ | t_3__18_;
  assign t_4__9_ = t_3__9_ | t_3__17_;
  assign t_4__8_ = t_3__8_ | t_3__16_;
  assign t_4__7_ = t_3__7_ | t_3__15_;
  assign t_4__6_ = t_3__6_ | t_3__14_;
  assign t_4__5_ = t_3__5_ | t_3__13_;
  assign t_4__4_ = t_3__4_ | t_3__12_;
  assign t_4__3_ = t_3__3_ | t_3__11_;
  assign t_4__2_ = t_3__2_ | t_3__10_;
  assign t_4__1_ = t_3__1_ | t_3__9_;
  assign t_4__0_ = t_3__0_ | t_3__8_;
  assign t_5__32_ = t_4__32_ | 1'b0;
  assign t_5__31_ = t_4__31_ | 1'b0;
  assign t_5__30_ = t_4__30_ | 1'b0;
  assign t_5__29_ = t_4__29_ | 1'b0;
  assign t_5__28_ = t_4__28_ | 1'b0;
  assign t_5__27_ = t_4__27_ | 1'b0;
  assign t_5__26_ = t_4__26_ | 1'b0;
  assign t_5__25_ = t_4__25_ | 1'b0;
  assign t_5__24_ = t_4__24_ | 1'b0;
  assign t_5__23_ = t_4__23_ | 1'b0;
  assign t_5__22_ = t_4__22_ | 1'b0;
  assign t_5__21_ = t_4__21_ | 1'b0;
  assign t_5__20_ = t_4__20_ | 1'b0;
  assign t_5__19_ = t_4__19_ | 1'b0;
  assign t_5__18_ = t_4__18_ | 1'b0;
  assign t_5__17_ = t_4__17_ | 1'b0;
  assign t_5__16_ = t_4__16_ | t_4__32_;
  assign t_5__15_ = t_4__15_ | t_4__31_;
  assign t_5__14_ = t_4__14_ | t_4__30_;
  assign t_5__13_ = t_4__13_ | t_4__29_;
  assign t_5__12_ = t_4__12_ | t_4__28_;
  assign t_5__11_ = t_4__11_ | t_4__27_;
  assign t_5__10_ = t_4__10_ | t_4__26_;
  assign t_5__9_ = t_4__9_ | t_4__25_;
  assign t_5__8_ = t_4__8_ | t_4__24_;
  assign t_5__7_ = t_4__7_ | t_4__23_;
  assign t_5__6_ = t_4__6_ | t_4__22_;
  assign t_5__5_ = t_4__5_ | t_4__21_;
  assign t_5__4_ = t_4__4_ | t_4__20_;
  assign t_5__3_ = t_4__3_ | t_4__19_;
  assign t_5__2_ = t_4__2_ | t_4__18_;
  assign t_5__1_ = t_4__1_ | t_4__17_;
  assign t_5__0_ = t_4__0_ | t_4__16_;
  assign o[0] = t_5__32_ | 1'b0;
  assign o[1] = t_5__31_ | 1'b0;
  assign o[2] = t_5__30_ | 1'b0;
  assign o[3] = t_5__29_ | 1'b0;
  assign o[4] = t_5__28_ | 1'b0;
  assign o[5] = t_5__27_ | 1'b0;
  assign o[6] = t_5__26_ | 1'b0;
  assign o[7] = t_5__25_ | 1'b0;
  assign o[8] = t_5__24_ | 1'b0;
  assign o[9] = t_5__23_ | 1'b0;
  assign o[10] = t_5__22_ | 1'b0;
  assign o[11] = t_5__21_ | 1'b0;
  assign o[12] = t_5__20_ | 1'b0;
  assign o[13] = t_5__19_ | 1'b0;
  assign o[14] = t_5__18_ | 1'b0;
  assign o[15] = t_5__17_ | 1'b0;
  assign o[16] = t_5__16_ | 1'b0;
  assign o[17] = t_5__15_ | 1'b0;
  assign o[18] = t_5__14_ | 1'b0;
  assign o[19] = t_5__13_ | 1'b0;
  assign o[20] = t_5__12_ | 1'b0;
  assign o[21] = t_5__11_ | 1'b0;
  assign o[22] = t_5__10_ | 1'b0;
  assign o[23] = t_5__9_ | 1'b0;
  assign o[24] = t_5__8_ | 1'b0;
  assign o[25] = t_5__7_ | 1'b0;
  assign o[26] = t_5__6_ | 1'b0;
  assign o[27] = t_5__5_ | 1'b0;
  assign o[28] = t_5__4_ | 1'b0;
  assign o[29] = t_5__3_ | 1'b0;
  assign o[30] = t_5__2_ | 1'b0;
  assign o[31] = t_5__1_ | 1'b0;
  assign o[32] = t_5__0_ | t_5__32_;

endmodule



module bsg_priority_encode_one_hot_out_width_p33_lo_to_hi_p1
(
  i,
  o,
  v_o
);

  input [32:0] i;
  output [32:0] o;
  output v_o;
  wire [32:0] o;
  wire v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31;
  wire [31:1] scan_lo;

  bsg_scan_width_p33_or_p1_lo_to_hi_p1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, scan_lo, o[0:0] })
  );

  assign o[32] = v_o & N0;
  assign N0 = ~scan_lo[31];
  assign o[31] = scan_lo[31] & N1;
  assign N1 = ~scan_lo[30];
  assign o[30] = scan_lo[30] & N2;
  assign N2 = ~scan_lo[29];
  assign o[29] = scan_lo[29] & N3;
  assign N3 = ~scan_lo[28];
  assign o[28] = scan_lo[28] & N4;
  assign N4 = ~scan_lo[27];
  assign o[27] = scan_lo[27] & N5;
  assign N5 = ~scan_lo[26];
  assign o[26] = scan_lo[26] & N6;
  assign N6 = ~scan_lo[25];
  assign o[25] = scan_lo[25] & N7;
  assign N7 = ~scan_lo[24];
  assign o[24] = scan_lo[24] & N8;
  assign N8 = ~scan_lo[23];
  assign o[23] = scan_lo[23] & N9;
  assign N9 = ~scan_lo[22];
  assign o[22] = scan_lo[22] & N10;
  assign N10 = ~scan_lo[21];
  assign o[21] = scan_lo[21] & N11;
  assign N11 = ~scan_lo[20];
  assign o[20] = scan_lo[20] & N12;
  assign N12 = ~scan_lo[19];
  assign o[19] = scan_lo[19] & N13;
  assign N13 = ~scan_lo[18];
  assign o[18] = scan_lo[18] & N14;
  assign N14 = ~scan_lo[17];
  assign o[17] = scan_lo[17] & N15;
  assign N15 = ~scan_lo[16];
  assign o[16] = scan_lo[16] & N16;
  assign N16 = ~scan_lo[15];
  assign o[15] = scan_lo[15] & N17;
  assign N17 = ~scan_lo[14];
  assign o[14] = scan_lo[14] & N18;
  assign N18 = ~scan_lo[13];
  assign o[13] = scan_lo[13] & N19;
  assign N19 = ~scan_lo[12];
  assign o[12] = scan_lo[12] & N20;
  assign N20 = ~scan_lo[11];
  assign o[11] = scan_lo[11] & N21;
  assign N21 = ~scan_lo[10];
  assign o[10] = scan_lo[10] & N22;
  assign N22 = ~scan_lo[9];
  assign o[9] = scan_lo[9] & N23;
  assign N23 = ~scan_lo[8];
  assign o[8] = scan_lo[8] & N24;
  assign N24 = ~scan_lo[7];
  assign o[7] = scan_lo[7] & N25;
  assign N25 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N26;
  assign N26 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N27;
  assign N27 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N28;
  assign N28 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N29;
  assign N29 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N30;
  assign N30 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N31;
  assign N31 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p33_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [32:0] i;
  output [5:0] addr_o;
  output v_o;
  wire [5:0] addr_o;
  wire v_o,v_5__0_,v_4__48_,v_4__32_,v_4__16_,v_4__0_,v_3__56_,v_3__48_,v_3__40_,
  v_3__32_,v_3__24_,v_3__16_,v_3__8_,v_3__0_,v_2__60_,v_2__56_,v_2__52_,v_2__48_,
  v_2__44_,v_2__40_,v_2__36_,v_2__32_,v_2__28_,v_2__24_,v_2__20_,v_2__16_,v_2__12_,
  v_2__8_,v_2__4_,v_2__0_,v_1__62_,v_1__60_,v_1__58_,v_1__56_,v_1__54_,v_1__52_,
  v_1__50_,v_1__48_,v_1__46_,v_1__44_,v_1__42_,v_1__40_,v_1__38_,v_1__36_,v_1__34_,
  v_1__32_,v_1__30_,v_1__28_,v_1__26_,v_1__24_,v_1__22_,v_1__20_,v_1__18_,v_1__16_,
  v_1__14_,v_1__12_,v_1__10_,v_1__8_,v_1__6_,v_1__4_,v_1__2_,v_1__0_,addr_5__35_,
  addr_5__34_,addr_5__33_,addr_5__32_,addr_5__3_,addr_5__2_,addr_5__1_,addr_5__0_,
  addr_4__50_,addr_4__49_,addr_4__48_,addr_4__34_,addr_4__33_,addr_4__32_,addr_4__18_,
  addr_4__17_,addr_4__16_,addr_4__2_,addr_4__1_,addr_4__0_,addr_3__57_,addr_3__56_,
  addr_3__49_,addr_3__48_,addr_3__41_,addr_3__40_,addr_3__33_,addr_3__32_,
  addr_3__25_,addr_3__24_,addr_3__17_,addr_3__16_,addr_3__9_,addr_3__8_,addr_3__1_,
  addr_3__0_,addr_2__60_,addr_2__56_,addr_2__52_,addr_2__48_,addr_2__44_,addr_2__40_,
  addr_2__36_,addr_2__32_,addr_2__28_,addr_2__24_,addr_2__20_,addr_2__16_,addr_2__12_,
  addr_2__8_,addr_2__4_,addr_2__0_;
  assign v_1__0_ = i[1] | i[0];
  assign v_1__2_ = i[3] | i[2];
  assign v_1__4_ = i[5] | i[4];
  assign v_1__6_ = i[7] | i[6];
  assign v_1__8_ = i[9] | i[8];
  assign v_1__10_ = i[11] | i[10];
  assign v_1__12_ = i[13] | i[12];
  assign v_1__14_ = i[15] | i[14];
  assign v_1__16_ = i[17] | i[16];
  assign v_1__18_ = i[19] | i[18];
  assign v_1__20_ = i[21] | i[20];
  assign v_1__22_ = i[23] | i[22];
  assign v_1__24_ = i[25] | i[24];
  assign v_1__26_ = i[27] | i[26];
  assign v_1__28_ = i[29] | i[28];
  assign v_1__30_ = i[31] | i[30];
  assign v_1__32_ = 1'b0 | i[32];
  assign v_1__34_ = 1'b0 | 1'b0;
  assign v_1__36_ = 1'b0 | 1'b0;
  assign v_1__38_ = 1'b0 | 1'b0;
  assign v_1__40_ = 1'b0 | 1'b0;
  assign v_1__42_ = 1'b0 | 1'b0;
  assign v_1__44_ = 1'b0 | 1'b0;
  assign v_1__46_ = 1'b0 | 1'b0;
  assign v_1__48_ = 1'b0 | 1'b0;
  assign v_1__50_ = 1'b0 | 1'b0;
  assign v_1__52_ = 1'b0 | 1'b0;
  assign v_1__54_ = 1'b0 | 1'b0;
  assign v_1__56_ = 1'b0 | 1'b0;
  assign v_1__58_ = 1'b0 | 1'b0;
  assign v_1__60_ = 1'b0 | 1'b0;
  assign v_1__62_ = 1'b0 | 1'b0;
  assign v_2__0_ = v_1__2_ | v_1__0_;
  assign addr_2__0_ = i[1] | i[3];
  assign v_2__4_ = v_1__6_ | v_1__4_;
  assign addr_2__4_ = i[5] | i[7];
  assign v_2__8_ = v_1__10_ | v_1__8_;
  assign addr_2__8_ = i[9] | i[11];
  assign v_2__12_ = v_1__14_ | v_1__12_;
  assign addr_2__12_ = i[13] | i[15];
  assign v_2__16_ = v_1__18_ | v_1__16_;
  assign addr_2__16_ = i[17] | i[19];
  assign v_2__20_ = v_1__22_ | v_1__20_;
  assign addr_2__20_ = i[21] | i[23];
  assign v_2__24_ = v_1__26_ | v_1__24_;
  assign addr_2__24_ = i[25] | i[27];
  assign v_2__28_ = v_1__30_ | v_1__28_;
  assign addr_2__28_ = i[29] | i[31];
  assign v_2__32_ = v_1__34_ | v_1__32_;
  assign addr_2__32_ = 1'b0 | 1'b0;
  assign v_2__36_ = v_1__38_ | v_1__36_;
  assign addr_2__36_ = 1'b0 | 1'b0;
  assign v_2__40_ = v_1__42_ | v_1__40_;
  assign addr_2__40_ = 1'b0 | 1'b0;
  assign v_2__44_ = v_1__46_ | v_1__44_;
  assign addr_2__44_ = 1'b0 | 1'b0;
  assign v_2__48_ = v_1__50_ | v_1__48_;
  assign addr_2__48_ = 1'b0 | 1'b0;
  assign v_2__52_ = v_1__54_ | v_1__52_;
  assign addr_2__52_ = 1'b0 | 1'b0;
  assign v_2__56_ = v_1__58_ | v_1__56_;
  assign addr_2__56_ = 1'b0 | 1'b0;
  assign v_2__60_ = v_1__62_ | v_1__60_;
  assign addr_2__60_ = 1'b0 | 1'b0;
  assign v_3__0_ = v_2__4_ | v_2__0_;
  assign addr_3__1_ = v_1__2_ | v_1__6_;
  assign addr_3__0_ = addr_2__0_ | addr_2__4_;
  assign v_3__8_ = v_2__12_ | v_2__8_;
  assign addr_3__9_ = v_1__10_ | v_1__14_;
  assign addr_3__8_ = addr_2__8_ | addr_2__12_;
  assign v_3__16_ = v_2__20_ | v_2__16_;
  assign addr_3__17_ = v_1__18_ | v_1__22_;
  assign addr_3__16_ = addr_2__16_ | addr_2__20_;
  assign v_3__24_ = v_2__28_ | v_2__24_;
  assign addr_3__25_ = v_1__26_ | v_1__30_;
  assign addr_3__24_ = addr_2__24_ | addr_2__28_;
  assign v_3__32_ = v_2__36_ | v_2__32_;
  assign addr_3__33_ = v_1__34_ | v_1__38_;
  assign addr_3__32_ = addr_2__32_ | addr_2__36_;
  assign v_3__40_ = v_2__44_ | v_2__40_;
  assign addr_3__41_ = v_1__42_ | v_1__46_;
  assign addr_3__40_ = addr_2__40_ | addr_2__44_;
  assign v_3__48_ = v_2__52_ | v_2__48_;
  assign addr_3__49_ = v_1__50_ | v_1__54_;
  assign addr_3__48_ = addr_2__48_ | addr_2__52_;
  assign v_3__56_ = v_2__60_ | v_2__56_;
  assign addr_3__57_ = v_1__58_ | v_1__62_;
  assign addr_3__56_ = addr_2__56_ | addr_2__60_;
  assign v_4__0_ = v_3__8_ | v_3__0_;
  assign addr_4__2_ = v_2__4_ | v_2__12_;
  assign addr_4__1_ = addr_3__1_ | addr_3__9_;
  assign addr_4__0_ = addr_3__0_ | addr_3__8_;
  assign v_4__16_ = v_3__24_ | v_3__16_;
  assign addr_4__18_ = v_2__20_ | v_2__28_;
  assign addr_4__17_ = addr_3__17_ | addr_3__25_;
  assign addr_4__16_ = addr_3__16_ | addr_3__24_;
  assign v_4__32_ = v_3__40_ | v_3__32_;
  assign addr_4__34_ = v_2__36_ | v_2__44_;
  assign addr_4__33_ = addr_3__33_ | addr_3__41_;
  assign addr_4__32_ = addr_3__32_ | addr_3__40_;
  assign v_4__48_ = v_3__56_ | v_3__48_;
  assign addr_4__50_ = v_2__52_ | v_2__60_;
  assign addr_4__49_ = addr_3__49_ | addr_3__57_;
  assign addr_4__48_ = addr_3__48_ | addr_3__56_;
  assign v_5__0_ = v_4__16_ | v_4__0_;
  assign addr_5__3_ = v_3__8_ | v_3__24_;
  assign addr_5__2_ = addr_4__2_ | addr_4__18_;
  assign addr_5__1_ = addr_4__1_ | addr_4__17_;
  assign addr_5__0_ = addr_4__0_ | addr_4__16_;
  assign addr_o[5] = v_4__48_ | v_4__32_;
  assign addr_5__35_ = v_3__40_ | v_3__56_;
  assign addr_5__34_ = addr_4__34_ | addr_4__50_;
  assign addr_5__33_ = addr_4__33_ | addr_4__49_;
  assign addr_5__32_ = addr_4__32_ | addr_4__48_;
  assign v_o = addr_o[5] | v_5__0_;
  assign addr_o[4] = v_4__16_ | v_4__48_;
  assign addr_o[3] = addr_5__3_ | addr_5__35_;
  assign addr_o[2] = addr_5__2_ | addr_5__34_;
  assign addr_o[1] = addr_5__1_ | addr_5__33_;
  assign addr_o[0] = addr_5__0_ | addr_5__32_;

endmodule



module bsg_priority_encode_width_p33_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [32:0] i;
  output [5:0] addr_o;
  output v_o;
  wire [5:0] addr_o;
  wire v_o;
  wire [32:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p33_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_width_p33_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o)
  );


endmodule



module bsg_counting_leading_zeros_width_p32
(
  a_i,
  num_zero_o
);

  input [31:0] a_i;
  output [5:0] num_zero_o;
  wire [5:0] num_zero_o;

  bsg_priority_encode_width_p33_lo_to_hi_p1
  pe0
  (
    .i({ 1'b1, a_i[0:0], a_i[1:1], a_i[2:2], a_i[3:3], a_i[4:4], a_i[5:5], a_i[6:6], a_i[7:7], a_i[8:8], a_i[9:9], a_i[10:10], a_i[11:11], a_i[12:12], a_i[13:13], a_i[14:14], a_i[15:15], a_i[16:16], a_i[17:17], a_i[18:18], a_i[19:19], a_i[20:20], a_i[21:21], a_i[22:22], a_i[23:23], a_i[24:24], a_i[25:25], a_i[26:26], a_i[27:27], a_i[28:28], a_i[29:29], a_i[30:30], a_i[31:31] }),
    .addr_o(num_zero_o)
  );


endmodule



module bp_be_int_box_00
(
  raw_i,
  tag_i,
  unsigned_i,
  reg_o
);

  input [63:0] raw_i;
  input [1:0] tag_i;
  output [65:0] reg_o;
  input unsigned_i;
  wire [65:0] reg_o;
  wire N0,N1,N2,N3,N4,reg_o_65_,reg_o_64_,reg_o_62_,reg_o_61_,reg_o_60_,reg_o_59_,
  reg_o_58_,reg_o_57_,reg_o_56_,reg_o_55_,reg_o_54_,reg_o_53_,reg_o_52_,reg_o_51_,
  reg_o_50_,reg_o_49_,reg_o_48_,reg_o_47_,reg_o_46_,reg_o_45_,reg_o_44_,reg_o_43_,
  reg_o_42_,reg_o_41_,reg_o_40_,reg_o_39_,reg_o_38_,reg_o_37_,reg_o_36_,reg_o_35_,
  reg_o_34_,reg_o_33_,reg_o_32_,reg_o_31_,reg_o_30_,reg_o_29_,reg_o_28_,reg_o_27_,
  reg_o_26_,reg_o_25_,reg_o_24_,reg_o_23_,reg_o_22_,reg_o_21_,reg_o_20_,reg_o_19_,
  reg_o_18_,reg_o_17_,reg_o_16_,reg_o_15_,reg_o_14_,reg_o_13_,reg_o_12_,reg_o_11_,
  reg_o_10_,reg_o_9_,reg_o_8_,reg_o_7_,reg_o_6_,reg_o_5_,reg_o_4_,reg_o_3_,reg_o_2_,
  reg_o_1_,reg_o_0_,N5,N6,N7,N8,N9,N10,N11,N12,sig,N13,N14,N15,N16;
  assign reg_o_65_ = tag_i[1];
  assign reg_o[65] = reg_o_65_;
  assign reg_o_64_ = tag_i[0];
  assign reg_o[64] = reg_o_64_;
  assign reg_o_62_ = raw_i[62];
  assign reg_o[62] = reg_o_62_;
  assign reg_o_61_ = raw_i[61];
  assign reg_o[61] = reg_o_61_;
  assign reg_o_60_ = raw_i[60];
  assign reg_o[60] = reg_o_60_;
  assign reg_o_59_ = raw_i[59];
  assign reg_o[59] = reg_o_59_;
  assign reg_o_58_ = raw_i[58];
  assign reg_o[58] = reg_o_58_;
  assign reg_o_57_ = raw_i[57];
  assign reg_o[57] = reg_o_57_;
  assign reg_o_56_ = raw_i[56];
  assign reg_o[56] = reg_o_56_;
  assign reg_o_55_ = raw_i[55];
  assign reg_o[55] = reg_o_55_;
  assign reg_o_54_ = raw_i[54];
  assign reg_o[54] = reg_o_54_;
  assign reg_o_53_ = raw_i[53];
  assign reg_o[53] = reg_o_53_;
  assign reg_o_52_ = raw_i[52];
  assign reg_o[52] = reg_o_52_;
  assign reg_o_51_ = raw_i[51];
  assign reg_o[51] = reg_o_51_;
  assign reg_o_50_ = raw_i[50];
  assign reg_o[50] = reg_o_50_;
  assign reg_o_49_ = raw_i[49];
  assign reg_o[49] = reg_o_49_;
  assign reg_o_48_ = raw_i[48];
  assign reg_o[48] = reg_o_48_;
  assign reg_o_47_ = raw_i[47];
  assign reg_o[47] = reg_o_47_;
  assign reg_o_46_ = raw_i[46];
  assign reg_o[46] = reg_o_46_;
  assign reg_o_45_ = raw_i[45];
  assign reg_o[45] = reg_o_45_;
  assign reg_o_44_ = raw_i[44];
  assign reg_o[44] = reg_o_44_;
  assign reg_o_43_ = raw_i[43];
  assign reg_o[43] = reg_o_43_;
  assign reg_o_42_ = raw_i[42];
  assign reg_o[42] = reg_o_42_;
  assign reg_o_41_ = raw_i[41];
  assign reg_o[41] = reg_o_41_;
  assign reg_o_40_ = raw_i[40];
  assign reg_o[40] = reg_o_40_;
  assign reg_o_39_ = raw_i[39];
  assign reg_o[39] = reg_o_39_;
  assign reg_o_38_ = raw_i[38];
  assign reg_o[38] = reg_o_38_;
  assign reg_o_37_ = raw_i[37];
  assign reg_o[37] = reg_o_37_;
  assign reg_o_36_ = raw_i[36];
  assign reg_o[36] = reg_o_36_;
  assign reg_o_35_ = raw_i[35];
  assign reg_o[35] = reg_o_35_;
  assign reg_o_34_ = raw_i[34];
  assign reg_o[34] = reg_o_34_;
  assign reg_o_33_ = raw_i[33];
  assign reg_o[33] = reg_o_33_;
  assign reg_o_32_ = raw_i[32];
  assign reg_o[32] = reg_o_32_;
  assign reg_o_31_ = raw_i[31];
  assign reg_o[31] = reg_o_31_;
  assign reg_o_30_ = raw_i[30];
  assign reg_o[30] = reg_o_30_;
  assign reg_o_29_ = raw_i[29];
  assign reg_o[29] = reg_o_29_;
  assign reg_o_28_ = raw_i[28];
  assign reg_o[28] = reg_o_28_;
  assign reg_o_27_ = raw_i[27];
  assign reg_o[27] = reg_o_27_;
  assign reg_o_26_ = raw_i[26];
  assign reg_o[26] = reg_o_26_;
  assign reg_o_25_ = raw_i[25];
  assign reg_o[25] = reg_o_25_;
  assign reg_o_24_ = raw_i[24];
  assign reg_o[24] = reg_o_24_;
  assign reg_o_23_ = raw_i[23];
  assign reg_o[23] = reg_o_23_;
  assign reg_o_22_ = raw_i[22];
  assign reg_o[22] = reg_o_22_;
  assign reg_o_21_ = raw_i[21];
  assign reg_o[21] = reg_o_21_;
  assign reg_o_20_ = raw_i[20];
  assign reg_o[20] = reg_o_20_;
  assign reg_o_19_ = raw_i[19];
  assign reg_o[19] = reg_o_19_;
  assign reg_o_18_ = raw_i[18];
  assign reg_o[18] = reg_o_18_;
  assign reg_o_17_ = raw_i[17];
  assign reg_o[17] = reg_o_17_;
  assign reg_o_16_ = raw_i[16];
  assign reg_o[16] = reg_o_16_;
  assign reg_o_15_ = raw_i[15];
  assign reg_o[15] = reg_o_15_;
  assign reg_o_14_ = raw_i[14];
  assign reg_o[14] = reg_o_14_;
  assign reg_o_13_ = raw_i[13];
  assign reg_o[13] = reg_o_13_;
  assign reg_o_12_ = raw_i[12];
  assign reg_o[12] = reg_o_12_;
  assign reg_o_11_ = raw_i[11];
  assign reg_o[11] = reg_o_11_;
  assign reg_o_10_ = raw_i[10];
  assign reg_o[10] = reg_o_10_;
  assign reg_o_9_ = raw_i[9];
  assign reg_o[9] = reg_o_9_;
  assign reg_o_8_ = raw_i[8];
  assign reg_o[8] = reg_o_8_;
  assign reg_o_7_ = raw_i[7];
  assign reg_o[7] = reg_o_7_;
  assign reg_o_6_ = raw_i[6];
  assign reg_o[6] = reg_o_6_;
  assign reg_o_5_ = raw_i[5];
  assign reg_o[5] = reg_o_5_;
  assign reg_o_4_ = raw_i[4];
  assign reg_o[4] = reg_o_4_;
  assign reg_o_3_ = raw_i[3];
  assign reg_o[3] = reg_o_3_;
  assign reg_o_2_ = raw_i[2];
  assign reg_o[2] = reg_o_2_;
  assign reg_o_1_ = raw_i[1];
  assign reg_o[1] = reg_o_1_;
  assign reg_o_0_ = raw_i[0];
  assign reg_o[0] = reg_o_0_;
  assign N5 = reg_o_65_ & reg_o_64_;
  assign N7 = N6 | reg_o_64_;
  assign N10 = reg_o_65_ | N9;
  assign N12 = N6 & N9;
  assign N15 = reg_o_64_ | reg_o_65_;
  assign sig = (N0)? reg_o_7_ : 
               (N1)? reg_o_15_ : 
               (N2)? reg_o_31_ : 
               (N3)? raw_i[63] : 1'b0;
  assign N0 = N5;
  assign N1 = N8;
  assign N2 = N11;
  assign N3 = N12;
  assign reg_o[63] = (N4)? N14 : 
                     (N13)? raw_i[63] : 1'b0;
  assign N4 = N15;
  assign N6 = ~reg_o_65_;
  assign N8 = ~N7;
  assign N9 = ~reg_o_64_;
  assign N11 = ~N10;
  assign N13 = ~N15;
  assign N14 = sig & N16;
  assign N16 = ~unsigned_i;

endmodule



module bp_be_pipe_int_00
(
  clk_i,
  reset_i,
  en_i,
  reservation_i,
  flush_i,
  data_o,
  v_o,
  branch_o,
  btaken_o,
  npc_o,
  instr_misaligned_v_o
);

  input [520:0] reservation_i;
  output [65:0] data_o;
  output [38:0] npc_o;
  input clk_i;
  input reset_i;
  input en_i;
  input flush_i;
  output v_o;
  output branch_o;
  output btaken_o;
  output instr_misaligned_v_o;
  wire [65:0] data_o,ird_data_lo;
  wire [38:0] npc_o,baddr,ntaken_tgt;
  wire v_o,branch_o,btaken_o,instr_misaligned_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,
  N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,
  N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,
  N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,
  N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,
  N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,
  N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,
  N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,
  N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,
  N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,
  N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,
  N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,
  N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,
  N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,
  N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,
  N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,
  N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,
  N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,
  N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,
  N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,
  N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
  N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,
  N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,
  N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,
  N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,
  N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,
  N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,
  N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,
  N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,
  N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,
  N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,
  N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,
  N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,
  N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,
  N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,
  N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,
  N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,carry,sum_zero,N599,N600,N601,
  N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,
  N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,
  N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,comp_result,N646,N647,
  N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,
  N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,
  N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,
  N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,
  N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,
  N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
  N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,
  N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,N774,N775,
  N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,N790,N791,
  N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,N806,N807,
  N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,N822,N823,
  N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,N838,N839,
  N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,N854,N855,
  N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,N870,N871,
  N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,N886,N887,
  N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,N902,N903,
  N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,N918,N919,
  N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,N934,N935,
  N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,N950,N951,
  N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,N966,N967,
  N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,N982,N983,
  N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,N998,N999,
  N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012,
  N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,N1025,
  N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038,N1039,
  N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,
  N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,N1065,
  N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079,
  N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091,N1092,
  N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,N1105,
  N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118,N1119,
  N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,N1131,N1132,
  N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,
  N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
  N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,N1171,N1172,
  N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,N1185,
  N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,N1198,N1199,
  N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,N1211,N1212,
  N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
  N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,N1238,N1239,
  N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,N1251,N1252,
  N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,N1265,
  N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,N1278,N1279,
  N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,N1291,N1292,
  N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,N1305,
  N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,N1318,N1319,
  N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,N1331,N1332,
  N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,N1345,
  N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,N1358,N1359,
  N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,N1371,N1372,
  N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,N1385,
  N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,
  N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,N1411,N1412,
  N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,N1425,
  N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,N1438,N1439,
  N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,N1451,N1452,
  N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,N1465,
  N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478,N1479,
  N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,
  N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,N1505,
  N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,N1518,N1519,
  N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,N1531,N1532,
  N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,N1545,
  N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,N1558,N1559,
  N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,N1571,N1572,
  N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,N1585,
  N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,N1598,N1599,
  N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,N1611,N1612,
  N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,N1625,
  N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,N1638,N1639,
  N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,N1651,N1652,
  N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,N1665,
  N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,N1678,N1679,
  N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,N1691,N1692,
  N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,N1705,
  N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,N1718,N1719,
  N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,N1731,N1732,
  N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,N1745,
  N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,N1758,N1759,
  N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,N1771,N1772,
  N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,N1785,
  N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798,N1799,
  N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,N1811,N1812,
  N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,N1825,
  N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,N1838,N1839,
  N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,N1851,N1852,
  N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,N1865,
  N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,
  N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,N1891,N1892,
  N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,N1905,
  N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,N1919,
  N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,N1931,N1932,
  N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1945,
  N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,N1958,N1959,
  N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,
  N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,N1985,
  N1986,N1987,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,
  sv2v_dc_8,sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,
  sv2v_dc_15,sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,sv2v_dc_21,
  sv2v_dc_22,sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,sv2v_dc_27,sv2v_dc_28,sv2v_dc_29,
  sv2v_dc_30,sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,sv2v_dc_34,sv2v_dc_35,sv2v_dc_36,
  sv2v_dc_37,sv2v_dc_38,sv2v_dc_39,sv2v_dc_40,sv2v_dc_41,sv2v_dc_42,sv2v_dc_43,
  sv2v_dc_44,sv2v_dc_45,sv2v_dc_46,sv2v_dc_47,sv2v_dc_48,sv2v_dc_49,sv2v_dc_50,sv2v_dc_51,
  sv2v_dc_52,sv2v_dc_53,sv2v_dc_54,sv2v_dc_55,sv2v_dc_56,sv2v_dc_57,sv2v_dc_58,
  sv2v_dc_59,sv2v_dc_60,sv2v_dc_61,sv2v_dc_62,sv2v_dc_63,sv2v_dc_64,sv2v_dc_65,
  sv2v_dc_66;
  wire [5:5] shmask;
  wire [5:0] shamt,shamtn,clzh,clz,clzl,bindex;
  wire [38:1] taken_raw;
  wire [63:0] src1,src2,orcb,alu_result;
  wire [64:0] sum;
  wire [6:0] popcount;
  assign instr_misaligned_v_o = 1'b0;
  assign N49 = N46 & N47;
  assign N50 = N49 & N48;
  assign N51 = N46 | reservation_i[399];
  assign N52 = N51 | N48;
  assign N54 = N58 | N48;
  assign N56 = N51 | reservation_i[398];
  assign N58 = reservation_i[400] | N47;
  assign N59 = N58 | reservation_i[398];
  assign N61 = reservation_i[400] | reservation_i[399];
  assign N62 = N61 | N48;
  assign N63 = reservation_i[400] & reservation_i[399];
  assign N261 = N258 & N259;
  assign N262 = N261 & N260;
  assign N263 = reservation_i[397] | N259;
  assign N264 = N263 | N260;
  assign N266 = N258 | reservation_i[396];
  assign N267 = N266 | reservation_i[395];
  assign N269 = N258 | N259;
  assign N270 = N269 | reservation_i[395];
  assign N272 = reservation_i[397] & reservation_i[395];
  assign N273 = N263 | reservation_i[395];
  assign N274 = N259 & reservation_i[395];
  assign { sv2v_dc_1, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405 } = $signed(reservation_i[389:325]) >>> shamt;
  assign { sv2v_dc_2, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469 } = $signed(reservation_i[389:325]) >>> shamtn;
  assign N600 = N637 | reservation_i[407];
  assign N601 = reservation_i[406] | N638;
  assign N602 = N600 | N601;
  assign N603 = N602 | reservation_i[404];
  assign N604 = reservation_i[408] | reservation_i[407];
  assign N605 = N604 | N601;
  assign N606 = N605 | reservation_i[404];
  assign N609 = N602 | N608;
  assign N610 = N605 | N608;
  assign N612 = N642 | reservation_i[405];
  assign N613 = N600 | N612;
  assign N614 = N613 | reservation_i[404];
  assign N615 = reservation_i[408] | N634;
  assign N616 = N615 | N601;
  assign N617 = N616 | reservation_i[404];
  assign N619 = N613 | N608;
  assign N620 = N616 | N608;
  assign N622 = N642 | N638;
  assign N623 = N615 | N622;
  assign N624 = N623 | reservation_i[404];
  assign N626 = reservation_i[408] & reservation_i[407];
  assign N627 = N626 & reservation_i[404];
  assign N628 = reservation_i[406] & reservation_i[405];
  assign N629 = N628 & reservation_i[404];
  assign N630 = N637 & reservation_i[406];
  assign N631 = N630 & reservation_i[404];
  assign N632 = reservation_i[408] & reservation_i[406];
  assign N633 = N632 & reservation_i[405];
  assign N635 = N634 & reservation_i[406];
  assign N636 = N635 & reservation_i[405];
  assign N639 = N637 & N638;
  assign N640 = reservation_i[407] & N638;
  assign N641 = N640 & N608;
  assign N643 = N642 & N638;
  assign N644 = N626 & N642;

  bsg_popcount_width_p64
  popc
  (
    .i(reservation_i[388:325]),
    .o(popcount)
  );


  bsg_counting_leading_zeros_width_p32
  bclzh
  (
    .a_i(reservation_i[388:357]),
    .num_zero_o(clzh)
  );


  bsg_counting_leading_zeros_width_p32
  bclzl
  (
    .a_i(reservation_i[356:325]),
    .num_zero_o(clzl)
  );

  assign N653 = N599 & N637;
  assign N654 = N653 & N643;
  assign N655 = N654 & N608;
  assign N656 = reservation_i[409] | reservation_i[408];
  assign N657 = N656 | N612;
  assign N658 = N657 | reservation_i[404];
  assign N660 = reservation_i[409] | reservation_i[408];
  assign N661 = N660 | N622;
  assign N662 = N661 | reservation_i[404];
  assign N664 = reservation_i[409] | reservation_i[408];
  assign N665 = N664 | N622;
  assign N666 = N665 | N608;
  assign N668 = reservation_i[409] | N637;
  assign N669 = reservation_i[406] | reservation_i[405];
  assign N670 = N668 | N669;
  assign N671 = N670 | reservation_i[404];
  assign N673 = reservation_i[409] | N637;
  assign N674 = reservation_i[406] | reservation_i[405];
  assign N675 = N673 | N674;
  assign N676 = N675 | N608;
  assign N678 = reservation_i[409] | N637;
  assign N679 = N678 | N612;
  assign N680 = N679 | reservation_i[404];
  assign N681 = reservation_i[409] | N637;
  assign N682 = N681 | N612;
  assign N683 = N682 | N608;
  assign N684 = reservation_i[409] | N637;
  assign N685 = N684 | N601;
  assign N686 = N685 | reservation_i[404];
  assign N687 = reservation_i[409] | N637;
  assign N688 = N687 | N601;
  assign N689 = N688 | N608;
  assign N691 = reservation_i[409] | N637;
  assign N692 = N691 | N622;
  assign N693 = N692 | reservation_i[404];
  assign N695 = reservation_i[409] | N637;
  assign N696 = N695 | N622;
  assign N697 = N696 | N608;
  assign N699 = N599 | reservation_i[408];
  assign N700 = reservation_i[406] | reservation_i[405];
  assign N701 = N699 | N700;
  assign N702 = N701 | reservation_i[404];
  assign N704 = N599 | reservation_i[408];
  assign N705 = reservation_i[406] | reservation_i[405];
  assign N706 = N704 | N705;
  assign N707 = N706 | N608;
  assign N709 = N599 | reservation_i[408];
  assign N710 = N709 | N601;
  assign N711 = N710 | reservation_i[404];
  assign N713 = N599 | reservation_i[408];
  assign N714 = N713 | N612;
  assign N715 = N714 | reservation_i[404];
  assign N717 = reservation_i[409] & reservation_i[406];
  assign N718 = N717 & reservation_i[405];
  assign N719 = N638 & reservation_i[404];
  assign N720 = N630 & N719;
  assign N721 = reservation_i[409] & reservation_i[408];
  assign N722 = N599 & N637;
  assign N723 = N642 & reservation_i[404];
  assign N724 = N722 & N723;
  assign N725 = N637 & N642;
  assign N726 = reservation_i[405] & reservation_i[404];
  assign N727 = N725 & N726;
  assign N728 = N599 & N637;
  assign N729 = N642 & reservation_i[405];
  assign N730 = N728 & N729;

  bp_be_int_box_00
  box
  (
    .raw_i(alu_result),
    .tag_i(reservation_i[402:401]),
    .unsigned_i(1'b0),
    .reg_o(ird_data_lo)
  );

  assign { sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36, sv2v_dc_37, sv2v_dc_38, sv2v_dc_39, sv2v_dc_40, sv2v_dc_41, sv2v_dc_42, sv2v_dc_43, sv2v_dc_44, sv2v_dc_45, sv2v_dc_46, sv2v_dc_47, sv2v_dc_48, sv2v_dc_49, sv2v_dc_50, sv2v_dc_51, sv2v_dc_52, sv2v_dc_53, sv2v_dc_54, sv2v_dc_55, sv2v_dc_56, sv2v_dc_57, sv2v_dc_58, sv2v_dc_59, sv2v_dc_60, sv2v_dc_61, sv2v_dc_62, sv2v_dc_63, sv2v_dc_64, sv2v_dc_65, N1117 } = reservation_i[388:325] >> bindex;
  assign { N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << bindex;
  assign { N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << bindex;
  assign { N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << bindex;
  assign { N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130 } = reservation_i[388:325] << shamt;
  assign { N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194 } = reservation_i[388:325] << shamtn;
  assign N1441 = ~reservation_i[416];
  assign N1442 = N1441 | reservation_i[417];
  assign N1443 = ~N1442;
  assign ntaken_tgt = reservation_i[519:481] + { reservation_i[391:390], 1'b0 };
  assign { taken_raw, sv2v_dc_66 } = baddr + reservation_i[233:195];
  assign shamtn = { N1443, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } - shamt;
  assign { N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533 } = { src1[63:63], src1 } + { src2[63:63], src2 };
  assign { carry, sum } = { N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533 } + reservation_i[419];
  assign baddr = (N0)? reservation_i[363:325] : 
                 (N45)? reservation_i[519:481] : 1'b0;
  assign N0 = reservation_i[431];
  assign { N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66 } = (N1)? reservation_i[388:325] : 
                                                                                                                                                                                                                                                                                                                                                                            (N65)? { reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:519], reservation_i[519:481] } : 1'b0;
  assign N1 = reservation_i[440];
  assign src1 = (N2)? { N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66 } : 
                (N3)? { reservation_i[325:325], reservation_i[326:326], reservation_i[327:327], reservation_i[328:328], reservation_i[329:329], reservation_i[330:330], reservation_i[331:331], reservation_i[332:332], reservation_i[333:333], reservation_i[334:334], reservation_i[335:335], reservation_i[336:336], reservation_i[337:337], reservation_i[338:338], reservation_i[339:339], reservation_i[340:340], reservation_i[341:341], reservation_i[342:342], reservation_i[343:343], reservation_i[344:344], reservation_i[345:345], reservation_i[346:346], reservation_i[347:347], reservation_i[348:348], reservation_i[349:349], reservation_i[350:350], reservation_i[351:351], reservation_i[352:352], reservation_i[353:353], reservation_i[354:354], reservation_i[355:355], reservation_i[356:356], reservation_i[357:357], reservation_i[358:358], reservation_i[359:359], reservation_i[360:360], reservation_i[361:361], reservation_i[362:362], reservation_i[363:363], reservation_i[364:364], reservation_i[365:365], reservation_i[366:366], reservation_i[367:367], reservation_i[368:368], reservation_i[369:369], reservation_i[370:370], reservation_i[371:371], reservation_i[372:372], reservation_i[373:373], reservation_i[374:374], reservation_i[375:375], reservation_i[376:376], reservation_i[377:377], reservation_i[378:378], reservation_i[379:379], reservation_i[380:380], reservation_i[381:381], reservation_i[382:382], reservation_i[383:383], reservation_i[384:384], reservation_i[385:385], reservation_i[386:386], reservation_i[387:387], reservation_i[388:388] } : 
                (N4)? { N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130 } : 
                (N5)? { N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194 } : 
                (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2 = N50;
  assign N3 = N53;
  assign N4 = N55;
  assign N5 = N57;
  assign N6 = N60;
  assign N7 = N64;
  assign { N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277 } = (N8)? reservation_i[323:260] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N276)? reservation_i[258:195] : 1'b0;
  assign N8 = reservation_i[439];
  assign src2 = (N9)? { N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277 } : 
                (N10)? { N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404 } : 
                (N11)? { N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405 } : 
                (N12)? { N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469 } : 
                (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N9 = N262;
  assign N10 = N265;
  assign N11 = N268;
  assign N12 = N271;
  assign N13 = N275;
  assign N649 = (N14)? sum[64] : 
                (N15)? N646 : 
                (N16)? N647 : 
                (N17)? carry : 
                (N18)? N648 : 
                (N19)? sum_zero : 1'b0;
  assign N14 = N607;
  assign N15 = N611;
  assign N16 = N618;
  assign N17 = N621;
  assign N18 = N625;
  assign N19 = N645;
  assign comp_result = (N20)? N649 : 
                       (N21)? sum_zero : 1'b0;
  assign N20 = N599;
  assign N21 = reservation_i[409];
  assign clz = (N22)? clzh : 
               (N23)? { N651, clzl[4:0] } : 1'b0;
  assign N22 = N650;
  assign N23 = clzh[5];
  assign { N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925 } = (N24)? reservation_i[388:325] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N25)? reservation_i[323:260] : 1'b0;
  assign N24 = comp_result;
  assign N25 = N924;
  assign { N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374 } = (N26)? sum[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N27)? { N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772, N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783, N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794, N795 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N28)? { N796, N797, N798, N799, N800, N801, N802, N803, N804, N805, N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816, N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827, N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838, N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849, N850, N851, N852, N853, N854, N855, N856, N857, N858, N859 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N29)? { N860, N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871, N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882, N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893, N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904, N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915, N916, N917, N918, N919, N920, N921, N922, N923 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N30)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, popcount } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N31)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, clz } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N32)? { N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N33)? orcb : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N34)? { reservation_i[332:325], reservation_i[340:333], reservation_i[348:341], reservation_i[356:349], reservation_i[364:357], reservation_i[372:365], reservation_i[380:373], reservation_i[388:381] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N35)? { N1053, N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063, N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072, N1073, N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083, N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093, N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102, N1103, N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113, N1114, N1115, N1116 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N36)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1117 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N37)? { N1182, N1183, N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202, N1203, N1204, N1205, N1206, N1207, N1208, N1209, N1210, N1211, N1212, N1213, N1214, N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222, N1223, N1224, N1225, N1226, N1227, N1228, N1229, N1230, N1231, N1232, N1233, N1234, N1235, N1236, N1237, N1238, N1239, N1240, N1241, N1242, N1243, N1244, N1245 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N38)? { N1310, N1311, N1312, N1313, N1314, N1315, N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323, N1324, N1325, N1326, N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334, N1335, N1336, N1337, N1338, N1339, N1340, N1341, N1342, N1343, N1344, N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1354, N1355, N1356, N1357, N1358, N1359, N1360, N1361, N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1369, N1370, N1371, N1372, N1373 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N39)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, comp_result } : 1'b0;
  assign N26 = N655;
  assign N27 = N659;
  assign N28 = N663;
  assign N29 = N667;
  assign N30 = N672;
  assign N31 = N677;
  assign N32 = N690;
  assign N33 = N694;
  assign N34 = N698;
  assign N35 = N703;
  assign N36 = N708;
  assign N37 = N712;
  assign N38 = N716;
  assign N39 = N731;
  assign alu_result = (N40)? { N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374 } : 
                      (N41)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, comp_result } : 1'b0;
  assign N40 = N634;
  assign N41 = reservation_i[407];
  assign data_o = (N42)? { 1'b0, 1'b0, ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt[38:38], ntaken_tgt } : 
                  (N1439)? ird_data_lo : 1'b0;
  assign N42 = N1438;
  assign npc_o = (N43)? { taken_raw, 1'b0 } : 
                 (N44)? ntaken_tgt : 1'b0;
  assign N43 = btaken_o;
  assign N44 = N1440;
  assign shmask[5] = ~N1443;
  assign shamt[5] = N282 & shmask[5];
  assign shamt[4] = N281 & 1'b1;
  assign shamt[3] = N280 & 1'b1;
  assign shamt[2] = N279 & 1'b1;
  assign shamt[1] = N278 & 1'b1;
  assign shamt[0] = N277 & 1'b1;
  assign N45 = ~reservation_i[431];
  assign N46 = ~reservation_i[400];
  assign N47 = ~reservation_i[399];
  assign N48 = ~reservation_i[398];
  assign N53 = ~N52;
  assign N55 = ~N54;
  assign N57 = ~N56;
  assign N60 = ~N59;
  assign N64 = N1444 | N63;
  assign N1444 = ~N62;
  assign N65 = ~reservation_i[440];
  assign N258 = ~reservation_i[397];
  assign N259 = ~reservation_i[396];
  assign N260 = ~reservation_i[395];
  assign N265 = ~N264;
  assign N268 = ~N267;
  assign N271 = ~N270;
  assign N275 = N272 | N1446;
  assign N1446 = N1445 | N274;
  assign N1445 = ~N273;
  assign N276 = ~reservation_i[439];
  assign N341 = ~reservation_i[323];
  assign N342 = ~reservation_i[322];
  assign N343 = ~reservation_i[321];
  assign N344 = ~reservation_i[320];
  assign N345 = ~reservation_i[319];
  assign N346 = ~reservation_i[318];
  assign N347 = ~reservation_i[317];
  assign N348 = ~reservation_i[316];
  assign N349 = ~reservation_i[315];
  assign N350 = ~reservation_i[314];
  assign N351 = ~reservation_i[313];
  assign N352 = ~reservation_i[312];
  assign N353 = ~reservation_i[311];
  assign N354 = ~reservation_i[310];
  assign N355 = ~reservation_i[309];
  assign N356 = ~reservation_i[308];
  assign N357 = ~reservation_i[307];
  assign N358 = ~reservation_i[306];
  assign N359 = ~reservation_i[305];
  assign N360 = ~reservation_i[304];
  assign N361 = ~reservation_i[303];
  assign N362 = ~reservation_i[302];
  assign N363 = ~reservation_i[301];
  assign N364 = ~reservation_i[300];
  assign N365 = ~reservation_i[299];
  assign N366 = ~reservation_i[298];
  assign N367 = ~reservation_i[297];
  assign N368 = ~reservation_i[296];
  assign N369 = ~reservation_i[295];
  assign N370 = ~reservation_i[294];
  assign N371 = ~reservation_i[293];
  assign N372 = ~reservation_i[292];
  assign N373 = ~reservation_i[291];
  assign N374 = ~reservation_i[290];
  assign N375 = ~reservation_i[289];
  assign N376 = ~reservation_i[288];
  assign N377 = ~reservation_i[287];
  assign N378 = ~reservation_i[286];
  assign N379 = ~reservation_i[285];
  assign N380 = ~reservation_i[284];
  assign N381 = ~reservation_i[283];
  assign N382 = ~reservation_i[282];
  assign N383 = ~reservation_i[281];
  assign N384 = ~reservation_i[280];
  assign N385 = ~reservation_i[279];
  assign N386 = ~reservation_i[278];
  assign N387 = ~reservation_i[277];
  assign N388 = ~reservation_i[276];
  assign N389 = ~reservation_i[275];
  assign N390 = ~reservation_i[274];
  assign N391 = ~reservation_i[273];
  assign N392 = ~reservation_i[272];
  assign N393 = ~reservation_i[271];
  assign N394 = ~reservation_i[270];
  assign N395 = ~reservation_i[269];
  assign N396 = ~reservation_i[268];
  assign N397 = ~reservation_i[267];
  assign N398 = ~reservation_i[266];
  assign N399 = ~reservation_i[265];
  assign N400 = ~reservation_i[264];
  assign N401 = ~reservation_i[263];
  assign N402 = ~reservation_i[262];
  assign N403 = ~reservation_i[261];
  assign N404 = ~reservation_i[260];
  assign sum_zero = ~N1510;
  assign N1510 = N1509 | sum[0];
  assign N1509 = N1508 | sum[1];
  assign N1508 = N1507 | sum[2];
  assign N1507 = N1506 | sum[3];
  assign N1506 = N1505 | sum[4];
  assign N1505 = N1504 | sum[5];
  assign N1504 = N1503 | sum[6];
  assign N1503 = N1502 | sum[7];
  assign N1502 = N1501 | sum[8];
  assign N1501 = N1500 | sum[9];
  assign N1500 = N1499 | sum[10];
  assign N1499 = N1498 | sum[11];
  assign N1498 = N1497 | sum[12];
  assign N1497 = N1496 | sum[13];
  assign N1496 = N1495 | sum[14];
  assign N1495 = N1494 | sum[15];
  assign N1494 = N1493 | sum[16];
  assign N1493 = N1492 | sum[17];
  assign N1492 = N1491 | sum[18];
  assign N1491 = N1490 | sum[19];
  assign N1490 = N1489 | sum[20];
  assign N1489 = N1488 | sum[21];
  assign N1488 = N1487 | sum[22];
  assign N1487 = N1486 | sum[23];
  assign N1486 = N1485 | sum[24];
  assign N1485 = N1484 | sum[25];
  assign N1484 = N1483 | sum[26];
  assign N1483 = N1482 | sum[27];
  assign N1482 = N1481 | sum[28];
  assign N1481 = N1480 | sum[29];
  assign N1480 = N1479 | sum[30];
  assign N1479 = N1478 | sum[31];
  assign N1478 = N1477 | sum[32];
  assign N1477 = N1476 | sum[33];
  assign N1476 = N1475 | sum[34];
  assign N1475 = N1474 | sum[35];
  assign N1474 = N1473 | sum[36];
  assign N1473 = N1472 | sum[37];
  assign N1472 = N1471 | sum[38];
  assign N1471 = N1470 | sum[39];
  assign N1470 = N1469 | sum[40];
  assign N1469 = N1468 | sum[41];
  assign N1468 = N1467 | sum[42];
  assign N1467 = N1466 | sum[43];
  assign N1466 = N1465 | sum[44];
  assign N1465 = N1464 | sum[45];
  assign N1464 = N1463 | sum[46];
  assign N1463 = N1462 | sum[47];
  assign N1462 = N1461 | sum[48];
  assign N1461 = N1460 | sum[49];
  assign N1460 = N1459 | sum[50];
  assign N1459 = N1458 | sum[51];
  assign N1458 = N1457 | sum[52];
  assign N1457 = N1456 | sum[53];
  assign N1456 = N1455 | sum[54];
  assign N1455 = N1454 | sum[55];
  assign N1454 = N1453 | sum[56];
  assign N1453 = N1452 | sum[57];
  assign N1452 = N1451 | sum[58];
  assign N1451 = N1450 | sum[59];
  assign N1450 = N1449 | sum[60];
  assign N1449 = N1448 | sum[61];
  assign N1448 = N1447 | sum[62];
  assign N1447 = sum[64] | sum[63];
  assign N599 = ~reservation_i[409];
  assign N607 = N1511 | N1512;
  assign N1511 = ~N603;
  assign N1512 = ~N606;
  assign N608 = ~reservation_i[404];
  assign N611 = N1513 | N1514;
  assign N1513 = ~N609;
  assign N1514 = ~N610;
  assign N618 = N1515 | N1516;
  assign N1515 = ~N614;
  assign N1516 = ~N617;
  assign N621 = N1517 | N1518;
  assign N1517 = ~N619;
  assign N1518 = ~N620;
  assign N625 = ~N624;
  assign N634 = ~reservation_i[407];
  assign N637 = ~reservation_i[408];
  assign N638 = ~reservation_i[405];
  assign N642 = ~reservation_i[406];
  assign N645 = N627 | N1525;
  assign N1525 = N629 | N1524;
  assign N1524 = N631 | N1523;
  assign N1523 = N633 | N1522;
  assign N1522 = N636 | N1521;
  assign N1521 = N639 | N1520;
  assign N1520 = N641 | N1519;
  assign N1519 = N643 | N644;
  assign N646 = ~carry;
  assign N647 = ~sum[64];
  assign N648 = ~sum_zero;
  assign N650 = ~clzh[5];
  assign N651 = N1442 | clzl[5];
  assign orcb[7] = N1531 | reservation_i[325];
  assign N1531 = N1530 | reservation_i[326];
  assign N1530 = N1529 | reservation_i[327];
  assign N1529 = N1528 | reservation_i[328];
  assign N1528 = N1527 | reservation_i[329];
  assign N1527 = N1526 | reservation_i[330];
  assign N1526 = reservation_i[332] | reservation_i[331];
  assign orcb[6] = N1537 | reservation_i[325];
  assign N1537 = N1536 | reservation_i[326];
  assign N1536 = N1535 | reservation_i[327];
  assign N1535 = N1534 | reservation_i[328];
  assign N1534 = N1533 | reservation_i[329];
  assign N1533 = N1532 | reservation_i[330];
  assign N1532 = reservation_i[332] | reservation_i[331];
  assign orcb[5] = N1543 | reservation_i[325];
  assign N1543 = N1542 | reservation_i[326];
  assign N1542 = N1541 | reservation_i[327];
  assign N1541 = N1540 | reservation_i[328];
  assign N1540 = N1539 | reservation_i[329];
  assign N1539 = N1538 | reservation_i[330];
  assign N1538 = reservation_i[332] | reservation_i[331];
  assign orcb[4] = N1549 | reservation_i[325];
  assign N1549 = N1548 | reservation_i[326];
  assign N1548 = N1547 | reservation_i[327];
  assign N1547 = N1546 | reservation_i[328];
  assign N1546 = N1545 | reservation_i[329];
  assign N1545 = N1544 | reservation_i[330];
  assign N1544 = reservation_i[332] | reservation_i[331];
  assign orcb[3] = N1555 | reservation_i[325];
  assign N1555 = N1554 | reservation_i[326];
  assign N1554 = N1553 | reservation_i[327];
  assign N1553 = N1552 | reservation_i[328];
  assign N1552 = N1551 | reservation_i[329];
  assign N1551 = N1550 | reservation_i[330];
  assign N1550 = reservation_i[332] | reservation_i[331];
  assign orcb[2] = N1561 | reservation_i[325];
  assign N1561 = N1560 | reservation_i[326];
  assign N1560 = N1559 | reservation_i[327];
  assign N1559 = N1558 | reservation_i[328];
  assign N1558 = N1557 | reservation_i[329];
  assign N1557 = N1556 | reservation_i[330];
  assign N1556 = reservation_i[332] | reservation_i[331];
  assign orcb[1] = N1567 | reservation_i[325];
  assign N1567 = N1566 | reservation_i[326];
  assign N1566 = N1565 | reservation_i[327];
  assign N1565 = N1564 | reservation_i[328];
  assign N1564 = N1563 | reservation_i[329];
  assign N1563 = N1562 | reservation_i[330];
  assign N1562 = reservation_i[332] | reservation_i[331];
  assign orcb[0] = N1573 | reservation_i[325];
  assign N1573 = N1572 | reservation_i[326];
  assign N1572 = N1571 | reservation_i[327];
  assign N1571 = N1570 | reservation_i[328];
  assign N1570 = N1569 | reservation_i[329];
  assign N1569 = N1568 | reservation_i[330];
  assign N1568 = reservation_i[332] | reservation_i[331];
  assign orcb[15] = N1579 | reservation_i[333];
  assign N1579 = N1578 | reservation_i[334];
  assign N1578 = N1577 | reservation_i[335];
  assign N1577 = N1576 | reservation_i[336];
  assign N1576 = N1575 | reservation_i[337];
  assign N1575 = N1574 | reservation_i[338];
  assign N1574 = reservation_i[340] | reservation_i[339];
  assign orcb[14] = N1585 | reservation_i[333];
  assign N1585 = N1584 | reservation_i[334];
  assign N1584 = N1583 | reservation_i[335];
  assign N1583 = N1582 | reservation_i[336];
  assign N1582 = N1581 | reservation_i[337];
  assign N1581 = N1580 | reservation_i[338];
  assign N1580 = reservation_i[340] | reservation_i[339];
  assign orcb[13] = N1591 | reservation_i[333];
  assign N1591 = N1590 | reservation_i[334];
  assign N1590 = N1589 | reservation_i[335];
  assign N1589 = N1588 | reservation_i[336];
  assign N1588 = N1587 | reservation_i[337];
  assign N1587 = N1586 | reservation_i[338];
  assign N1586 = reservation_i[340] | reservation_i[339];
  assign orcb[12] = N1597 | reservation_i[333];
  assign N1597 = N1596 | reservation_i[334];
  assign N1596 = N1595 | reservation_i[335];
  assign N1595 = N1594 | reservation_i[336];
  assign N1594 = N1593 | reservation_i[337];
  assign N1593 = N1592 | reservation_i[338];
  assign N1592 = reservation_i[340] | reservation_i[339];
  assign orcb[11] = N1603 | reservation_i[333];
  assign N1603 = N1602 | reservation_i[334];
  assign N1602 = N1601 | reservation_i[335];
  assign N1601 = N1600 | reservation_i[336];
  assign N1600 = N1599 | reservation_i[337];
  assign N1599 = N1598 | reservation_i[338];
  assign N1598 = reservation_i[340] | reservation_i[339];
  assign orcb[10] = N1609 | reservation_i[333];
  assign N1609 = N1608 | reservation_i[334];
  assign N1608 = N1607 | reservation_i[335];
  assign N1607 = N1606 | reservation_i[336];
  assign N1606 = N1605 | reservation_i[337];
  assign N1605 = N1604 | reservation_i[338];
  assign N1604 = reservation_i[340] | reservation_i[339];
  assign orcb[9] = N1615 | reservation_i[333];
  assign N1615 = N1614 | reservation_i[334];
  assign N1614 = N1613 | reservation_i[335];
  assign N1613 = N1612 | reservation_i[336];
  assign N1612 = N1611 | reservation_i[337];
  assign N1611 = N1610 | reservation_i[338];
  assign N1610 = reservation_i[340] | reservation_i[339];
  assign orcb[8] = N1621 | reservation_i[333];
  assign N1621 = N1620 | reservation_i[334];
  assign N1620 = N1619 | reservation_i[335];
  assign N1619 = N1618 | reservation_i[336];
  assign N1618 = N1617 | reservation_i[337];
  assign N1617 = N1616 | reservation_i[338];
  assign N1616 = reservation_i[340] | reservation_i[339];
  assign orcb[23] = N1627 | reservation_i[341];
  assign N1627 = N1626 | reservation_i[342];
  assign N1626 = N1625 | reservation_i[343];
  assign N1625 = N1624 | reservation_i[344];
  assign N1624 = N1623 | reservation_i[345];
  assign N1623 = N1622 | reservation_i[346];
  assign N1622 = reservation_i[348] | reservation_i[347];
  assign orcb[22] = N1633 | reservation_i[341];
  assign N1633 = N1632 | reservation_i[342];
  assign N1632 = N1631 | reservation_i[343];
  assign N1631 = N1630 | reservation_i[344];
  assign N1630 = N1629 | reservation_i[345];
  assign N1629 = N1628 | reservation_i[346];
  assign N1628 = reservation_i[348] | reservation_i[347];
  assign orcb[21] = N1639 | reservation_i[341];
  assign N1639 = N1638 | reservation_i[342];
  assign N1638 = N1637 | reservation_i[343];
  assign N1637 = N1636 | reservation_i[344];
  assign N1636 = N1635 | reservation_i[345];
  assign N1635 = N1634 | reservation_i[346];
  assign N1634 = reservation_i[348] | reservation_i[347];
  assign orcb[20] = N1645 | reservation_i[341];
  assign N1645 = N1644 | reservation_i[342];
  assign N1644 = N1643 | reservation_i[343];
  assign N1643 = N1642 | reservation_i[344];
  assign N1642 = N1641 | reservation_i[345];
  assign N1641 = N1640 | reservation_i[346];
  assign N1640 = reservation_i[348] | reservation_i[347];
  assign orcb[19] = N1651 | reservation_i[341];
  assign N1651 = N1650 | reservation_i[342];
  assign N1650 = N1649 | reservation_i[343];
  assign N1649 = N1648 | reservation_i[344];
  assign N1648 = N1647 | reservation_i[345];
  assign N1647 = N1646 | reservation_i[346];
  assign N1646 = reservation_i[348] | reservation_i[347];
  assign orcb[18] = N1657 | reservation_i[341];
  assign N1657 = N1656 | reservation_i[342];
  assign N1656 = N1655 | reservation_i[343];
  assign N1655 = N1654 | reservation_i[344];
  assign N1654 = N1653 | reservation_i[345];
  assign N1653 = N1652 | reservation_i[346];
  assign N1652 = reservation_i[348] | reservation_i[347];
  assign orcb[17] = N1663 | reservation_i[341];
  assign N1663 = N1662 | reservation_i[342];
  assign N1662 = N1661 | reservation_i[343];
  assign N1661 = N1660 | reservation_i[344];
  assign N1660 = N1659 | reservation_i[345];
  assign N1659 = N1658 | reservation_i[346];
  assign N1658 = reservation_i[348] | reservation_i[347];
  assign orcb[16] = N1669 | reservation_i[341];
  assign N1669 = N1668 | reservation_i[342];
  assign N1668 = N1667 | reservation_i[343];
  assign N1667 = N1666 | reservation_i[344];
  assign N1666 = N1665 | reservation_i[345];
  assign N1665 = N1664 | reservation_i[346];
  assign N1664 = reservation_i[348] | reservation_i[347];
  assign orcb[31] = N1675 | reservation_i[349];
  assign N1675 = N1674 | reservation_i[350];
  assign N1674 = N1673 | reservation_i[351];
  assign N1673 = N1672 | reservation_i[352];
  assign N1672 = N1671 | reservation_i[353];
  assign N1671 = N1670 | reservation_i[354];
  assign N1670 = reservation_i[356] | reservation_i[355];
  assign orcb[30] = N1681 | reservation_i[349];
  assign N1681 = N1680 | reservation_i[350];
  assign N1680 = N1679 | reservation_i[351];
  assign N1679 = N1678 | reservation_i[352];
  assign N1678 = N1677 | reservation_i[353];
  assign N1677 = N1676 | reservation_i[354];
  assign N1676 = reservation_i[356] | reservation_i[355];
  assign orcb[29] = N1687 | reservation_i[349];
  assign N1687 = N1686 | reservation_i[350];
  assign N1686 = N1685 | reservation_i[351];
  assign N1685 = N1684 | reservation_i[352];
  assign N1684 = N1683 | reservation_i[353];
  assign N1683 = N1682 | reservation_i[354];
  assign N1682 = reservation_i[356] | reservation_i[355];
  assign orcb[28] = N1693 | reservation_i[349];
  assign N1693 = N1692 | reservation_i[350];
  assign N1692 = N1691 | reservation_i[351];
  assign N1691 = N1690 | reservation_i[352];
  assign N1690 = N1689 | reservation_i[353];
  assign N1689 = N1688 | reservation_i[354];
  assign N1688 = reservation_i[356] | reservation_i[355];
  assign orcb[27] = N1699 | reservation_i[349];
  assign N1699 = N1698 | reservation_i[350];
  assign N1698 = N1697 | reservation_i[351];
  assign N1697 = N1696 | reservation_i[352];
  assign N1696 = N1695 | reservation_i[353];
  assign N1695 = N1694 | reservation_i[354];
  assign N1694 = reservation_i[356] | reservation_i[355];
  assign orcb[26] = N1705 | reservation_i[349];
  assign N1705 = N1704 | reservation_i[350];
  assign N1704 = N1703 | reservation_i[351];
  assign N1703 = N1702 | reservation_i[352];
  assign N1702 = N1701 | reservation_i[353];
  assign N1701 = N1700 | reservation_i[354];
  assign N1700 = reservation_i[356] | reservation_i[355];
  assign orcb[25] = N1711 | reservation_i[349];
  assign N1711 = N1710 | reservation_i[350];
  assign N1710 = N1709 | reservation_i[351];
  assign N1709 = N1708 | reservation_i[352];
  assign N1708 = N1707 | reservation_i[353];
  assign N1707 = N1706 | reservation_i[354];
  assign N1706 = reservation_i[356] | reservation_i[355];
  assign orcb[24] = N1717 | reservation_i[349];
  assign N1717 = N1716 | reservation_i[350];
  assign N1716 = N1715 | reservation_i[351];
  assign N1715 = N1714 | reservation_i[352];
  assign N1714 = N1713 | reservation_i[353];
  assign N1713 = N1712 | reservation_i[354];
  assign N1712 = reservation_i[356] | reservation_i[355];
  assign orcb[39] = N1723 | reservation_i[357];
  assign N1723 = N1722 | reservation_i[358];
  assign N1722 = N1721 | reservation_i[359];
  assign N1721 = N1720 | reservation_i[360];
  assign N1720 = N1719 | reservation_i[361];
  assign N1719 = N1718 | reservation_i[362];
  assign N1718 = reservation_i[364] | reservation_i[363];
  assign orcb[38] = N1729 | reservation_i[357];
  assign N1729 = N1728 | reservation_i[358];
  assign N1728 = N1727 | reservation_i[359];
  assign N1727 = N1726 | reservation_i[360];
  assign N1726 = N1725 | reservation_i[361];
  assign N1725 = N1724 | reservation_i[362];
  assign N1724 = reservation_i[364] | reservation_i[363];
  assign orcb[37] = N1735 | reservation_i[357];
  assign N1735 = N1734 | reservation_i[358];
  assign N1734 = N1733 | reservation_i[359];
  assign N1733 = N1732 | reservation_i[360];
  assign N1732 = N1731 | reservation_i[361];
  assign N1731 = N1730 | reservation_i[362];
  assign N1730 = reservation_i[364] | reservation_i[363];
  assign orcb[36] = N1741 | reservation_i[357];
  assign N1741 = N1740 | reservation_i[358];
  assign N1740 = N1739 | reservation_i[359];
  assign N1739 = N1738 | reservation_i[360];
  assign N1738 = N1737 | reservation_i[361];
  assign N1737 = N1736 | reservation_i[362];
  assign N1736 = reservation_i[364] | reservation_i[363];
  assign orcb[35] = N1747 | reservation_i[357];
  assign N1747 = N1746 | reservation_i[358];
  assign N1746 = N1745 | reservation_i[359];
  assign N1745 = N1744 | reservation_i[360];
  assign N1744 = N1743 | reservation_i[361];
  assign N1743 = N1742 | reservation_i[362];
  assign N1742 = reservation_i[364] | reservation_i[363];
  assign orcb[34] = N1753 | reservation_i[357];
  assign N1753 = N1752 | reservation_i[358];
  assign N1752 = N1751 | reservation_i[359];
  assign N1751 = N1750 | reservation_i[360];
  assign N1750 = N1749 | reservation_i[361];
  assign N1749 = N1748 | reservation_i[362];
  assign N1748 = reservation_i[364] | reservation_i[363];
  assign orcb[33] = N1759 | reservation_i[357];
  assign N1759 = N1758 | reservation_i[358];
  assign N1758 = N1757 | reservation_i[359];
  assign N1757 = N1756 | reservation_i[360];
  assign N1756 = N1755 | reservation_i[361];
  assign N1755 = N1754 | reservation_i[362];
  assign N1754 = reservation_i[364] | reservation_i[363];
  assign orcb[32] = N1765 | reservation_i[357];
  assign N1765 = N1764 | reservation_i[358];
  assign N1764 = N1763 | reservation_i[359];
  assign N1763 = N1762 | reservation_i[360];
  assign N1762 = N1761 | reservation_i[361];
  assign N1761 = N1760 | reservation_i[362];
  assign N1760 = reservation_i[364] | reservation_i[363];
  assign orcb[47] = N1771 | reservation_i[365];
  assign N1771 = N1770 | reservation_i[366];
  assign N1770 = N1769 | reservation_i[367];
  assign N1769 = N1768 | reservation_i[368];
  assign N1768 = N1767 | reservation_i[369];
  assign N1767 = N1766 | reservation_i[370];
  assign N1766 = reservation_i[372] | reservation_i[371];
  assign orcb[46] = N1777 | reservation_i[365];
  assign N1777 = N1776 | reservation_i[366];
  assign N1776 = N1775 | reservation_i[367];
  assign N1775 = N1774 | reservation_i[368];
  assign N1774 = N1773 | reservation_i[369];
  assign N1773 = N1772 | reservation_i[370];
  assign N1772 = reservation_i[372] | reservation_i[371];
  assign orcb[45] = N1783 | reservation_i[365];
  assign N1783 = N1782 | reservation_i[366];
  assign N1782 = N1781 | reservation_i[367];
  assign N1781 = N1780 | reservation_i[368];
  assign N1780 = N1779 | reservation_i[369];
  assign N1779 = N1778 | reservation_i[370];
  assign N1778 = reservation_i[372] | reservation_i[371];
  assign orcb[44] = N1789 | reservation_i[365];
  assign N1789 = N1788 | reservation_i[366];
  assign N1788 = N1787 | reservation_i[367];
  assign N1787 = N1786 | reservation_i[368];
  assign N1786 = N1785 | reservation_i[369];
  assign N1785 = N1784 | reservation_i[370];
  assign N1784 = reservation_i[372] | reservation_i[371];
  assign orcb[43] = N1795 | reservation_i[365];
  assign N1795 = N1794 | reservation_i[366];
  assign N1794 = N1793 | reservation_i[367];
  assign N1793 = N1792 | reservation_i[368];
  assign N1792 = N1791 | reservation_i[369];
  assign N1791 = N1790 | reservation_i[370];
  assign N1790 = reservation_i[372] | reservation_i[371];
  assign orcb[42] = N1801 | reservation_i[365];
  assign N1801 = N1800 | reservation_i[366];
  assign N1800 = N1799 | reservation_i[367];
  assign N1799 = N1798 | reservation_i[368];
  assign N1798 = N1797 | reservation_i[369];
  assign N1797 = N1796 | reservation_i[370];
  assign N1796 = reservation_i[372] | reservation_i[371];
  assign orcb[41] = N1807 | reservation_i[365];
  assign N1807 = N1806 | reservation_i[366];
  assign N1806 = N1805 | reservation_i[367];
  assign N1805 = N1804 | reservation_i[368];
  assign N1804 = N1803 | reservation_i[369];
  assign N1803 = N1802 | reservation_i[370];
  assign N1802 = reservation_i[372] | reservation_i[371];
  assign orcb[40] = N1813 | reservation_i[365];
  assign N1813 = N1812 | reservation_i[366];
  assign N1812 = N1811 | reservation_i[367];
  assign N1811 = N1810 | reservation_i[368];
  assign N1810 = N1809 | reservation_i[369];
  assign N1809 = N1808 | reservation_i[370];
  assign N1808 = reservation_i[372] | reservation_i[371];
  assign orcb[55] = N1819 | reservation_i[373];
  assign N1819 = N1818 | reservation_i[374];
  assign N1818 = N1817 | reservation_i[375];
  assign N1817 = N1816 | reservation_i[376];
  assign N1816 = N1815 | reservation_i[377];
  assign N1815 = N1814 | reservation_i[378];
  assign N1814 = reservation_i[380] | reservation_i[379];
  assign orcb[54] = N1825 | reservation_i[373];
  assign N1825 = N1824 | reservation_i[374];
  assign N1824 = N1823 | reservation_i[375];
  assign N1823 = N1822 | reservation_i[376];
  assign N1822 = N1821 | reservation_i[377];
  assign N1821 = N1820 | reservation_i[378];
  assign N1820 = reservation_i[380] | reservation_i[379];
  assign orcb[53] = N1831 | reservation_i[373];
  assign N1831 = N1830 | reservation_i[374];
  assign N1830 = N1829 | reservation_i[375];
  assign N1829 = N1828 | reservation_i[376];
  assign N1828 = N1827 | reservation_i[377];
  assign N1827 = N1826 | reservation_i[378];
  assign N1826 = reservation_i[380] | reservation_i[379];
  assign orcb[52] = N1837 | reservation_i[373];
  assign N1837 = N1836 | reservation_i[374];
  assign N1836 = N1835 | reservation_i[375];
  assign N1835 = N1834 | reservation_i[376];
  assign N1834 = N1833 | reservation_i[377];
  assign N1833 = N1832 | reservation_i[378];
  assign N1832 = reservation_i[380] | reservation_i[379];
  assign orcb[51] = N1843 | reservation_i[373];
  assign N1843 = N1842 | reservation_i[374];
  assign N1842 = N1841 | reservation_i[375];
  assign N1841 = N1840 | reservation_i[376];
  assign N1840 = N1839 | reservation_i[377];
  assign N1839 = N1838 | reservation_i[378];
  assign N1838 = reservation_i[380] | reservation_i[379];
  assign orcb[50] = N1849 | reservation_i[373];
  assign N1849 = N1848 | reservation_i[374];
  assign N1848 = N1847 | reservation_i[375];
  assign N1847 = N1846 | reservation_i[376];
  assign N1846 = N1845 | reservation_i[377];
  assign N1845 = N1844 | reservation_i[378];
  assign N1844 = reservation_i[380] | reservation_i[379];
  assign orcb[49] = N1855 | reservation_i[373];
  assign N1855 = N1854 | reservation_i[374];
  assign N1854 = N1853 | reservation_i[375];
  assign N1853 = N1852 | reservation_i[376];
  assign N1852 = N1851 | reservation_i[377];
  assign N1851 = N1850 | reservation_i[378];
  assign N1850 = reservation_i[380] | reservation_i[379];
  assign orcb[48] = N1861 | reservation_i[373];
  assign N1861 = N1860 | reservation_i[374];
  assign N1860 = N1859 | reservation_i[375];
  assign N1859 = N1858 | reservation_i[376];
  assign N1858 = N1857 | reservation_i[377];
  assign N1857 = N1856 | reservation_i[378];
  assign N1856 = reservation_i[380] | reservation_i[379];
  assign orcb[63] = N1867 | reservation_i[381];
  assign N1867 = N1866 | reservation_i[382];
  assign N1866 = N1865 | reservation_i[383];
  assign N1865 = N1864 | reservation_i[384];
  assign N1864 = N1863 | reservation_i[385];
  assign N1863 = N1862 | reservation_i[386];
  assign N1862 = reservation_i[388] | reservation_i[387];
  assign orcb[62] = N1873 | reservation_i[381];
  assign N1873 = N1872 | reservation_i[382];
  assign N1872 = N1871 | reservation_i[383];
  assign N1871 = N1870 | reservation_i[384];
  assign N1870 = N1869 | reservation_i[385];
  assign N1869 = N1868 | reservation_i[386];
  assign N1868 = reservation_i[388] | reservation_i[387];
  assign orcb[61] = N1879 | reservation_i[381];
  assign N1879 = N1878 | reservation_i[382];
  assign N1878 = N1877 | reservation_i[383];
  assign N1877 = N1876 | reservation_i[384];
  assign N1876 = N1875 | reservation_i[385];
  assign N1875 = N1874 | reservation_i[386];
  assign N1874 = reservation_i[388] | reservation_i[387];
  assign orcb[60] = N1885 | reservation_i[381];
  assign N1885 = N1884 | reservation_i[382];
  assign N1884 = N1883 | reservation_i[383];
  assign N1883 = N1882 | reservation_i[384];
  assign N1882 = N1881 | reservation_i[385];
  assign N1881 = N1880 | reservation_i[386];
  assign N1880 = reservation_i[388] | reservation_i[387];
  assign orcb[59] = N1891 | reservation_i[381];
  assign N1891 = N1890 | reservation_i[382];
  assign N1890 = N1889 | reservation_i[383];
  assign N1889 = N1888 | reservation_i[384];
  assign N1888 = N1887 | reservation_i[385];
  assign N1887 = N1886 | reservation_i[386];
  assign N1886 = reservation_i[388] | reservation_i[387];
  assign orcb[58] = N1897 | reservation_i[381];
  assign N1897 = N1896 | reservation_i[382];
  assign N1896 = N1895 | reservation_i[383];
  assign N1895 = N1894 | reservation_i[384];
  assign N1894 = N1893 | reservation_i[385];
  assign N1893 = N1892 | reservation_i[386];
  assign N1892 = reservation_i[388] | reservation_i[387];
  assign orcb[57] = N1903 | reservation_i[381];
  assign N1903 = N1902 | reservation_i[382];
  assign N1902 = N1901 | reservation_i[383];
  assign N1901 = N1900 | reservation_i[384];
  assign N1900 = N1899 | reservation_i[385];
  assign N1899 = N1898 | reservation_i[386];
  assign N1898 = reservation_i[388] | reservation_i[387];
  assign orcb[56] = N1909 | reservation_i[381];
  assign N1909 = N1908 | reservation_i[382];
  assign N1908 = N1907 | reservation_i[383];
  assign N1907 = N1906 | reservation_i[384];
  assign N1906 = N1905 | reservation_i[385];
  assign N1905 = N1904 | reservation_i[386];
  assign N1904 = reservation_i[388] | reservation_i[387];
  assign bindex[5] = src2[5] & shmask[5];
  assign bindex[4] = src2[4] & 1'b1;
  assign bindex[3] = src2[3] & 1'b1;
  assign bindex[2] = src2[2] & 1'b1;
  assign bindex[1] = src2[1] & 1'b1;
  assign bindex[0] = src2[0] & 1'b1;
  assign N652 = N634;
  assign N659 = ~N658;
  assign N663 = ~N662;
  assign N667 = ~N666;
  assign N672 = ~N671;
  assign N677 = ~N676;
  assign N690 = N1914 | N1915;
  assign N1914 = N1912 | N1913;
  assign N1912 = N1910 | N1911;
  assign N1910 = ~N680;
  assign N1911 = ~N683;
  assign N1913 = ~N686;
  assign N1915 = ~N689;
  assign N694 = ~N693;
  assign N698 = ~N697;
  assign N703 = ~N702;
  assign N708 = ~N707;
  assign N712 = ~N711;
  assign N716 = ~N715;
  assign N731 = N718 | N1919;
  assign N1919 = N720 | N1918;
  assign N1918 = N721 | N1917;
  assign N1917 = N724 | N1916;
  assign N1916 = N727 | N730;
  assign N732 = src1[63] ^ src2[63];
  assign N733 = src1[62] ^ src2[62];
  assign N734 = src1[61] ^ src2[61];
  assign N735 = src1[60] ^ src2[60];
  assign N736 = src1[59] ^ src2[59];
  assign N737 = src1[58] ^ src2[58];
  assign N738 = src1[57] ^ src2[57];
  assign N739 = src1[56] ^ src2[56];
  assign N740 = src1[55] ^ src2[55];
  assign N741 = src1[54] ^ src2[54];
  assign N742 = src1[53] ^ src2[53];
  assign N743 = src1[52] ^ src2[52];
  assign N744 = src1[51] ^ src2[51];
  assign N745 = src1[50] ^ src2[50];
  assign N746 = src1[49] ^ src2[49];
  assign N747 = src1[48] ^ src2[48];
  assign N748 = src1[47] ^ src2[47];
  assign N749 = src1[46] ^ src2[46];
  assign N750 = src1[45] ^ src2[45];
  assign N751 = src1[44] ^ src2[44];
  assign N752 = src1[43] ^ src2[43];
  assign N753 = src1[42] ^ src2[42];
  assign N754 = src1[41] ^ src2[41];
  assign N755 = src1[40] ^ src2[40];
  assign N756 = src1[39] ^ src2[39];
  assign N757 = src1[38] ^ src2[38];
  assign N758 = src1[37] ^ src2[37];
  assign N759 = src1[36] ^ src2[36];
  assign N760 = src1[35] ^ src2[35];
  assign N761 = src1[34] ^ src2[34];
  assign N762 = src1[33] ^ src2[33];
  assign N763 = src1[32] ^ src2[32];
  assign N764 = src1[31] ^ src2[31];
  assign N765 = src1[30] ^ src2[30];
  assign N766 = src1[29] ^ src2[29];
  assign N767 = src1[28] ^ src2[28];
  assign N768 = src1[27] ^ src2[27];
  assign N769 = src1[26] ^ src2[26];
  assign N770 = src1[25] ^ src2[25];
  assign N771 = src1[24] ^ src2[24];
  assign N772 = src1[23] ^ src2[23];
  assign N773 = src1[22] ^ src2[22];
  assign N774 = src1[21] ^ src2[21];
  assign N775 = src1[20] ^ src2[20];
  assign N776 = src1[19] ^ src2[19];
  assign N777 = src1[18] ^ src2[18];
  assign N778 = src1[17] ^ src2[17];
  assign N779 = src1[16] ^ src2[16];
  assign N780 = src1[15] ^ src2[15];
  assign N781 = src1[14] ^ src2[14];
  assign N782 = src1[13] ^ src2[13];
  assign N783 = src1[12] ^ src2[12];
  assign N784 = src1[11] ^ src2[11];
  assign N785 = src1[10] ^ src2[10];
  assign N786 = src1[9] ^ src2[9];
  assign N787 = src1[8] ^ src2[8];
  assign N788 = src1[7] ^ src2[7];
  assign N789 = src1[6] ^ src2[6];
  assign N790 = src1[5] ^ src2[5];
  assign N791 = src1[4] ^ src2[4];
  assign N792 = src1[3] ^ src2[3];
  assign N793 = src1[2] ^ src2[2];
  assign N794 = src1[1] ^ src2[1];
  assign N795 = src1[0] ^ src2[0];
  assign N796 = src1[63] | src2[63];
  assign N797 = src1[62] | src2[62];
  assign N798 = src1[61] | src2[61];
  assign N799 = src1[60] | src2[60];
  assign N800 = src1[59] | src2[59];
  assign N801 = src1[58] | src2[58];
  assign N802 = src1[57] | src2[57];
  assign N803 = src1[56] | src2[56];
  assign N804 = src1[55] | src2[55];
  assign N805 = src1[54] | src2[54];
  assign N806 = src1[53] | src2[53];
  assign N807 = src1[52] | src2[52];
  assign N808 = src1[51] | src2[51];
  assign N809 = src1[50] | src2[50];
  assign N810 = src1[49] | src2[49];
  assign N811 = src1[48] | src2[48];
  assign N812 = src1[47] | src2[47];
  assign N813 = src1[46] | src2[46];
  assign N814 = src1[45] | src2[45];
  assign N815 = src1[44] | src2[44];
  assign N816 = src1[43] | src2[43];
  assign N817 = src1[42] | src2[42];
  assign N818 = src1[41] | src2[41];
  assign N819 = src1[40] | src2[40];
  assign N820 = src1[39] | src2[39];
  assign N821 = src1[38] | src2[38];
  assign N822 = src1[37] | src2[37];
  assign N823 = src1[36] | src2[36];
  assign N824 = src1[35] | src2[35];
  assign N825 = src1[34] | src2[34];
  assign N826 = src1[33] | src2[33];
  assign N827 = src1[32] | src2[32];
  assign N828 = src1[31] | src2[31];
  assign N829 = src1[30] | src2[30];
  assign N830 = src1[29] | src2[29];
  assign N831 = src1[28] | src2[28];
  assign N832 = src1[27] | src2[27];
  assign N833 = src1[26] | src2[26];
  assign N834 = src1[25] | src2[25];
  assign N835 = src1[24] | src2[24];
  assign N836 = src1[23] | src2[23];
  assign N837 = src1[22] | src2[22];
  assign N838 = src1[21] | src2[21];
  assign N839 = src1[20] | src2[20];
  assign N840 = src1[19] | src2[19];
  assign N841 = src1[18] | src2[18];
  assign N842 = src1[17] | src2[17];
  assign N843 = src1[16] | src2[16];
  assign N844 = src1[15] | src2[15];
  assign N845 = src1[14] | src2[14];
  assign N846 = src1[13] | src2[13];
  assign N847 = src1[12] | src2[12];
  assign N848 = src1[11] | src2[11];
  assign N849 = src1[10] | src2[10];
  assign N850 = src1[9] | src2[9];
  assign N851 = src1[8] | src2[8];
  assign N852 = src1[7] | src2[7];
  assign N853 = src1[6] | src2[6];
  assign N854 = src1[5] | src2[5];
  assign N855 = src1[4] | src2[4];
  assign N856 = src1[3] | src2[3];
  assign N857 = src1[2] | src2[2];
  assign N858 = src1[1] | src2[1];
  assign N859 = src1[0] | src2[0];
  assign N860 = src1[63] & src2[63];
  assign N861 = src1[62] & src2[62];
  assign N862 = src1[61] & src2[61];
  assign N863 = src1[60] & src2[60];
  assign N864 = src1[59] & src2[59];
  assign N865 = src1[58] & src2[58];
  assign N866 = src1[57] & src2[57];
  assign N867 = src1[56] & src2[56];
  assign N868 = src1[55] & src2[55];
  assign N869 = src1[54] & src2[54];
  assign N870 = src1[53] & src2[53];
  assign N871 = src1[52] & src2[52];
  assign N872 = src1[51] & src2[51];
  assign N873 = src1[50] & src2[50];
  assign N874 = src1[49] & src2[49];
  assign N875 = src1[48] & src2[48];
  assign N876 = src1[47] & src2[47];
  assign N877 = src1[46] & src2[46];
  assign N878 = src1[45] & src2[45];
  assign N879 = src1[44] & src2[44];
  assign N880 = src1[43] & src2[43];
  assign N881 = src1[42] & src2[42];
  assign N882 = src1[41] & src2[41];
  assign N883 = src1[40] & src2[40];
  assign N884 = src1[39] & src2[39];
  assign N885 = src1[38] & src2[38];
  assign N886 = src1[37] & src2[37];
  assign N887 = src1[36] & src2[36];
  assign N888 = src1[35] & src2[35];
  assign N889 = src1[34] & src2[34];
  assign N890 = src1[33] & src2[33];
  assign N891 = src1[32] & src2[32];
  assign N892 = src1[31] & src2[31];
  assign N893 = src1[30] & src2[30];
  assign N894 = src1[29] & src2[29];
  assign N895 = src1[28] & src2[28];
  assign N896 = src1[27] & src2[27];
  assign N897 = src1[26] & src2[26];
  assign N898 = src1[25] & src2[25];
  assign N899 = src1[24] & src2[24];
  assign N900 = src1[23] & src2[23];
  assign N901 = src1[22] & src2[22];
  assign N902 = src1[21] & src2[21];
  assign N903 = src1[20] & src2[20];
  assign N904 = src1[19] & src2[19];
  assign N905 = src1[18] & src2[18];
  assign N906 = src1[17] & src2[17];
  assign N907 = src1[16] & src2[16];
  assign N908 = src1[15] & src2[15];
  assign N909 = src1[14] & src2[14];
  assign N910 = src1[13] & src2[13];
  assign N911 = src1[12] & src2[12];
  assign N912 = src1[11] & src2[11];
  assign N913 = src1[10] & src2[10];
  assign N914 = src1[9] & src2[9];
  assign N915 = src1[8] & src2[8];
  assign N916 = src1[7] & src2[7];
  assign N917 = src1[6] & src2[6];
  assign N918 = src1[5] & src2[5];
  assign N919 = src1[4] & src2[4];
  assign N920 = src1[3] & src2[3];
  assign N921 = src1[2] & src2[2];
  assign N922 = src1[1] & src2[1];
  assign N923 = src1[0] & src2[0];
  assign N924 = ~comp_result;
  assign N1053 = reservation_i[388] & N1920;
  assign N1920 = ~N1052;
  assign N1054 = reservation_i[387] & N1921;
  assign N1921 = ~N1051;
  assign N1055 = reservation_i[386] & N1922;
  assign N1922 = ~N1050;
  assign N1056 = reservation_i[385] & N1923;
  assign N1923 = ~N1049;
  assign N1057 = reservation_i[384] & N1924;
  assign N1924 = ~N1048;
  assign N1058 = reservation_i[383] & N1925;
  assign N1925 = ~N1047;
  assign N1059 = reservation_i[382] & N1926;
  assign N1926 = ~N1046;
  assign N1060 = reservation_i[381] & N1927;
  assign N1927 = ~N1045;
  assign N1061 = reservation_i[380] & N1928;
  assign N1928 = ~N1044;
  assign N1062 = reservation_i[379] & N1929;
  assign N1929 = ~N1043;
  assign N1063 = reservation_i[378] & N1930;
  assign N1930 = ~N1042;
  assign N1064 = reservation_i[377] & N1931;
  assign N1931 = ~N1041;
  assign N1065 = reservation_i[376] & N1932;
  assign N1932 = ~N1040;
  assign N1066 = reservation_i[375] & N1933;
  assign N1933 = ~N1039;
  assign N1067 = reservation_i[374] & N1934;
  assign N1934 = ~N1038;
  assign N1068 = reservation_i[373] & N1935;
  assign N1935 = ~N1037;
  assign N1069 = reservation_i[372] & N1936;
  assign N1936 = ~N1036;
  assign N1070 = reservation_i[371] & N1937;
  assign N1937 = ~N1035;
  assign N1071 = reservation_i[370] & N1938;
  assign N1938 = ~N1034;
  assign N1072 = reservation_i[369] & N1939;
  assign N1939 = ~N1033;
  assign N1073 = reservation_i[368] & N1940;
  assign N1940 = ~N1032;
  assign N1074 = reservation_i[367] & N1941;
  assign N1941 = ~N1031;
  assign N1075 = reservation_i[366] & N1942;
  assign N1942 = ~N1030;
  assign N1076 = reservation_i[365] & N1943;
  assign N1943 = ~N1029;
  assign N1077 = reservation_i[364] & N1944;
  assign N1944 = ~N1028;
  assign N1078 = reservation_i[363] & N1945;
  assign N1945 = ~N1027;
  assign N1079 = reservation_i[362] & N1946;
  assign N1946 = ~N1026;
  assign N1080 = reservation_i[361] & N1947;
  assign N1947 = ~N1025;
  assign N1081 = reservation_i[360] & N1948;
  assign N1948 = ~N1024;
  assign N1082 = reservation_i[359] & N1949;
  assign N1949 = ~N1023;
  assign N1083 = reservation_i[358] & N1950;
  assign N1950 = ~N1022;
  assign N1084 = reservation_i[357] & N1951;
  assign N1951 = ~N1021;
  assign N1085 = reservation_i[356] & N1952;
  assign N1952 = ~N1020;
  assign N1086 = reservation_i[355] & N1953;
  assign N1953 = ~N1019;
  assign N1087 = reservation_i[354] & N1954;
  assign N1954 = ~N1018;
  assign N1088 = reservation_i[353] & N1955;
  assign N1955 = ~N1017;
  assign N1089 = reservation_i[352] & N1956;
  assign N1956 = ~N1016;
  assign N1090 = reservation_i[351] & N1957;
  assign N1957 = ~N1015;
  assign N1091 = reservation_i[350] & N1958;
  assign N1958 = ~N1014;
  assign N1092 = reservation_i[349] & N1959;
  assign N1959 = ~N1013;
  assign N1093 = reservation_i[348] & N1960;
  assign N1960 = ~N1012;
  assign N1094 = reservation_i[347] & N1961;
  assign N1961 = ~N1011;
  assign N1095 = reservation_i[346] & N1962;
  assign N1962 = ~N1010;
  assign N1096 = reservation_i[345] & N1963;
  assign N1963 = ~N1009;
  assign N1097 = reservation_i[344] & N1964;
  assign N1964 = ~N1008;
  assign N1098 = reservation_i[343] & N1965;
  assign N1965 = ~N1007;
  assign N1099 = reservation_i[342] & N1966;
  assign N1966 = ~N1006;
  assign N1100 = reservation_i[341] & N1967;
  assign N1967 = ~N1005;
  assign N1101 = reservation_i[340] & N1968;
  assign N1968 = ~N1004;
  assign N1102 = reservation_i[339] & N1969;
  assign N1969 = ~N1003;
  assign N1103 = reservation_i[338] & N1970;
  assign N1970 = ~N1002;
  assign N1104 = reservation_i[337] & N1971;
  assign N1971 = ~N1001;
  assign N1105 = reservation_i[336] & N1972;
  assign N1972 = ~N1000;
  assign N1106 = reservation_i[335] & N1973;
  assign N1973 = ~N999;
  assign N1107 = reservation_i[334] & N1974;
  assign N1974 = ~N998;
  assign N1108 = reservation_i[333] & N1975;
  assign N1975 = ~N997;
  assign N1109 = reservation_i[332] & N1976;
  assign N1976 = ~N996;
  assign N1110 = reservation_i[331] & N1977;
  assign N1977 = ~N995;
  assign N1111 = reservation_i[330] & N1978;
  assign N1978 = ~N994;
  assign N1112 = reservation_i[329] & N1979;
  assign N1979 = ~N993;
  assign N1113 = reservation_i[328] & N1980;
  assign N1980 = ~N992;
  assign N1114 = reservation_i[327] & N1981;
  assign N1981 = ~N991;
  assign N1115 = reservation_i[326] & N1982;
  assign N1982 = ~N990;
  assign N1116 = reservation_i[325] & N1983;
  assign N1983 = ~N989;
  assign N1182 = reservation_i[388] ^ N1181;
  assign N1183 = reservation_i[387] ^ N1180;
  assign N1184 = reservation_i[386] ^ N1179;
  assign N1185 = reservation_i[385] ^ N1178;
  assign N1186 = reservation_i[384] ^ N1177;
  assign N1187 = reservation_i[383] ^ N1176;
  assign N1188 = reservation_i[382] ^ N1175;
  assign N1189 = reservation_i[381] ^ N1174;
  assign N1190 = reservation_i[380] ^ N1173;
  assign N1191 = reservation_i[379] ^ N1172;
  assign N1192 = reservation_i[378] ^ N1171;
  assign N1193 = reservation_i[377] ^ N1170;
  assign N1194 = reservation_i[376] ^ N1169;
  assign N1195 = reservation_i[375] ^ N1168;
  assign N1196 = reservation_i[374] ^ N1167;
  assign N1197 = reservation_i[373] ^ N1166;
  assign N1198 = reservation_i[372] ^ N1165;
  assign N1199 = reservation_i[371] ^ N1164;
  assign N1200 = reservation_i[370] ^ N1163;
  assign N1201 = reservation_i[369] ^ N1162;
  assign N1202 = reservation_i[368] ^ N1161;
  assign N1203 = reservation_i[367] ^ N1160;
  assign N1204 = reservation_i[366] ^ N1159;
  assign N1205 = reservation_i[365] ^ N1158;
  assign N1206 = reservation_i[364] ^ N1157;
  assign N1207 = reservation_i[363] ^ N1156;
  assign N1208 = reservation_i[362] ^ N1155;
  assign N1209 = reservation_i[361] ^ N1154;
  assign N1210 = reservation_i[360] ^ N1153;
  assign N1211 = reservation_i[359] ^ N1152;
  assign N1212 = reservation_i[358] ^ N1151;
  assign N1213 = reservation_i[357] ^ N1150;
  assign N1214 = reservation_i[356] ^ N1149;
  assign N1215 = reservation_i[355] ^ N1148;
  assign N1216 = reservation_i[354] ^ N1147;
  assign N1217 = reservation_i[353] ^ N1146;
  assign N1218 = reservation_i[352] ^ N1145;
  assign N1219 = reservation_i[351] ^ N1144;
  assign N1220 = reservation_i[350] ^ N1143;
  assign N1221 = reservation_i[349] ^ N1142;
  assign N1222 = reservation_i[348] ^ N1141;
  assign N1223 = reservation_i[347] ^ N1140;
  assign N1224 = reservation_i[346] ^ N1139;
  assign N1225 = reservation_i[345] ^ N1138;
  assign N1226 = reservation_i[344] ^ N1137;
  assign N1227 = reservation_i[343] ^ N1136;
  assign N1228 = reservation_i[342] ^ N1135;
  assign N1229 = reservation_i[341] ^ N1134;
  assign N1230 = reservation_i[340] ^ N1133;
  assign N1231 = reservation_i[339] ^ N1132;
  assign N1232 = reservation_i[338] ^ N1131;
  assign N1233 = reservation_i[337] ^ N1130;
  assign N1234 = reservation_i[336] ^ N1129;
  assign N1235 = reservation_i[335] ^ N1128;
  assign N1236 = reservation_i[334] ^ N1127;
  assign N1237 = reservation_i[333] ^ N1126;
  assign N1238 = reservation_i[332] ^ N1125;
  assign N1239 = reservation_i[331] ^ N1124;
  assign N1240 = reservation_i[330] ^ N1123;
  assign N1241 = reservation_i[329] ^ N1122;
  assign N1242 = reservation_i[328] ^ N1121;
  assign N1243 = reservation_i[327] ^ N1120;
  assign N1244 = reservation_i[326] ^ N1119;
  assign N1245 = reservation_i[325] ^ N1118;
  assign N1310 = reservation_i[388] | N1309;
  assign N1311 = reservation_i[387] | N1308;
  assign N1312 = reservation_i[386] | N1307;
  assign N1313 = reservation_i[385] | N1306;
  assign N1314 = reservation_i[384] | N1305;
  assign N1315 = reservation_i[383] | N1304;
  assign N1316 = reservation_i[382] | N1303;
  assign N1317 = reservation_i[381] | N1302;
  assign N1318 = reservation_i[380] | N1301;
  assign N1319 = reservation_i[379] | N1300;
  assign N1320 = reservation_i[378] | N1299;
  assign N1321 = reservation_i[377] | N1298;
  assign N1322 = reservation_i[376] | N1297;
  assign N1323 = reservation_i[375] | N1296;
  assign N1324 = reservation_i[374] | N1295;
  assign N1325 = reservation_i[373] | N1294;
  assign N1326 = reservation_i[372] | N1293;
  assign N1327 = reservation_i[371] | N1292;
  assign N1328 = reservation_i[370] | N1291;
  assign N1329 = reservation_i[369] | N1290;
  assign N1330 = reservation_i[368] | N1289;
  assign N1331 = reservation_i[367] | N1288;
  assign N1332 = reservation_i[366] | N1287;
  assign N1333 = reservation_i[365] | N1286;
  assign N1334 = reservation_i[364] | N1285;
  assign N1335 = reservation_i[363] | N1284;
  assign N1336 = reservation_i[362] | N1283;
  assign N1337 = reservation_i[361] | N1282;
  assign N1338 = reservation_i[360] | N1281;
  assign N1339 = reservation_i[359] | N1280;
  assign N1340 = reservation_i[358] | N1279;
  assign N1341 = reservation_i[357] | N1278;
  assign N1342 = reservation_i[356] | N1277;
  assign N1343 = reservation_i[355] | N1276;
  assign N1344 = reservation_i[354] | N1275;
  assign N1345 = reservation_i[353] | N1274;
  assign N1346 = reservation_i[352] | N1273;
  assign N1347 = reservation_i[351] | N1272;
  assign N1348 = reservation_i[350] | N1271;
  assign N1349 = reservation_i[349] | N1270;
  assign N1350 = reservation_i[348] | N1269;
  assign N1351 = reservation_i[347] | N1268;
  assign N1352 = reservation_i[346] | N1267;
  assign N1353 = reservation_i[345] | N1266;
  assign N1354 = reservation_i[344] | N1265;
  assign N1355 = reservation_i[343] | N1264;
  assign N1356 = reservation_i[342] | N1263;
  assign N1357 = reservation_i[341] | N1262;
  assign N1358 = reservation_i[340] | N1261;
  assign N1359 = reservation_i[339] | N1260;
  assign N1360 = reservation_i[338] | N1259;
  assign N1361 = reservation_i[337] | N1258;
  assign N1362 = reservation_i[336] | N1257;
  assign N1363 = reservation_i[335] | N1256;
  assign N1364 = reservation_i[334] | N1255;
  assign N1365 = reservation_i[333] | N1254;
  assign N1366 = reservation_i[332] | N1253;
  assign N1367 = reservation_i[331] | N1252;
  assign N1368 = reservation_i[330] | N1251;
  assign N1369 = reservation_i[329] | N1250;
  assign N1370 = reservation_i[328] | N1249;
  assign N1371 = reservation_i[327] | N1248;
  assign N1372 = reservation_i[326] | N1247;
  assign N1373 = reservation_i[325] | N1246;
  assign N1438 = reservation_i[432] | reservation_i[431];
  assign N1439 = ~N1438;
  assign v_o = N1984 & reservation_i[448];
  assign N1984 = en_i & reservation_i[520];
  assign branch_o = N1985 | reservation_i[431];
  assign N1985 = reservation_i[433] | reservation_i[432];
  assign btaken_o = N1987 | reservation_i[431];
  assign N1987 = N1986 | reservation_i[432];
  assign N1986 = reservation_i[433] & comp_result;
  assign N1440 = ~btaken_o;

endmodule



module bsg_dff_width_p521
(
  clk_i,
  data_i,
  data_o
);

  input [520:0] data_i;
  output [520:0] data_o;
  input clk_i;
  wire [520:0] data_o;
  reg data_o_520_sv2v_reg,data_o_519_sv2v_reg,data_o_518_sv2v_reg,data_o_517_sv2v_reg,
  data_o_516_sv2v_reg,data_o_515_sv2v_reg,data_o_514_sv2v_reg,data_o_513_sv2v_reg,
  data_o_512_sv2v_reg,data_o_511_sv2v_reg,data_o_510_sv2v_reg,data_o_509_sv2v_reg,
  data_o_508_sv2v_reg,data_o_507_sv2v_reg,data_o_506_sv2v_reg,data_o_505_sv2v_reg,
  data_o_504_sv2v_reg,data_o_503_sv2v_reg,data_o_502_sv2v_reg,data_o_501_sv2v_reg,
  data_o_500_sv2v_reg,data_o_499_sv2v_reg,data_o_498_sv2v_reg,data_o_497_sv2v_reg,
  data_o_496_sv2v_reg,data_o_495_sv2v_reg,data_o_494_sv2v_reg,data_o_493_sv2v_reg,
  data_o_492_sv2v_reg,data_o_491_sv2v_reg,data_o_490_sv2v_reg,data_o_489_sv2v_reg,
  data_o_488_sv2v_reg,data_o_487_sv2v_reg,data_o_486_sv2v_reg,data_o_485_sv2v_reg,
  data_o_484_sv2v_reg,data_o_483_sv2v_reg,data_o_482_sv2v_reg,data_o_481_sv2v_reg,
  data_o_480_sv2v_reg,data_o_479_sv2v_reg,data_o_478_sv2v_reg,data_o_477_sv2v_reg,
  data_o_476_sv2v_reg,data_o_475_sv2v_reg,data_o_474_sv2v_reg,data_o_473_sv2v_reg,
  data_o_472_sv2v_reg,data_o_471_sv2v_reg,data_o_470_sv2v_reg,data_o_469_sv2v_reg,
  data_o_468_sv2v_reg,data_o_467_sv2v_reg,data_o_466_sv2v_reg,data_o_465_sv2v_reg,
  data_o_464_sv2v_reg,data_o_463_sv2v_reg,data_o_462_sv2v_reg,data_o_461_sv2v_reg,
  data_o_460_sv2v_reg,data_o_459_sv2v_reg,data_o_458_sv2v_reg,data_o_457_sv2v_reg,
  data_o_456_sv2v_reg,data_o_455_sv2v_reg,data_o_454_sv2v_reg,data_o_453_sv2v_reg,
  data_o_452_sv2v_reg,data_o_451_sv2v_reg,data_o_450_sv2v_reg,data_o_449_sv2v_reg,
  data_o_448_sv2v_reg,data_o_447_sv2v_reg,data_o_446_sv2v_reg,data_o_445_sv2v_reg,
  data_o_444_sv2v_reg,data_o_443_sv2v_reg,data_o_442_sv2v_reg,data_o_441_sv2v_reg,
  data_o_440_sv2v_reg,data_o_439_sv2v_reg,data_o_438_sv2v_reg,data_o_437_sv2v_reg,
  data_o_436_sv2v_reg,data_o_435_sv2v_reg,data_o_434_sv2v_reg,data_o_433_sv2v_reg,
  data_o_432_sv2v_reg,data_o_431_sv2v_reg,data_o_430_sv2v_reg,data_o_429_sv2v_reg,
  data_o_428_sv2v_reg,data_o_427_sv2v_reg,data_o_426_sv2v_reg,data_o_425_sv2v_reg,
  data_o_424_sv2v_reg,data_o_423_sv2v_reg,data_o_422_sv2v_reg,data_o_421_sv2v_reg,
  data_o_420_sv2v_reg,data_o_419_sv2v_reg,data_o_418_sv2v_reg,data_o_417_sv2v_reg,
  data_o_416_sv2v_reg,data_o_415_sv2v_reg,data_o_414_sv2v_reg,data_o_413_sv2v_reg,
  data_o_412_sv2v_reg,data_o_411_sv2v_reg,data_o_410_sv2v_reg,data_o_409_sv2v_reg,
  data_o_408_sv2v_reg,data_o_407_sv2v_reg,data_o_406_sv2v_reg,data_o_405_sv2v_reg,
  data_o_404_sv2v_reg,data_o_403_sv2v_reg,data_o_402_sv2v_reg,data_o_401_sv2v_reg,
  data_o_400_sv2v_reg,data_o_399_sv2v_reg,data_o_398_sv2v_reg,data_o_397_sv2v_reg,
  data_o_396_sv2v_reg,data_o_395_sv2v_reg,data_o_394_sv2v_reg,data_o_393_sv2v_reg,
  data_o_392_sv2v_reg,data_o_391_sv2v_reg,data_o_390_sv2v_reg,data_o_389_sv2v_reg,
  data_o_388_sv2v_reg,data_o_387_sv2v_reg,data_o_386_sv2v_reg,data_o_385_sv2v_reg,
  data_o_384_sv2v_reg,data_o_383_sv2v_reg,data_o_382_sv2v_reg,data_o_381_sv2v_reg,
  data_o_380_sv2v_reg,data_o_379_sv2v_reg,data_o_378_sv2v_reg,data_o_377_sv2v_reg,
  data_o_376_sv2v_reg,data_o_375_sv2v_reg,data_o_374_sv2v_reg,data_o_373_sv2v_reg,
  data_o_372_sv2v_reg,data_o_371_sv2v_reg,data_o_370_sv2v_reg,data_o_369_sv2v_reg,
  data_o_368_sv2v_reg,data_o_367_sv2v_reg,data_o_366_sv2v_reg,data_o_365_sv2v_reg,
  data_o_364_sv2v_reg,data_o_363_sv2v_reg,data_o_362_sv2v_reg,data_o_361_sv2v_reg,
  data_o_360_sv2v_reg,data_o_359_sv2v_reg,data_o_358_sv2v_reg,data_o_357_sv2v_reg,
  data_o_356_sv2v_reg,data_o_355_sv2v_reg,data_o_354_sv2v_reg,data_o_353_sv2v_reg,
  data_o_352_sv2v_reg,data_o_351_sv2v_reg,data_o_350_sv2v_reg,data_o_349_sv2v_reg,
  data_o_348_sv2v_reg,data_o_347_sv2v_reg,data_o_346_sv2v_reg,data_o_345_sv2v_reg,
  data_o_344_sv2v_reg,data_o_343_sv2v_reg,data_o_342_sv2v_reg,data_o_341_sv2v_reg,
  data_o_340_sv2v_reg,data_o_339_sv2v_reg,data_o_338_sv2v_reg,data_o_337_sv2v_reg,
  data_o_336_sv2v_reg,data_o_335_sv2v_reg,data_o_334_sv2v_reg,data_o_333_sv2v_reg,
  data_o_332_sv2v_reg,data_o_331_sv2v_reg,data_o_330_sv2v_reg,data_o_329_sv2v_reg,
  data_o_328_sv2v_reg,data_o_327_sv2v_reg,data_o_326_sv2v_reg,data_o_325_sv2v_reg,
  data_o_324_sv2v_reg,data_o_323_sv2v_reg,data_o_322_sv2v_reg,data_o_321_sv2v_reg,
  data_o_320_sv2v_reg,data_o_319_sv2v_reg,data_o_318_sv2v_reg,data_o_317_sv2v_reg,
  data_o_316_sv2v_reg,data_o_315_sv2v_reg,data_o_314_sv2v_reg,data_o_313_sv2v_reg,
  data_o_312_sv2v_reg,data_o_311_sv2v_reg,data_o_310_sv2v_reg,data_o_309_sv2v_reg,
  data_o_308_sv2v_reg,data_o_307_sv2v_reg,data_o_306_sv2v_reg,data_o_305_sv2v_reg,
  data_o_304_sv2v_reg,data_o_303_sv2v_reg,data_o_302_sv2v_reg,data_o_301_sv2v_reg,
  data_o_300_sv2v_reg,data_o_299_sv2v_reg,data_o_298_sv2v_reg,data_o_297_sv2v_reg,
  data_o_296_sv2v_reg,data_o_295_sv2v_reg,data_o_294_sv2v_reg,data_o_293_sv2v_reg,
  data_o_292_sv2v_reg,data_o_291_sv2v_reg,data_o_290_sv2v_reg,data_o_289_sv2v_reg,
  data_o_288_sv2v_reg,data_o_287_sv2v_reg,data_o_286_sv2v_reg,data_o_285_sv2v_reg,
  data_o_284_sv2v_reg,data_o_283_sv2v_reg,data_o_282_sv2v_reg,data_o_281_sv2v_reg,
  data_o_280_sv2v_reg,data_o_279_sv2v_reg,data_o_278_sv2v_reg,data_o_277_sv2v_reg,
  data_o_276_sv2v_reg,data_o_275_sv2v_reg,data_o_274_sv2v_reg,data_o_273_sv2v_reg,
  data_o_272_sv2v_reg,data_o_271_sv2v_reg,data_o_270_sv2v_reg,data_o_269_sv2v_reg,
  data_o_268_sv2v_reg,data_o_267_sv2v_reg,data_o_266_sv2v_reg,data_o_265_sv2v_reg,
  data_o_264_sv2v_reg,data_o_263_sv2v_reg,data_o_262_sv2v_reg,data_o_261_sv2v_reg,
  data_o_260_sv2v_reg,data_o_259_sv2v_reg,data_o_258_sv2v_reg,data_o_257_sv2v_reg,
  data_o_256_sv2v_reg,data_o_255_sv2v_reg,data_o_254_sv2v_reg,data_o_253_sv2v_reg,
  data_o_252_sv2v_reg,data_o_251_sv2v_reg,data_o_250_sv2v_reg,data_o_249_sv2v_reg,
  data_o_248_sv2v_reg,data_o_247_sv2v_reg,data_o_246_sv2v_reg,data_o_245_sv2v_reg,
  data_o_244_sv2v_reg,data_o_243_sv2v_reg,data_o_242_sv2v_reg,data_o_241_sv2v_reg,
  data_o_240_sv2v_reg,data_o_239_sv2v_reg,data_o_238_sv2v_reg,data_o_237_sv2v_reg,
  data_o_236_sv2v_reg,data_o_235_sv2v_reg,data_o_234_sv2v_reg,data_o_233_sv2v_reg,
  data_o_232_sv2v_reg,data_o_231_sv2v_reg,data_o_230_sv2v_reg,data_o_229_sv2v_reg,
  data_o_228_sv2v_reg,data_o_227_sv2v_reg,data_o_226_sv2v_reg,data_o_225_sv2v_reg,
  data_o_224_sv2v_reg,data_o_223_sv2v_reg,data_o_222_sv2v_reg,data_o_221_sv2v_reg,
  data_o_220_sv2v_reg,data_o_219_sv2v_reg,data_o_218_sv2v_reg,data_o_217_sv2v_reg,
  data_o_216_sv2v_reg,data_o_215_sv2v_reg,data_o_214_sv2v_reg,data_o_213_sv2v_reg,
  data_o_212_sv2v_reg,data_o_211_sv2v_reg,data_o_210_sv2v_reg,data_o_209_sv2v_reg,
  data_o_208_sv2v_reg,data_o_207_sv2v_reg,data_o_206_sv2v_reg,data_o_205_sv2v_reg,
  data_o_204_sv2v_reg,data_o_203_sv2v_reg,data_o_202_sv2v_reg,data_o_201_sv2v_reg,
  data_o_200_sv2v_reg,data_o_199_sv2v_reg,data_o_198_sv2v_reg,data_o_197_sv2v_reg,
  data_o_196_sv2v_reg,data_o_195_sv2v_reg,data_o_194_sv2v_reg,data_o_193_sv2v_reg,
  data_o_192_sv2v_reg,data_o_191_sv2v_reg,data_o_190_sv2v_reg,data_o_189_sv2v_reg,
  data_o_188_sv2v_reg,data_o_187_sv2v_reg,data_o_186_sv2v_reg,data_o_185_sv2v_reg,
  data_o_184_sv2v_reg,data_o_183_sv2v_reg,data_o_182_sv2v_reg,data_o_181_sv2v_reg,
  data_o_180_sv2v_reg,data_o_179_sv2v_reg,data_o_178_sv2v_reg,data_o_177_sv2v_reg,
  data_o_176_sv2v_reg,data_o_175_sv2v_reg,data_o_174_sv2v_reg,data_o_173_sv2v_reg,
  data_o_172_sv2v_reg,data_o_171_sv2v_reg,data_o_170_sv2v_reg,data_o_169_sv2v_reg,
  data_o_168_sv2v_reg,data_o_167_sv2v_reg,data_o_166_sv2v_reg,data_o_165_sv2v_reg,
  data_o_164_sv2v_reg,data_o_163_sv2v_reg,data_o_162_sv2v_reg,data_o_161_sv2v_reg,
  data_o_160_sv2v_reg,data_o_159_sv2v_reg,data_o_158_sv2v_reg,data_o_157_sv2v_reg,
  data_o_156_sv2v_reg,data_o_155_sv2v_reg,data_o_154_sv2v_reg,data_o_153_sv2v_reg,
  data_o_152_sv2v_reg,data_o_151_sv2v_reg,data_o_150_sv2v_reg,data_o_149_sv2v_reg,
  data_o_148_sv2v_reg,data_o_147_sv2v_reg,data_o_146_sv2v_reg,data_o_145_sv2v_reg,
  data_o_144_sv2v_reg,data_o_143_sv2v_reg,data_o_142_sv2v_reg,data_o_141_sv2v_reg,
  data_o_140_sv2v_reg,data_o_139_sv2v_reg,data_o_138_sv2v_reg,data_o_137_sv2v_reg,
  data_o_136_sv2v_reg,data_o_135_sv2v_reg,data_o_134_sv2v_reg,data_o_133_sv2v_reg,
  data_o_132_sv2v_reg,data_o_131_sv2v_reg,data_o_130_sv2v_reg,data_o_129_sv2v_reg,
  data_o_128_sv2v_reg,data_o_127_sv2v_reg,data_o_126_sv2v_reg,data_o_125_sv2v_reg,
  data_o_124_sv2v_reg,data_o_123_sv2v_reg,data_o_122_sv2v_reg,data_o_121_sv2v_reg,
  data_o_120_sv2v_reg,data_o_119_sv2v_reg,data_o_118_sv2v_reg,data_o_117_sv2v_reg,
  data_o_116_sv2v_reg,data_o_115_sv2v_reg,data_o_114_sv2v_reg,data_o_113_sv2v_reg,
  data_o_112_sv2v_reg,data_o_111_sv2v_reg,data_o_110_sv2v_reg,data_o_109_sv2v_reg,
  data_o_108_sv2v_reg,data_o_107_sv2v_reg,data_o_106_sv2v_reg,data_o_105_sv2v_reg,
  data_o_104_sv2v_reg,data_o_103_sv2v_reg,data_o_102_sv2v_reg,data_o_101_sv2v_reg,
  data_o_100_sv2v_reg,data_o_99_sv2v_reg,data_o_98_sv2v_reg,data_o_97_sv2v_reg,
  data_o_96_sv2v_reg,data_o_95_sv2v_reg,data_o_94_sv2v_reg,data_o_93_sv2v_reg,
  data_o_92_sv2v_reg,data_o_91_sv2v_reg,data_o_90_sv2v_reg,data_o_89_sv2v_reg,
  data_o_88_sv2v_reg,data_o_87_sv2v_reg,data_o_86_sv2v_reg,data_o_85_sv2v_reg,
  data_o_84_sv2v_reg,data_o_83_sv2v_reg,data_o_82_sv2v_reg,data_o_81_sv2v_reg,data_o_80_sv2v_reg,
  data_o_79_sv2v_reg,data_o_78_sv2v_reg,data_o_77_sv2v_reg,data_o_76_sv2v_reg,
  data_o_75_sv2v_reg,data_o_74_sv2v_reg,data_o_73_sv2v_reg,data_o_72_sv2v_reg,
  data_o_71_sv2v_reg,data_o_70_sv2v_reg,data_o_69_sv2v_reg,data_o_68_sv2v_reg,
  data_o_67_sv2v_reg,data_o_66_sv2v_reg,data_o_65_sv2v_reg,data_o_64_sv2v_reg,
  data_o_63_sv2v_reg,data_o_62_sv2v_reg,data_o_61_sv2v_reg,data_o_60_sv2v_reg,data_o_59_sv2v_reg,
  data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,data_o_55_sv2v_reg,
  data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,data_o_51_sv2v_reg,
  data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,data_o_47_sv2v_reg,
  data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,data_o_43_sv2v_reg,
  data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,
  data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,
  data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,
  data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,
  data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,
  data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,
  data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,
  data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,
  data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[520] = data_o_520_sv2v_reg;
  assign data_o[519] = data_o_519_sv2v_reg;
  assign data_o[518] = data_o_518_sv2v_reg;
  assign data_o[517] = data_o_517_sv2v_reg;
  assign data_o[516] = data_o_516_sv2v_reg;
  assign data_o[515] = data_o_515_sv2v_reg;
  assign data_o[514] = data_o_514_sv2v_reg;
  assign data_o[513] = data_o_513_sv2v_reg;
  assign data_o[512] = data_o_512_sv2v_reg;
  assign data_o[511] = data_o_511_sv2v_reg;
  assign data_o[510] = data_o_510_sv2v_reg;
  assign data_o[509] = data_o_509_sv2v_reg;
  assign data_o[508] = data_o_508_sv2v_reg;
  assign data_o[507] = data_o_507_sv2v_reg;
  assign data_o[506] = data_o_506_sv2v_reg;
  assign data_o[505] = data_o_505_sv2v_reg;
  assign data_o[504] = data_o_504_sv2v_reg;
  assign data_o[503] = data_o_503_sv2v_reg;
  assign data_o[502] = data_o_502_sv2v_reg;
  assign data_o[501] = data_o_501_sv2v_reg;
  assign data_o[500] = data_o_500_sv2v_reg;
  assign data_o[499] = data_o_499_sv2v_reg;
  assign data_o[498] = data_o_498_sv2v_reg;
  assign data_o[497] = data_o_497_sv2v_reg;
  assign data_o[496] = data_o_496_sv2v_reg;
  assign data_o[495] = data_o_495_sv2v_reg;
  assign data_o[494] = data_o_494_sv2v_reg;
  assign data_o[493] = data_o_493_sv2v_reg;
  assign data_o[492] = data_o_492_sv2v_reg;
  assign data_o[491] = data_o_491_sv2v_reg;
  assign data_o[490] = data_o_490_sv2v_reg;
  assign data_o[489] = data_o_489_sv2v_reg;
  assign data_o[488] = data_o_488_sv2v_reg;
  assign data_o[487] = data_o_487_sv2v_reg;
  assign data_o[486] = data_o_486_sv2v_reg;
  assign data_o[485] = data_o_485_sv2v_reg;
  assign data_o[484] = data_o_484_sv2v_reg;
  assign data_o[483] = data_o_483_sv2v_reg;
  assign data_o[482] = data_o_482_sv2v_reg;
  assign data_o[481] = data_o_481_sv2v_reg;
  assign data_o[480] = data_o_480_sv2v_reg;
  assign data_o[479] = data_o_479_sv2v_reg;
  assign data_o[478] = data_o_478_sv2v_reg;
  assign data_o[477] = data_o_477_sv2v_reg;
  assign data_o[476] = data_o_476_sv2v_reg;
  assign data_o[475] = data_o_475_sv2v_reg;
  assign data_o[474] = data_o_474_sv2v_reg;
  assign data_o[473] = data_o_473_sv2v_reg;
  assign data_o[472] = data_o_472_sv2v_reg;
  assign data_o[471] = data_o_471_sv2v_reg;
  assign data_o[470] = data_o_470_sv2v_reg;
  assign data_o[469] = data_o_469_sv2v_reg;
  assign data_o[468] = data_o_468_sv2v_reg;
  assign data_o[467] = data_o_467_sv2v_reg;
  assign data_o[466] = data_o_466_sv2v_reg;
  assign data_o[465] = data_o_465_sv2v_reg;
  assign data_o[464] = data_o_464_sv2v_reg;
  assign data_o[463] = data_o_463_sv2v_reg;
  assign data_o[462] = data_o_462_sv2v_reg;
  assign data_o[461] = data_o_461_sv2v_reg;
  assign data_o[460] = data_o_460_sv2v_reg;
  assign data_o[459] = data_o_459_sv2v_reg;
  assign data_o[458] = data_o_458_sv2v_reg;
  assign data_o[457] = data_o_457_sv2v_reg;
  assign data_o[456] = data_o_456_sv2v_reg;
  assign data_o[455] = data_o_455_sv2v_reg;
  assign data_o[454] = data_o_454_sv2v_reg;
  assign data_o[453] = data_o_453_sv2v_reg;
  assign data_o[452] = data_o_452_sv2v_reg;
  assign data_o[451] = data_o_451_sv2v_reg;
  assign data_o[450] = data_o_450_sv2v_reg;
  assign data_o[449] = data_o_449_sv2v_reg;
  assign data_o[448] = data_o_448_sv2v_reg;
  assign data_o[447] = data_o_447_sv2v_reg;
  assign data_o[446] = data_o_446_sv2v_reg;
  assign data_o[445] = data_o_445_sv2v_reg;
  assign data_o[444] = data_o_444_sv2v_reg;
  assign data_o[443] = data_o_443_sv2v_reg;
  assign data_o[442] = data_o_442_sv2v_reg;
  assign data_o[441] = data_o_441_sv2v_reg;
  assign data_o[440] = data_o_440_sv2v_reg;
  assign data_o[439] = data_o_439_sv2v_reg;
  assign data_o[438] = data_o_438_sv2v_reg;
  assign data_o[437] = data_o_437_sv2v_reg;
  assign data_o[436] = data_o_436_sv2v_reg;
  assign data_o[435] = data_o_435_sv2v_reg;
  assign data_o[434] = data_o_434_sv2v_reg;
  assign data_o[433] = data_o_433_sv2v_reg;
  assign data_o[432] = data_o_432_sv2v_reg;
  assign data_o[431] = data_o_431_sv2v_reg;
  assign data_o[430] = data_o_430_sv2v_reg;
  assign data_o[429] = data_o_429_sv2v_reg;
  assign data_o[428] = data_o_428_sv2v_reg;
  assign data_o[427] = data_o_427_sv2v_reg;
  assign data_o[426] = data_o_426_sv2v_reg;
  assign data_o[425] = data_o_425_sv2v_reg;
  assign data_o[424] = data_o_424_sv2v_reg;
  assign data_o[423] = data_o_423_sv2v_reg;
  assign data_o[422] = data_o_422_sv2v_reg;
  assign data_o[421] = data_o_421_sv2v_reg;
  assign data_o[420] = data_o_420_sv2v_reg;
  assign data_o[419] = data_o_419_sv2v_reg;
  assign data_o[418] = data_o_418_sv2v_reg;
  assign data_o[417] = data_o_417_sv2v_reg;
  assign data_o[416] = data_o_416_sv2v_reg;
  assign data_o[415] = data_o_415_sv2v_reg;
  assign data_o[414] = data_o_414_sv2v_reg;
  assign data_o[413] = data_o_413_sv2v_reg;
  assign data_o[412] = data_o_412_sv2v_reg;
  assign data_o[411] = data_o_411_sv2v_reg;
  assign data_o[410] = data_o_410_sv2v_reg;
  assign data_o[409] = data_o_409_sv2v_reg;
  assign data_o[408] = data_o_408_sv2v_reg;
  assign data_o[407] = data_o_407_sv2v_reg;
  assign data_o[406] = data_o_406_sv2v_reg;
  assign data_o[405] = data_o_405_sv2v_reg;
  assign data_o[404] = data_o_404_sv2v_reg;
  assign data_o[403] = data_o_403_sv2v_reg;
  assign data_o[402] = data_o_402_sv2v_reg;
  assign data_o[401] = data_o_401_sv2v_reg;
  assign data_o[400] = data_o_400_sv2v_reg;
  assign data_o[399] = data_o_399_sv2v_reg;
  assign data_o[398] = data_o_398_sv2v_reg;
  assign data_o[397] = data_o_397_sv2v_reg;
  assign data_o[396] = data_o_396_sv2v_reg;
  assign data_o[395] = data_o_395_sv2v_reg;
  assign data_o[394] = data_o_394_sv2v_reg;
  assign data_o[393] = data_o_393_sv2v_reg;
  assign data_o[392] = data_o_392_sv2v_reg;
  assign data_o[391] = data_o_391_sv2v_reg;
  assign data_o[390] = data_o_390_sv2v_reg;
  assign data_o[389] = data_o_389_sv2v_reg;
  assign data_o[388] = data_o_388_sv2v_reg;
  assign data_o[387] = data_o_387_sv2v_reg;
  assign data_o[386] = data_o_386_sv2v_reg;
  assign data_o[385] = data_o_385_sv2v_reg;
  assign data_o[384] = data_o_384_sv2v_reg;
  assign data_o[383] = data_o_383_sv2v_reg;
  assign data_o[382] = data_o_382_sv2v_reg;
  assign data_o[381] = data_o_381_sv2v_reg;
  assign data_o[380] = data_o_380_sv2v_reg;
  assign data_o[379] = data_o_379_sv2v_reg;
  assign data_o[378] = data_o_378_sv2v_reg;
  assign data_o[377] = data_o_377_sv2v_reg;
  assign data_o[376] = data_o_376_sv2v_reg;
  assign data_o[375] = data_o_375_sv2v_reg;
  assign data_o[374] = data_o_374_sv2v_reg;
  assign data_o[373] = data_o_373_sv2v_reg;
  assign data_o[372] = data_o_372_sv2v_reg;
  assign data_o[371] = data_o_371_sv2v_reg;
  assign data_o[370] = data_o_370_sv2v_reg;
  assign data_o[369] = data_o_369_sv2v_reg;
  assign data_o[368] = data_o_368_sv2v_reg;
  assign data_o[367] = data_o_367_sv2v_reg;
  assign data_o[366] = data_o_366_sv2v_reg;
  assign data_o[365] = data_o_365_sv2v_reg;
  assign data_o[364] = data_o_364_sv2v_reg;
  assign data_o[363] = data_o_363_sv2v_reg;
  assign data_o[362] = data_o_362_sv2v_reg;
  assign data_o[361] = data_o_361_sv2v_reg;
  assign data_o[360] = data_o_360_sv2v_reg;
  assign data_o[359] = data_o_359_sv2v_reg;
  assign data_o[358] = data_o_358_sv2v_reg;
  assign data_o[357] = data_o_357_sv2v_reg;
  assign data_o[356] = data_o_356_sv2v_reg;
  assign data_o[355] = data_o_355_sv2v_reg;
  assign data_o[354] = data_o_354_sv2v_reg;
  assign data_o[353] = data_o_353_sv2v_reg;
  assign data_o[352] = data_o_352_sv2v_reg;
  assign data_o[351] = data_o_351_sv2v_reg;
  assign data_o[350] = data_o_350_sv2v_reg;
  assign data_o[349] = data_o_349_sv2v_reg;
  assign data_o[348] = data_o_348_sv2v_reg;
  assign data_o[347] = data_o_347_sv2v_reg;
  assign data_o[346] = data_o_346_sv2v_reg;
  assign data_o[345] = data_o_345_sv2v_reg;
  assign data_o[344] = data_o_344_sv2v_reg;
  assign data_o[343] = data_o_343_sv2v_reg;
  assign data_o[342] = data_o_342_sv2v_reg;
  assign data_o[341] = data_o_341_sv2v_reg;
  assign data_o[340] = data_o_340_sv2v_reg;
  assign data_o[339] = data_o_339_sv2v_reg;
  assign data_o[338] = data_o_338_sv2v_reg;
  assign data_o[337] = data_o_337_sv2v_reg;
  assign data_o[336] = data_o_336_sv2v_reg;
  assign data_o[335] = data_o_335_sv2v_reg;
  assign data_o[334] = data_o_334_sv2v_reg;
  assign data_o[333] = data_o_333_sv2v_reg;
  assign data_o[332] = data_o_332_sv2v_reg;
  assign data_o[331] = data_o_331_sv2v_reg;
  assign data_o[330] = data_o_330_sv2v_reg;
  assign data_o[329] = data_o_329_sv2v_reg;
  assign data_o[328] = data_o_328_sv2v_reg;
  assign data_o[327] = data_o_327_sv2v_reg;
  assign data_o[326] = data_o_326_sv2v_reg;
  assign data_o[325] = data_o_325_sv2v_reg;
  assign data_o[324] = data_o_324_sv2v_reg;
  assign data_o[323] = data_o_323_sv2v_reg;
  assign data_o[322] = data_o_322_sv2v_reg;
  assign data_o[321] = data_o_321_sv2v_reg;
  assign data_o[320] = data_o_320_sv2v_reg;
  assign data_o[319] = data_o_319_sv2v_reg;
  assign data_o[318] = data_o_318_sv2v_reg;
  assign data_o[317] = data_o_317_sv2v_reg;
  assign data_o[316] = data_o_316_sv2v_reg;
  assign data_o[315] = data_o_315_sv2v_reg;
  assign data_o[314] = data_o_314_sv2v_reg;
  assign data_o[313] = data_o_313_sv2v_reg;
  assign data_o[312] = data_o_312_sv2v_reg;
  assign data_o[311] = data_o_311_sv2v_reg;
  assign data_o[310] = data_o_310_sv2v_reg;
  assign data_o[309] = data_o_309_sv2v_reg;
  assign data_o[308] = data_o_308_sv2v_reg;
  assign data_o[307] = data_o_307_sv2v_reg;
  assign data_o[306] = data_o_306_sv2v_reg;
  assign data_o[305] = data_o_305_sv2v_reg;
  assign data_o[304] = data_o_304_sv2v_reg;
  assign data_o[303] = data_o_303_sv2v_reg;
  assign data_o[302] = data_o_302_sv2v_reg;
  assign data_o[301] = data_o_301_sv2v_reg;
  assign data_o[300] = data_o_300_sv2v_reg;
  assign data_o[299] = data_o_299_sv2v_reg;
  assign data_o[298] = data_o_298_sv2v_reg;
  assign data_o[297] = data_o_297_sv2v_reg;
  assign data_o[296] = data_o_296_sv2v_reg;
  assign data_o[295] = data_o_295_sv2v_reg;
  assign data_o[294] = data_o_294_sv2v_reg;
  assign data_o[293] = data_o_293_sv2v_reg;
  assign data_o[292] = data_o_292_sv2v_reg;
  assign data_o[291] = data_o_291_sv2v_reg;
  assign data_o[290] = data_o_290_sv2v_reg;
  assign data_o[289] = data_o_289_sv2v_reg;
  assign data_o[288] = data_o_288_sv2v_reg;
  assign data_o[287] = data_o_287_sv2v_reg;
  assign data_o[286] = data_o_286_sv2v_reg;
  assign data_o[285] = data_o_285_sv2v_reg;
  assign data_o[284] = data_o_284_sv2v_reg;
  assign data_o[283] = data_o_283_sv2v_reg;
  assign data_o[282] = data_o_282_sv2v_reg;
  assign data_o[281] = data_o_281_sv2v_reg;
  assign data_o[280] = data_o_280_sv2v_reg;
  assign data_o[279] = data_o_279_sv2v_reg;
  assign data_o[278] = data_o_278_sv2v_reg;
  assign data_o[277] = data_o_277_sv2v_reg;
  assign data_o[276] = data_o_276_sv2v_reg;
  assign data_o[275] = data_o_275_sv2v_reg;
  assign data_o[274] = data_o_274_sv2v_reg;
  assign data_o[273] = data_o_273_sv2v_reg;
  assign data_o[272] = data_o_272_sv2v_reg;
  assign data_o[271] = data_o_271_sv2v_reg;
  assign data_o[270] = data_o_270_sv2v_reg;
  assign data_o[269] = data_o_269_sv2v_reg;
  assign data_o[268] = data_o_268_sv2v_reg;
  assign data_o[267] = data_o_267_sv2v_reg;
  assign data_o[266] = data_o_266_sv2v_reg;
  assign data_o[265] = data_o_265_sv2v_reg;
  assign data_o[264] = data_o_264_sv2v_reg;
  assign data_o[263] = data_o_263_sv2v_reg;
  assign data_o[262] = data_o_262_sv2v_reg;
  assign data_o[261] = data_o_261_sv2v_reg;
  assign data_o[260] = data_o_260_sv2v_reg;
  assign data_o[259] = data_o_259_sv2v_reg;
  assign data_o[258] = data_o_258_sv2v_reg;
  assign data_o[257] = data_o_257_sv2v_reg;
  assign data_o[256] = data_o_256_sv2v_reg;
  assign data_o[255] = data_o_255_sv2v_reg;
  assign data_o[254] = data_o_254_sv2v_reg;
  assign data_o[253] = data_o_253_sv2v_reg;
  assign data_o[252] = data_o_252_sv2v_reg;
  assign data_o[251] = data_o_251_sv2v_reg;
  assign data_o[250] = data_o_250_sv2v_reg;
  assign data_o[249] = data_o_249_sv2v_reg;
  assign data_o[248] = data_o_248_sv2v_reg;
  assign data_o[247] = data_o_247_sv2v_reg;
  assign data_o[246] = data_o_246_sv2v_reg;
  assign data_o[245] = data_o_245_sv2v_reg;
  assign data_o[244] = data_o_244_sv2v_reg;
  assign data_o[243] = data_o_243_sv2v_reg;
  assign data_o[242] = data_o_242_sv2v_reg;
  assign data_o[241] = data_o_241_sv2v_reg;
  assign data_o[240] = data_o_240_sv2v_reg;
  assign data_o[239] = data_o_239_sv2v_reg;
  assign data_o[238] = data_o_238_sv2v_reg;
  assign data_o[237] = data_o_237_sv2v_reg;
  assign data_o[236] = data_o_236_sv2v_reg;
  assign data_o[235] = data_o_235_sv2v_reg;
  assign data_o[234] = data_o_234_sv2v_reg;
  assign data_o[233] = data_o_233_sv2v_reg;
  assign data_o[232] = data_o_232_sv2v_reg;
  assign data_o[231] = data_o_231_sv2v_reg;
  assign data_o[230] = data_o_230_sv2v_reg;
  assign data_o[229] = data_o_229_sv2v_reg;
  assign data_o[228] = data_o_228_sv2v_reg;
  assign data_o[227] = data_o_227_sv2v_reg;
  assign data_o[226] = data_o_226_sv2v_reg;
  assign data_o[225] = data_o_225_sv2v_reg;
  assign data_o[224] = data_o_224_sv2v_reg;
  assign data_o[223] = data_o_223_sv2v_reg;
  assign data_o[222] = data_o_222_sv2v_reg;
  assign data_o[221] = data_o_221_sv2v_reg;
  assign data_o[220] = data_o_220_sv2v_reg;
  assign data_o[219] = data_o_219_sv2v_reg;
  assign data_o[218] = data_o_218_sv2v_reg;
  assign data_o[217] = data_o_217_sv2v_reg;
  assign data_o[216] = data_o_216_sv2v_reg;
  assign data_o[215] = data_o_215_sv2v_reg;
  assign data_o[214] = data_o_214_sv2v_reg;
  assign data_o[213] = data_o_213_sv2v_reg;
  assign data_o[212] = data_o_212_sv2v_reg;
  assign data_o[211] = data_o_211_sv2v_reg;
  assign data_o[210] = data_o_210_sv2v_reg;
  assign data_o[209] = data_o_209_sv2v_reg;
  assign data_o[208] = data_o_208_sv2v_reg;
  assign data_o[207] = data_o_207_sv2v_reg;
  assign data_o[206] = data_o_206_sv2v_reg;
  assign data_o[205] = data_o_205_sv2v_reg;
  assign data_o[204] = data_o_204_sv2v_reg;
  assign data_o[203] = data_o_203_sv2v_reg;
  assign data_o[202] = data_o_202_sv2v_reg;
  assign data_o[201] = data_o_201_sv2v_reg;
  assign data_o[200] = data_o_200_sv2v_reg;
  assign data_o[199] = data_o_199_sv2v_reg;
  assign data_o[198] = data_o_198_sv2v_reg;
  assign data_o[197] = data_o_197_sv2v_reg;
  assign data_o[196] = data_o_196_sv2v_reg;
  assign data_o[195] = data_o_195_sv2v_reg;
  assign data_o[194] = data_o_194_sv2v_reg;
  assign data_o[193] = data_o_193_sv2v_reg;
  assign data_o[192] = data_o_192_sv2v_reg;
  assign data_o[191] = data_o_191_sv2v_reg;
  assign data_o[190] = data_o_190_sv2v_reg;
  assign data_o[189] = data_o_189_sv2v_reg;
  assign data_o[188] = data_o_188_sv2v_reg;
  assign data_o[187] = data_o_187_sv2v_reg;
  assign data_o[186] = data_o_186_sv2v_reg;
  assign data_o[185] = data_o_185_sv2v_reg;
  assign data_o[184] = data_o_184_sv2v_reg;
  assign data_o[183] = data_o_183_sv2v_reg;
  assign data_o[182] = data_o_182_sv2v_reg;
  assign data_o[181] = data_o_181_sv2v_reg;
  assign data_o[180] = data_o_180_sv2v_reg;
  assign data_o[179] = data_o_179_sv2v_reg;
  assign data_o[178] = data_o_178_sv2v_reg;
  assign data_o[177] = data_o_177_sv2v_reg;
  assign data_o[176] = data_o_176_sv2v_reg;
  assign data_o[175] = data_o_175_sv2v_reg;
  assign data_o[174] = data_o_174_sv2v_reg;
  assign data_o[173] = data_o_173_sv2v_reg;
  assign data_o[172] = data_o_172_sv2v_reg;
  assign data_o[171] = data_o_171_sv2v_reg;
  assign data_o[170] = data_o_170_sv2v_reg;
  assign data_o[169] = data_o_169_sv2v_reg;
  assign data_o[168] = data_o_168_sv2v_reg;
  assign data_o[167] = data_o_167_sv2v_reg;
  assign data_o[166] = data_o_166_sv2v_reg;
  assign data_o[165] = data_o_165_sv2v_reg;
  assign data_o[164] = data_o_164_sv2v_reg;
  assign data_o[163] = data_o_163_sv2v_reg;
  assign data_o[162] = data_o_162_sv2v_reg;
  assign data_o[161] = data_o_161_sv2v_reg;
  assign data_o[160] = data_o_160_sv2v_reg;
  assign data_o[159] = data_o_159_sv2v_reg;
  assign data_o[158] = data_o_158_sv2v_reg;
  assign data_o[157] = data_o_157_sv2v_reg;
  assign data_o[156] = data_o_156_sv2v_reg;
  assign data_o[155] = data_o_155_sv2v_reg;
  assign data_o[154] = data_o_154_sv2v_reg;
  assign data_o[153] = data_o_153_sv2v_reg;
  assign data_o[152] = data_o_152_sv2v_reg;
  assign data_o[151] = data_o_151_sv2v_reg;
  assign data_o[150] = data_o_150_sv2v_reg;
  assign data_o[149] = data_o_149_sv2v_reg;
  assign data_o[148] = data_o_148_sv2v_reg;
  assign data_o[147] = data_o_147_sv2v_reg;
  assign data_o[146] = data_o_146_sv2v_reg;
  assign data_o[145] = data_o_145_sv2v_reg;
  assign data_o[144] = data_o_144_sv2v_reg;
  assign data_o[143] = data_o_143_sv2v_reg;
  assign data_o[142] = data_o_142_sv2v_reg;
  assign data_o[141] = data_o_141_sv2v_reg;
  assign data_o[140] = data_o_140_sv2v_reg;
  assign data_o[139] = data_o_139_sv2v_reg;
  assign data_o[138] = data_o_138_sv2v_reg;
  assign data_o[137] = data_o_137_sv2v_reg;
  assign data_o[136] = data_o_136_sv2v_reg;
  assign data_o[135] = data_o_135_sv2v_reg;
  assign data_o[134] = data_o_134_sv2v_reg;
  assign data_o[133] = data_o_133_sv2v_reg;
  assign data_o[132] = data_o_132_sv2v_reg;
  assign data_o[131] = data_o_131_sv2v_reg;
  assign data_o[130] = data_o_130_sv2v_reg;
  assign data_o[129] = data_o_129_sv2v_reg;
  assign data_o[128] = data_o_128_sv2v_reg;
  assign data_o[127] = data_o_127_sv2v_reg;
  assign data_o[126] = data_o_126_sv2v_reg;
  assign data_o[125] = data_o_125_sv2v_reg;
  assign data_o[124] = data_o_124_sv2v_reg;
  assign data_o[123] = data_o_123_sv2v_reg;
  assign data_o[122] = data_o_122_sv2v_reg;
  assign data_o[121] = data_o_121_sv2v_reg;
  assign data_o[120] = data_o_120_sv2v_reg;
  assign data_o[119] = data_o_119_sv2v_reg;
  assign data_o[118] = data_o_118_sv2v_reg;
  assign data_o[117] = data_o_117_sv2v_reg;
  assign data_o[116] = data_o_116_sv2v_reg;
  assign data_o[115] = data_o_115_sv2v_reg;
  assign data_o[114] = data_o_114_sv2v_reg;
  assign data_o[113] = data_o_113_sv2v_reg;
  assign data_o[112] = data_o_112_sv2v_reg;
  assign data_o[111] = data_o_111_sv2v_reg;
  assign data_o[110] = data_o_110_sv2v_reg;
  assign data_o[109] = data_o_109_sv2v_reg;
  assign data_o[108] = data_o_108_sv2v_reg;
  assign data_o[107] = data_o_107_sv2v_reg;
  assign data_o[106] = data_o_106_sv2v_reg;
  assign data_o[105] = data_o_105_sv2v_reg;
  assign data_o[104] = data_o_104_sv2v_reg;
  assign data_o[103] = data_o_103_sv2v_reg;
  assign data_o[102] = data_o_102_sv2v_reg;
  assign data_o[101] = data_o_101_sv2v_reg;
  assign data_o[100] = data_o_100_sv2v_reg;
  assign data_o[99] = data_o_99_sv2v_reg;
  assign data_o[98] = data_o_98_sv2v_reg;
  assign data_o[97] = data_o_97_sv2v_reg;
  assign data_o[96] = data_o_96_sv2v_reg;
  assign data_o[95] = data_o_95_sv2v_reg;
  assign data_o[94] = data_o_94_sv2v_reg;
  assign data_o[93] = data_o_93_sv2v_reg;
  assign data_o[92] = data_o_92_sv2v_reg;
  assign data_o[91] = data_o_91_sv2v_reg;
  assign data_o[90] = data_o_90_sv2v_reg;
  assign data_o[89] = data_o_89_sv2v_reg;
  assign data_o[88] = data_o_88_sv2v_reg;
  assign data_o[87] = data_o_87_sv2v_reg;
  assign data_o[86] = data_o_86_sv2v_reg;
  assign data_o[85] = data_o_85_sv2v_reg;
  assign data_o[84] = data_o_84_sv2v_reg;
  assign data_o[83] = data_o_83_sv2v_reg;
  assign data_o[82] = data_o_82_sv2v_reg;
  assign data_o[81] = data_o_81_sv2v_reg;
  assign data_o[80] = data_o_80_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_520_sv2v_reg <= data_i[520];
      data_o_519_sv2v_reg <= data_i[519];
      data_o_518_sv2v_reg <= data_i[518];
      data_o_517_sv2v_reg <= data_i[517];
      data_o_516_sv2v_reg <= data_i[516];
      data_o_515_sv2v_reg <= data_i[515];
      data_o_514_sv2v_reg <= data_i[514];
      data_o_513_sv2v_reg <= data_i[513];
      data_o_512_sv2v_reg <= data_i[512];
      data_o_511_sv2v_reg <= data_i[511];
      data_o_510_sv2v_reg <= data_i[510];
      data_o_509_sv2v_reg <= data_i[509];
      data_o_508_sv2v_reg <= data_i[508];
      data_o_507_sv2v_reg <= data_i[507];
      data_o_506_sv2v_reg <= data_i[506];
      data_o_505_sv2v_reg <= data_i[505];
      data_o_504_sv2v_reg <= data_i[504];
      data_o_503_sv2v_reg <= data_i[503];
      data_o_502_sv2v_reg <= data_i[502];
      data_o_501_sv2v_reg <= data_i[501];
      data_o_500_sv2v_reg <= data_i[500];
      data_o_499_sv2v_reg <= data_i[499];
      data_o_498_sv2v_reg <= data_i[498];
      data_o_497_sv2v_reg <= data_i[497];
      data_o_496_sv2v_reg <= data_i[496];
      data_o_495_sv2v_reg <= data_i[495];
      data_o_494_sv2v_reg <= data_i[494];
      data_o_493_sv2v_reg <= data_i[493];
      data_o_492_sv2v_reg <= data_i[492];
      data_o_491_sv2v_reg <= data_i[491];
      data_o_490_sv2v_reg <= data_i[490];
      data_o_489_sv2v_reg <= data_i[489];
      data_o_488_sv2v_reg <= data_i[488];
      data_o_487_sv2v_reg <= data_i[487];
      data_o_486_sv2v_reg <= data_i[486];
      data_o_485_sv2v_reg <= data_i[485];
      data_o_484_sv2v_reg <= data_i[484];
      data_o_483_sv2v_reg <= data_i[483];
      data_o_482_sv2v_reg <= data_i[482];
      data_o_481_sv2v_reg <= data_i[481];
      data_o_480_sv2v_reg <= data_i[480];
      data_o_479_sv2v_reg <= data_i[479];
      data_o_478_sv2v_reg <= data_i[478];
      data_o_477_sv2v_reg <= data_i[477];
      data_o_476_sv2v_reg <= data_i[476];
      data_o_475_sv2v_reg <= data_i[475];
      data_o_474_sv2v_reg <= data_i[474];
      data_o_473_sv2v_reg <= data_i[473];
      data_o_472_sv2v_reg <= data_i[472];
      data_o_471_sv2v_reg <= data_i[471];
      data_o_470_sv2v_reg <= data_i[470];
      data_o_469_sv2v_reg <= data_i[469];
      data_o_468_sv2v_reg <= data_i[468];
      data_o_467_sv2v_reg <= data_i[467];
      data_o_466_sv2v_reg <= data_i[466];
      data_o_465_sv2v_reg <= data_i[465];
      data_o_464_sv2v_reg <= data_i[464];
      data_o_463_sv2v_reg <= data_i[463];
      data_o_462_sv2v_reg <= data_i[462];
      data_o_461_sv2v_reg <= data_i[461];
      data_o_460_sv2v_reg <= data_i[460];
      data_o_459_sv2v_reg <= data_i[459];
      data_o_458_sv2v_reg <= data_i[458];
      data_o_457_sv2v_reg <= data_i[457];
      data_o_456_sv2v_reg <= data_i[456];
      data_o_455_sv2v_reg <= data_i[455];
      data_o_454_sv2v_reg <= data_i[454];
      data_o_453_sv2v_reg <= data_i[453];
      data_o_452_sv2v_reg <= data_i[452];
      data_o_451_sv2v_reg <= data_i[451];
      data_o_450_sv2v_reg <= data_i[450];
      data_o_449_sv2v_reg <= data_i[449];
      data_o_448_sv2v_reg <= data_i[448];
      data_o_447_sv2v_reg <= data_i[447];
      data_o_446_sv2v_reg <= data_i[446];
      data_o_445_sv2v_reg <= data_i[445];
      data_o_444_sv2v_reg <= data_i[444];
      data_o_443_sv2v_reg <= data_i[443];
      data_o_442_sv2v_reg <= data_i[442];
      data_o_441_sv2v_reg <= data_i[441];
      data_o_440_sv2v_reg <= data_i[440];
      data_o_439_sv2v_reg <= data_i[439];
      data_o_438_sv2v_reg <= data_i[438];
      data_o_437_sv2v_reg <= data_i[437];
      data_o_436_sv2v_reg <= data_i[436];
      data_o_435_sv2v_reg <= data_i[435];
      data_o_434_sv2v_reg <= data_i[434];
      data_o_433_sv2v_reg <= data_i[433];
      data_o_432_sv2v_reg <= data_i[432];
      data_o_431_sv2v_reg <= data_i[431];
      data_o_430_sv2v_reg <= data_i[430];
      data_o_429_sv2v_reg <= data_i[429];
      data_o_428_sv2v_reg <= data_i[428];
      data_o_427_sv2v_reg <= data_i[427];
      data_o_426_sv2v_reg <= data_i[426];
      data_o_425_sv2v_reg <= data_i[425];
      data_o_424_sv2v_reg <= data_i[424];
      data_o_423_sv2v_reg <= data_i[423];
      data_o_422_sv2v_reg <= data_i[422];
      data_o_421_sv2v_reg <= data_i[421];
      data_o_420_sv2v_reg <= data_i[420];
      data_o_419_sv2v_reg <= data_i[419];
      data_o_418_sv2v_reg <= data_i[418];
      data_o_417_sv2v_reg <= data_i[417];
      data_o_416_sv2v_reg <= data_i[416];
      data_o_415_sv2v_reg <= data_i[415];
      data_o_414_sv2v_reg <= data_i[414];
      data_o_413_sv2v_reg <= data_i[413];
      data_o_412_sv2v_reg <= data_i[412];
      data_o_411_sv2v_reg <= data_i[411];
      data_o_410_sv2v_reg <= data_i[410];
      data_o_409_sv2v_reg <= data_i[409];
      data_o_408_sv2v_reg <= data_i[408];
      data_o_407_sv2v_reg <= data_i[407];
      data_o_406_sv2v_reg <= data_i[406];
      data_o_405_sv2v_reg <= data_i[405];
      data_o_404_sv2v_reg <= data_i[404];
      data_o_403_sv2v_reg <= data_i[403];
      data_o_402_sv2v_reg <= data_i[402];
      data_o_401_sv2v_reg <= data_i[401];
      data_o_400_sv2v_reg <= data_i[400];
      data_o_399_sv2v_reg <= data_i[399];
      data_o_398_sv2v_reg <= data_i[398];
      data_o_397_sv2v_reg <= data_i[397];
      data_o_396_sv2v_reg <= data_i[396];
      data_o_395_sv2v_reg <= data_i[395];
      data_o_394_sv2v_reg <= data_i[394];
      data_o_393_sv2v_reg <= data_i[393];
      data_o_392_sv2v_reg <= data_i[392];
      data_o_391_sv2v_reg <= data_i[391];
      data_o_390_sv2v_reg <= data_i[390];
      data_o_389_sv2v_reg <= data_i[389];
      data_o_388_sv2v_reg <= data_i[388];
      data_o_387_sv2v_reg <= data_i[387];
      data_o_386_sv2v_reg <= data_i[386];
      data_o_385_sv2v_reg <= data_i[385];
      data_o_384_sv2v_reg <= data_i[384];
      data_o_383_sv2v_reg <= data_i[383];
      data_o_382_sv2v_reg <= data_i[382];
      data_o_381_sv2v_reg <= data_i[381];
      data_o_380_sv2v_reg <= data_i[380];
      data_o_379_sv2v_reg <= data_i[379];
      data_o_378_sv2v_reg <= data_i[378];
      data_o_377_sv2v_reg <= data_i[377];
      data_o_376_sv2v_reg <= data_i[376];
      data_o_375_sv2v_reg <= data_i[375];
      data_o_374_sv2v_reg <= data_i[374];
      data_o_373_sv2v_reg <= data_i[373];
      data_o_372_sv2v_reg <= data_i[372];
      data_o_371_sv2v_reg <= data_i[371];
      data_o_370_sv2v_reg <= data_i[370];
      data_o_369_sv2v_reg <= data_i[369];
      data_o_368_sv2v_reg <= data_i[368];
      data_o_367_sv2v_reg <= data_i[367];
      data_o_366_sv2v_reg <= data_i[366];
      data_o_365_sv2v_reg <= data_i[365];
      data_o_364_sv2v_reg <= data_i[364];
      data_o_363_sv2v_reg <= data_i[363];
      data_o_362_sv2v_reg <= data_i[362];
      data_o_361_sv2v_reg <= data_i[361];
      data_o_360_sv2v_reg <= data_i[360];
      data_o_359_sv2v_reg <= data_i[359];
      data_o_358_sv2v_reg <= data_i[358];
      data_o_357_sv2v_reg <= data_i[357];
      data_o_356_sv2v_reg <= data_i[356];
      data_o_355_sv2v_reg <= data_i[355];
      data_o_354_sv2v_reg <= data_i[354];
      data_o_353_sv2v_reg <= data_i[353];
      data_o_352_sv2v_reg <= data_i[352];
      data_o_351_sv2v_reg <= data_i[351];
      data_o_350_sv2v_reg <= data_i[350];
      data_o_349_sv2v_reg <= data_i[349];
      data_o_348_sv2v_reg <= data_i[348];
      data_o_347_sv2v_reg <= data_i[347];
      data_o_346_sv2v_reg <= data_i[346];
      data_o_345_sv2v_reg <= data_i[345];
      data_o_344_sv2v_reg <= data_i[344];
      data_o_343_sv2v_reg <= data_i[343];
      data_o_342_sv2v_reg <= data_i[342];
      data_o_341_sv2v_reg <= data_i[341];
      data_o_340_sv2v_reg <= data_i[340];
      data_o_339_sv2v_reg <= data_i[339];
      data_o_338_sv2v_reg <= data_i[338];
      data_o_337_sv2v_reg <= data_i[337];
      data_o_336_sv2v_reg <= data_i[336];
      data_o_335_sv2v_reg <= data_i[335];
      data_o_334_sv2v_reg <= data_i[334];
      data_o_333_sv2v_reg <= data_i[333];
      data_o_332_sv2v_reg <= data_i[332];
      data_o_331_sv2v_reg <= data_i[331];
      data_o_330_sv2v_reg <= data_i[330];
      data_o_329_sv2v_reg <= data_i[329];
      data_o_328_sv2v_reg <= data_i[328];
      data_o_327_sv2v_reg <= data_i[327];
      data_o_326_sv2v_reg <= data_i[326];
      data_o_325_sv2v_reg <= data_i[325];
      data_o_324_sv2v_reg <= data_i[324];
      data_o_323_sv2v_reg <= data_i[323];
      data_o_322_sv2v_reg <= data_i[322];
      data_o_321_sv2v_reg <= data_i[321];
      data_o_320_sv2v_reg <= data_i[320];
      data_o_319_sv2v_reg <= data_i[319];
      data_o_318_sv2v_reg <= data_i[318];
      data_o_317_sv2v_reg <= data_i[317];
      data_o_316_sv2v_reg <= data_i[316];
      data_o_315_sv2v_reg <= data_i[315];
      data_o_314_sv2v_reg <= data_i[314];
      data_o_313_sv2v_reg <= data_i[313];
      data_o_312_sv2v_reg <= data_i[312];
      data_o_311_sv2v_reg <= data_i[311];
      data_o_310_sv2v_reg <= data_i[310];
      data_o_309_sv2v_reg <= data_i[309];
      data_o_308_sv2v_reg <= data_i[308];
      data_o_307_sv2v_reg <= data_i[307];
      data_o_306_sv2v_reg <= data_i[306];
      data_o_305_sv2v_reg <= data_i[305];
      data_o_304_sv2v_reg <= data_i[304];
      data_o_303_sv2v_reg <= data_i[303];
      data_o_302_sv2v_reg <= data_i[302];
      data_o_301_sv2v_reg <= data_i[301];
      data_o_300_sv2v_reg <= data_i[300];
      data_o_299_sv2v_reg <= data_i[299];
      data_o_298_sv2v_reg <= data_i[298];
      data_o_297_sv2v_reg <= data_i[297];
      data_o_296_sv2v_reg <= data_i[296];
      data_o_295_sv2v_reg <= data_i[295];
      data_o_294_sv2v_reg <= data_i[294];
      data_o_293_sv2v_reg <= data_i[293];
      data_o_292_sv2v_reg <= data_i[292];
      data_o_291_sv2v_reg <= data_i[291];
      data_o_290_sv2v_reg <= data_i[290];
      data_o_289_sv2v_reg <= data_i[289];
      data_o_288_sv2v_reg <= data_i[288];
      data_o_287_sv2v_reg <= data_i[287];
      data_o_286_sv2v_reg <= data_i[286];
      data_o_285_sv2v_reg <= data_i[285];
      data_o_284_sv2v_reg <= data_i[284];
      data_o_283_sv2v_reg <= data_i[283];
      data_o_282_sv2v_reg <= data_i[282];
      data_o_281_sv2v_reg <= data_i[281];
      data_o_280_sv2v_reg <= data_i[280];
      data_o_279_sv2v_reg <= data_i[279];
      data_o_278_sv2v_reg <= data_i[278];
      data_o_277_sv2v_reg <= data_i[277];
      data_o_276_sv2v_reg <= data_i[276];
      data_o_275_sv2v_reg <= data_i[275];
      data_o_274_sv2v_reg <= data_i[274];
      data_o_273_sv2v_reg <= data_i[273];
      data_o_272_sv2v_reg <= data_i[272];
      data_o_271_sv2v_reg <= data_i[271];
      data_o_270_sv2v_reg <= data_i[270];
      data_o_269_sv2v_reg <= data_i[269];
      data_o_268_sv2v_reg <= data_i[268];
      data_o_267_sv2v_reg <= data_i[267];
      data_o_266_sv2v_reg <= data_i[266];
      data_o_265_sv2v_reg <= data_i[265];
      data_o_264_sv2v_reg <= data_i[264];
      data_o_263_sv2v_reg <= data_i[263];
      data_o_262_sv2v_reg <= data_i[262];
      data_o_261_sv2v_reg <= data_i[261];
      data_o_260_sv2v_reg <= data_i[260];
      data_o_259_sv2v_reg <= data_i[259];
      data_o_258_sv2v_reg <= data_i[258];
      data_o_257_sv2v_reg <= data_i[257];
      data_o_256_sv2v_reg <= data_i[256];
      data_o_255_sv2v_reg <= data_i[255];
      data_o_254_sv2v_reg <= data_i[254];
      data_o_253_sv2v_reg <= data_i[253];
      data_o_252_sv2v_reg <= data_i[252];
      data_o_251_sv2v_reg <= data_i[251];
      data_o_250_sv2v_reg <= data_i[250];
      data_o_249_sv2v_reg <= data_i[249];
      data_o_248_sv2v_reg <= data_i[248];
      data_o_247_sv2v_reg <= data_i[247];
      data_o_246_sv2v_reg <= data_i[246];
      data_o_245_sv2v_reg <= data_i[245];
      data_o_244_sv2v_reg <= data_i[244];
      data_o_243_sv2v_reg <= data_i[243];
      data_o_242_sv2v_reg <= data_i[242];
      data_o_241_sv2v_reg <= data_i[241];
      data_o_240_sv2v_reg <= data_i[240];
      data_o_239_sv2v_reg <= data_i[239];
      data_o_238_sv2v_reg <= data_i[238];
      data_o_237_sv2v_reg <= data_i[237];
      data_o_236_sv2v_reg <= data_i[236];
      data_o_235_sv2v_reg <= data_i[235];
      data_o_234_sv2v_reg <= data_i[234];
      data_o_233_sv2v_reg <= data_i[233];
      data_o_232_sv2v_reg <= data_i[232];
      data_o_231_sv2v_reg <= data_i[231];
      data_o_230_sv2v_reg <= data_i[230];
      data_o_229_sv2v_reg <= data_i[229];
      data_o_228_sv2v_reg <= data_i[228];
      data_o_227_sv2v_reg <= data_i[227];
      data_o_226_sv2v_reg <= data_i[226];
      data_o_225_sv2v_reg <= data_i[225];
      data_o_224_sv2v_reg <= data_i[224];
      data_o_223_sv2v_reg <= data_i[223];
      data_o_222_sv2v_reg <= data_i[222];
      data_o_221_sv2v_reg <= data_i[221];
      data_o_220_sv2v_reg <= data_i[220];
      data_o_219_sv2v_reg <= data_i[219];
      data_o_218_sv2v_reg <= data_i[218];
      data_o_217_sv2v_reg <= data_i[217];
      data_o_216_sv2v_reg <= data_i[216];
      data_o_215_sv2v_reg <= data_i[215];
      data_o_214_sv2v_reg <= data_i[214];
      data_o_213_sv2v_reg <= data_i[213];
      data_o_212_sv2v_reg <= data_i[212];
      data_o_211_sv2v_reg <= data_i[211];
      data_o_210_sv2v_reg <= data_i[210];
      data_o_209_sv2v_reg <= data_i[209];
      data_o_208_sv2v_reg <= data_i[208];
      data_o_207_sv2v_reg <= data_i[207];
      data_o_206_sv2v_reg <= data_i[206];
      data_o_205_sv2v_reg <= data_i[205];
      data_o_204_sv2v_reg <= data_i[204];
      data_o_203_sv2v_reg <= data_i[203];
      data_o_202_sv2v_reg <= data_i[202];
      data_o_201_sv2v_reg <= data_i[201];
      data_o_200_sv2v_reg <= data_i[200];
      data_o_199_sv2v_reg <= data_i[199];
      data_o_198_sv2v_reg <= data_i[198];
      data_o_197_sv2v_reg <= data_i[197];
      data_o_196_sv2v_reg <= data_i[196];
      data_o_195_sv2v_reg <= data_i[195];
      data_o_194_sv2v_reg <= data_i[194];
      data_o_193_sv2v_reg <= data_i[193];
      data_o_192_sv2v_reg <= data_i[192];
      data_o_191_sv2v_reg <= data_i[191];
      data_o_190_sv2v_reg <= data_i[190];
      data_o_189_sv2v_reg <= data_i[189];
      data_o_188_sv2v_reg <= data_i[188];
      data_o_187_sv2v_reg <= data_i[187];
      data_o_186_sv2v_reg <= data_i[186];
      data_o_185_sv2v_reg <= data_i[185];
      data_o_184_sv2v_reg <= data_i[184];
      data_o_183_sv2v_reg <= data_i[183];
      data_o_182_sv2v_reg <= data_i[182];
      data_o_181_sv2v_reg <= data_i[181];
      data_o_180_sv2v_reg <= data_i[180];
      data_o_179_sv2v_reg <= data_i[179];
      data_o_178_sv2v_reg <= data_i[178];
      data_o_177_sv2v_reg <= data_i[177];
      data_o_176_sv2v_reg <= data_i[176];
      data_o_175_sv2v_reg <= data_i[175];
      data_o_174_sv2v_reg <= data_i[174];
      data_o_173_sv2v_reg <= data_i[173];
      data_o_172_sv2v_reg <= data_i[172];
      data_o_171_sv2v_reg <= data_i[171];
      data_o_170_sv2v_reg <= data_i[170];
      data_o_169_sv2v_reg <= data_i[169];
      data_o_168_sv2v_reg <= data_i[168];
      data_o_167_sv2v_reg <= data_i[167];
      data_o_166_sv2v_reg <= data_i[166];
      data_o_165_sv2v_reg <= data_i[165];
      data_o_164_sv2v_reg <= data_i[164];
      data_o_163_sv2v_reg <= data_i[163];
      data_o_162_sv2v_reg <= data_i[162];
      data_o_161_sv2v_reg <= data_i[161];
      data_o_160_sv2v_reg <= data_i[160];
      data_o_159_sv2v_reg <= data_i[159];
      data_o_158_sv2v_reg <= data_i[158];
      data_o_157_sv2v_reg <= data_i[157];
      data_o_156_sv2v_reg <= data_i[156];
      data_o_155_sv2v_reg <= data_i[155];
      data_o_154_sv2v_reg <= data_i[154];
      data_o_153_sv2v_reg <= data_i[153];
      data_o_152_sv2v_reg <= data_i[152];
      data_o_151_sv2v_reg <= data_i[151];
      data_o_150_sv2v_reg <= data_i[150];
      data_o_149_sv2v_reg <= data_i[149];
      data_o_148_sv2v_reg <= data_i[148];
      data_o_147_sv2v_reg <= data_i[147];
      data_o_146_sv2v_reg <= data_i[146];
      data_o_145_sv2v_reg <= data_i[145];
      data_o_144_sv2v_reg <= data_i[144];
      data_o_143_sv2v_reg <= data_i[143];
      data_o_142_sv2v_reg <= data_i[142];
      data_o_141_sv2v_reg <= data_i[141];
      data_o_140_sv2v_reg <= data_i[140];
      data_o_139_sv2v_reg <= data_i[139];
      data_o_138_sv2v_reg <= data_i[138];
      data_o_137_sv2v_reg <= data_i[137];
      data_o_136_sv2v_reg <= data_i[136];
      data_o_135_sv2v_reg <= data_i[135];
      data_o_134_sv2v_reg <= data_i[134];
      data_o_133_sv2v_reg <= data_i[133];
      data_o_132_sv2v_reg <= data_i[132];
      data_o_131_sv2v_reg <= data_i[131];
      data_o_130_sv2v_reg <= data_i[130];
      data_o_129_sv2v_reg <= data_i[129];
      data_o_128_sv2v_reg <= data_i[128];
      data_o_127_sv2v_reg <= data_i[127];
      data_o_126_sv2v_reg <= data_i[126];
      data_o_125_sv2v_reg <= data_i[125];
      data_o_124_sv2v_reg <= data_i[124];
      data_o_123_sv2v_reg <= data_i[123];
      data_o_122_sv2v_reg <= data_i[122];
      data_o_121_sv2v_reg <= data_i[121];
      data_o_120_sv2v_reg <= data_i[120];
      data_o_119_sv2v_reg <= data_i[119];
      data_o_118_sv2v_reg <= data_i[118];
      data_o_117_sv2v_reg <= data_i[117];
      data_o_116_sv2v_reg <= data_i[116];
      data_o_115_sv2v_reg <= data_i[115];
      data_o_114_sv2v_reg <= data_i[114];
      data_o_113_sv2v_reg <= data_i[113];
      data_o_112_sv2v_reg <= data_i[112];
      data_o_111_sv2v_reg <= data_i[111];
      data_o_110_sv2v_reg <= data_i[110];
      data_o_109_sv2v_reg <= data_i[109];
      data_o_108_sv2v_reg <= data_i[108];
      data_o_107_sv2v_reg <= data_i[107];
      data_o_106_sv2v_reg <= data_i[106];
      data_o_105_sv2v_reg <= data_i[105];
      data_o_104_sv2v_reg <= data_i[104];
      data_o_103_sv2v_reg <= data_i[103];
      data_o_102_sv2v_reg <= data_i[102];
      data_o_101_sv2v_reg <= data_i[101];
      data_o_100_sv2v_reg <= data_i[100];
      data_o_99_sv2v_reg <= data_i[99];
      data_o_98_sv2v_reg <= data_i[98];
      data_o_97_sv2v_reg <= data_i[97];
      data_o_96_sv2v_reg <= data_i[96];
      data_o_95_sv2v_reg <= data_i[95];
      data_o_94_sv2v_reg <= data_i[94];
      data_o_93_sv2v_reg <= data_i[93];
      data_o_92_sv2v_reg <= data_i[92];
      data_o_91_sv2v_reg <= data_i[91];
      data_o_90_sv2v_reg <= data_i[90];
      data_o_89_sv2v_reg <= data_i[89];
      data_o_88_sv2v_reg <= data_i[88];
      data_o_87_sv2v_reg <= data_i[87];
      data_o_86_sv2v_reg <= data_i[86];
      data_o_85_sv2v_reg <= data_i[85];
      data_o_84_sv2v_reg <= data_i[84];
      data_o_83_sv2v_reg <= data_i[83];
      data_o_82_sv2v_reg <= data_i[82];
      data_o_81_sv2v_reg <= data_i[81];
      data_o_80_sv2v_reg <= data_i[80];
      data_o_79_sv2v_reg <= data_i[79];
      data_o_78_sv2v_reg <= data_i[78];
      data_o_77_sv2v_reg <= data_i[77];
      data_o_76_sv2v_reg <= data_i[76];
      data_o_75_sv2v_reg <= data_i[75];
      data_o_74_sv2v_reg <= data_i[74];
      data_o_73_sv2v_reg <= data_i[73];
      data_o_72_sv2v_reg <= data_i[72];
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module isSigNaNRecFN_expWidth11_sigWidth53
(
  in,
  isSigNaN
);

  input [64:0] in;
  output isSigNaN;
  wire isSigNaN,N0,N1,N2;
  assign N0 = in[62] & in[63];
  assign N1 = in[61] & N0;
  assign isSigNaN = N1 & N2;
  assign N2 = ~in[51];

endmodule



module bp_be_rec_to_raw_00
(
  rec_i,
  tag_i,
  raw_o
);

  input [64:0] rec_i;
  output [74:0] raw_o;
  input tag_i;
  wire [74:0] raw_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;
  wire [8:0] biased_sp;
  assign raw_o[0] = 1'b0;
  assign raw_o[1] = 1'b0;

  recFNToRawFN_expWidth11_sigWidth53
  rec2raw
  (
    .in(rec_i),
    .isNaN(raw_o[74]),
    .isInf(raw_o[73]),
    .isZero(raw_o[72]),
    .sign(raw_o[69]),
    .sExp(raw_o[68:56]),
    .sig(raw_o[55:2])
  );


  isSigNaNRecFN_expWidth11_sigWidth53
  is_snan
  (
    .in(rec_i),
    .isSigNaN(raw_o[71])
  );

  assign N3 = biased_sp < { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 };
  assign N5 = raw_o[67:56] < { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 };
  assign biased_sp = raw_o[64:56] + { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign raw_o[70] = (N0)? N4 : 
                     (N1)? N6 : 1'b0;
  assign N0 = tag_i;
  assign N1 = N2;
  assign N2 = ~tag_i;
  assign N4 = N11 & N3;
  assign N11 = N9 & N10;
  assign N9 = N7 & N8;
  assign N7 = ~raw_o[72];
  assign N8 = ~raw_o[73];
  assign N10 = ~raw_o[74];
  assign N6 = N13 & N5;
  assign N13 = N12 & N10;
  assign N12 = N7 & N8;

endmodule



module bsg_scan_width_p65_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [64:0] i;
  output [64:0] o;
  wire [64:0] o;
  wire t_6__64_,t_6__63_,t_6__62_,t_6__61_,t_6__60_,t_6__59_,t_6__58_,t_6__57_,
  t_6__56_,t_6__55_,t_6__54_,t_6__53_,t_6__52_,t_6__51_,t_6__50_,t_6__49_,t_6__48_,
  t_6__47_,t_6__46_,t_6__45_,t_6__44_,t_6__43_,t_6__42_,t_6__41_,t_6__40_,t_6__39_,
  t_6__38_,t_6__37_,t_6__36_,t_6__35_,t_6__34_,t_6__33_,t_6__32_,t_6__31_,t_6__30_,
  t_6__29_,t_6__28_,t_6__27_,t_6__26_,t_6__25_,t_6__24_,t_6__23_,t_6__22_,t_6__21_,
  t_6__20_,t_6__19_,t_6__18_,t_6__17_,t_6__16_,t_6__15_,t_6__14_,t_6__13_,t_6__12_,
  t_6__11_,t_6__10_,t_6__9_,t_6__8_,t_6__7_,t_6__6_,t_6__5_,t_6__4_,t_6__3_,t_6__2_,
  t_6__1_,t_6__0_,t_5__64_,t_5__63_,t_5__62_,t_5__61_,t_5__60_,t_5__59_,t_5__58_,
  t_5__57_,t_5__56_,t_5__55_,t_5__54_,t_5__53_,t_5__52_,t_5__51_,t_5__50_,t_5__49_,
  t_5__48_,t_5__47_,t_5__46_,t_5__45_,t_5__44_,t_5__43_,t_5__42_,t_5__41_,t_5__40_,
  t_5__39_,t_5__38_,t_5__37_,t_5__36_,t_5__35_,t_5__34_,t_5__33_,t_5__32_,
  t_5__31_,t_5__30_,t_5__29_,t_5__28_,t_5__27_,t_5__26_,t_5__25_,t_5__24_,t_5__23_,
  t_5__22_,t_5__21_,t_5__20_,t_5__19_,t_5__18_,t_5__17_,t_5__16_,t_5__15_,t_5__14_,
  t_5__13_,t_5__12_,t_5__11_,t_5__10_,t_5__9_,t_5__8_,t_5__7_,t_5__6_,t_5__5_,t_5__4_,
  t_5__3_,t_5__2_,t_5__1_,t_5__0_,t_4__64_,t_4__63_,t_4__62_,t_4__61_,t_4__60_,
  t_4__59_,t_4__58_,t_4__57_,t_4__56_,t_4__55_,t_4__54_,t_4__53_,t_4__52_,t_4__51_,
  t_4__50_,t_4__49_,t_4__48_,t_4__47_,t_4__46_,t_4__45_,t_4__44_,t_4__43_,t_4__42_,
  t_4__41_,t_4__40_,t_4__39_,t_4__38_,t_4__37_,t_4__36_,t_4__35_,t_4__34_,t_4__33_,
  t_4__32_,t_4__31_,t_4__30_,t_4__29_,t_4__28_,t_4__27_,t_4__26_,t_4__25_,t_4__24_,
  t_4__23_,t_4__22_,t_4__21_,t_4__20_,t_4__19_,t_4__18_,t_4__17_,t_4__16_,t_4__15_,
  t_4__14_,t_4__13_,t_4__12_,t_4__11_,t_4__10_,t_4__9_,t_4__8_,t_4__7_,t_4__6_,
  t_4__5_,t_4__4_,t_4__3_,t_4__2_,t_4__1_,t_4__0_,t_3__64_,t_3__63_,t_3__62_,
  t_3__61_,t_3__60_,t_3__59_,t_3__58_,t_3__57_,t_3__56_,t_3__55_,t_3__54_,t_3__53_,
  t_3__52_,t_3__51_,t_3__50_,t_3__49_,t_3__48_,t_3__47_,t_3__46_,t_3__45_,t_3__44_,
  t_3__43_,t_3__42_,t_3__41_,t_3__40_,t_3__39_,t_3__38_,t_3__37_,t_3__36_,t_3__35_,
  t_3__34_,t_3__33_,t_3__32_,t_3__31_,t_3__30_,t_3__29_,t_3__28_,t_3__27_,t_3__26_,
  t_3__25_,t_3__24_,t_3__23_,t_3__22_,t_3__21_,t_3__20_,t_3__19_,t_3__18_,t_3__17_,
  t_3__16_,t_3__15_,t_3__14_,t_3__13_,t_3__12_,t_3__11_,t_3__10_,t_3__9_,t_3__8_,
  t_3__7_,t_3__6_,t_3__5_,t_3__4_,t_3__3_,t_3__2_,t_3__1_,t_3__0_,t_2__64_,t_2__63_,
  t_2__62_,t_2__61_,t_2__60_,t_2__59_,t_2__58_,t_2__57_,t_2__56_,t_2__55_,t_2__54_,
  t_2__53_,t_2__52_,t_2__51_,t_2__50_,t_2__49_,t_2__48_,t_2__47_,t_2__46_,t_2__45_,
  t_2__44_,t_2__43_,t_2__42_,t_2__41_,t_2__40_,t_2__39_,t_2__38_,t_2__37_,
  t_2__36_,t_2__35_,t_2__34_,t_2__33_,t_2__32_,t_2__31_,t_2__30_,t_2__29_,t_2__28_,
  t_2__27_,t_2__26_,t_2__25_,t_2__24_,t_2__23_,t_2__22_,t_2__21_,t_2__20_,t_2__19_,
  t_2__18_,t_2__17_,t_2__16_,t_2__15_,t_2__14_,t_2__13_,t_2__12_,t_2__11_,t_2__10_,
  t_2__9_,t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,
  t_1__64_,t_1__63_,t_1__62_,t_1__61_,t_1__60_,t_1__59_,t_1__58_,t_1__57_,t_1__56_,
  t_1__55_,t_1__54_,t_1__53_,t_1__52_,t_1__51_,t_1__50_,t_1__49_,t_1__48_,t_1__47_,
  t_1__46_,t_1__45_,t_1__44_,t_1__43_,t_1__42_,t_1__41_,t_1__40_,t_1__39_,t_1__38_,
  t_1__37_,t_1__36_,t_1__35_,t_1__34_,t_1__33_,t_1__32_,t_1__31_,t_1__30_,t_1__29_,
  t_1__28_,t_1__27_,t_1__26_,t_1__25_,t_1__24_,t_1__23_,t_1__22_,t_1__21_,t_1__20_,
  t_1__19_,t_1__18_,t_1__17_,t_1__16_,t_1__15_,t_1__14_,t_1__13_,t_1__12_,
  t_1__11_,t_1__10_,t_1__9_,t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,
  t_1__1_,t_1__0_;
  assign t_1__64_ = i[0] | 1'b0;
  assign t_1__63_ = i[1] | i[0];
  assign t_1__62_ = i[2] | i[1];
  assign t_1__61_ = i[3] | i[2];
  assign t_1__60_ = i[4] | i[3];
  assign t_1__59_ = i[5] | i[4];
  assign t_1__58_ = i[6] | i[5];
  assign t_1__57_ = i[7] | i[6];
  assign t_1__56_ = i[8] | i[7];
  assign t_1__55_ = i[9] | i[8];
  assign t_1__54_ = i[10] | i[9];
  assign t_1__53_ = i[11] | i[10];
  assign t_1__52_ = i[12] | i[11];
  assign t_1__51_ = i[13] | i[12];
  assign t_1__50_ = i[14] | i[13];
  assign t_1__49_ = i[15] | i[14];
  assign t_1__48_ = i[16] | i[15];
  assign t_1__47_ = i[17] | i[16];
  assign t_1__46_ = i[18] | i[17];
  assign t_1__45_ = i[19] | i[18];
  assign t_1__44_ = i[20] | i[19];
  assign t_1__43_ = i[21] | i[20];
  assign t_1__42_ = i[22] | i[21];
  assign t_1__41_ = i[23] | i[22];
  assign t_1__40_ = i[24] | i[23];
  assign t_1__39_ = i[25] | i[24];
  assign t_1__38_ = i[26] | i[25];
  assign t_1__37_ = i[27] | i[26];
  assign t_1__36_ = i[28] | i[27];
  assign t_1__35_ = i[29] | i[28];
  assign t_1__34_ = i[30] | i[29];
  assign t_1__33_ = i[31] | i[30];
  assign t_1__32_ = i[32] | i[31];
  assign t_1__31_ = i[33] | i[32];
  assign t_1__30_ = i[34] | i[33];
  assign t_1__29_ = i[35] | i[34];
  assign t_1__28_ = i[36] | i[35];
  assign t_1__27_ = i[37] | i[36];
  assign t_1__26_ = i[38] | i[37];
  assign t_1__25_ = i[39] | i[38];
  assign t_1__24_ = i[40] | i[39];
  assign t_1__23_ = i[41] | i[40];
  assign t_1__22_ = i[42] | i[41];
  assign t_1__21_ = i[43] | i[42];
  assign t_1__20_ = i[44] | i[43];
  assign t_1__19_ = i[45] | i[44];
  assign t_1__18_ = i[46] | i[45];
  assign t_1__17_ = i[47] | i[46];
  assign t_1__16_ = i[48] | i[47];
  assign t_1__15_ = i[49] | i[48];
  assign t_1__14_ = i[50] | i[49];
  assign t_1__13_ = i[51] | i[50];
  assign t_1__12_ = i[52] | i[51];
  assign t_1__11_ = i[53] | i[52];
  assign t_1__10_ = i[54] | i[53];
  assign t_1__9_ = i[55] | i[54];
  assign t_1__8_ = i[56] | i[55];
  assign t_1__7_ = i[57] | i[56];
  assign t_1__6_ = i[58] | i[57];
  assign t_1__5_ = i[59] | i[58];
  assign t_1__4_ = i[60] | i[59];
  assign t_1__3_ = i[61] | i[60];
  assign t_1__2_ = i[62] | i[61];
  assign t_1__1_ = i[63] | i[62];
  assign t_1__0_ = i[64] | i[63];
  assign t_2__64_ = t_1__64_ | 1'b0;
  assign t_2__63_ = t_1__63_ | 1'b0;
  assign t_2__62_ = t_1__62_ | t_1__64_;
  assign t_2__61_ = t_1__61_ | t_1__63_;
  assign t_2__60_ = t_1__60_ | t_1__62_;
  assign t_2__59_ = t_1__59_ | t_1__61_;
  assign t_2__58_ = t_1__58_ | t_1__60_;
  assign t_2__57_ = t_1__57_ | t_1__59_;
  assign t_2__56_ = t_1__56_ | t_1__58_;
  assign t_2__55_ = t_1__55_ | t_1__57_;
  assign t_2__54_ = t_1__54_ | t_1__56_;
  assign t_2__53_ = t_1__53_ | t_1__55_;
  assign t_2__52_ = t_1__52_ | t_1__54_;
  assign t_2__51_ = t_1__51_ | t_1__53_;
  assign t_2__50_ = t_1__50_ | t_1__52_;
  assign t_2__49_ = t_1__49_ | t_1__51_;
  assign t_2__48_ = t_1__48_ | t_1__50_;
  assign t_2__47_ = t_1__47_ | t_1__49_;
  assign t_2__46_ = t_1__46_ | t_1__48_;
  assign t_2__45_ = t_1__45_ | t_1__47_;
  assign t_2__44_ = t_1__44_ | t_1__46_;
  assign t_2__43_ = t_1__43_ | t_1__45_;
  assign t_2__42_ = t_1__42_ | t_1__44_;
  assign t_2__41_ = t_1__41_ | t_1__43_;
  assign t_2__40_ = t_1__40_ | t_1__42_;
  assign t_2__39_ = t_1__39_ | t_1__41_;
  assign t_2__38_ = t_1__38_ | t_1__40_;
  assign t_2__37_ = t_1__37_ | t_1__39_;
  assign t_2__36_ = t_1__36_ | t_1__38_;
  assign t_2__35_ = t_1__35_ | t_1__37_;
  assign t_2__34_ = t_1__34_ | t_1__36_;
  assign t_2__33_ = t_1__33_ | t_1__35_;
  assign t_2__32_ = t_1__32_ | t_1__34_;
  assign t_2__31_ = t_1__31_ | t_1__33_;
  assign t_2__30_ = t_1__30_ | t_1__32_;
  assign t_2__29_ = t_1__29_ | t_1__31_;
  assign t_2__28_ = t_1__28_ | t_1__30_;
  assign t_2__27_ = t_1__27_ | t_1__29_;
  assign t_2__26_ = t_1__26_ | t_1__28_;
  assign t_2__25_ = t_1__25_ | t_1__27_;
  assign t_2__24_ = t_1__24_ | t_1__26_;
  assign t_2__23_ = t_1__23_ | t_1__25_;
  assign t_2__22_ = t_1__22_ | t_1__24_;
  assign t_2__21_ = t_1__21_ | t_1__23_;
  assign t_2__20_ = t_1__20_ | t_1__22_;
  assign t_2__19_ = t_1__19_ | t_1__21_;
  assign t_2__18_ = t_1__18_ | t_1__20_;
  assign t_2__17_ = t_1__17_ | t_1__19_;
  assign t_2__16_ = t_1__16_ | t_1__18_;
  assign t_2__15_ = t_1__15_ | t_1__17_;
  assign t_2__14_ = t_1__14_ | t_1__16_;
  assign t_2__13_ = t_1__13_ | t_1__15_;
  assign t_2__12_ = t_1__12_ | t_1__14_;
  assign t_2__11_ = t_1__11_ | t_1__13_;
  assign t_2__10_ = t_1__10_ | t_1__12_;
  assign t_2__9_ = t_1__9_ | t_1__11_;
  assign t_2__8_ = t_1__8_ | t_1__10_;
  assign t_2__7_ = t_1__7_ | t_1__9_;
  assign t_2__6_ = t_1__6_ | t_1__8_;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign t_3__64_ = t_2__64_ | 1'b0;
  assign t_3__63_ = t_2__63_ | 1'b0;
  assign t_3__62_ = t_2__62_ | 1'b0;
  assign t_3__61_ = t_2__61_ | 1'b0;
  assign t_3__60_ = t_2__60_ | t_2__64_;
  assign t_3__59_ = t_2__59_ | t_2__63_;
  assign t_3__58_ = t_2__58_ | t_2__62_;
  assign t_3__57_ = t_2__57_ | t_2__61_;
  assign t_3__56_ = t_2__56_ | t_2__60_;
  assign t_3__55_ = t_2__55_ | t_2__59_;
  assign t_3__54_ = t_2__54_ | t_2__58_;
  assign t_3__53_ = t_2__53_ | t_2__57_;
  assign t_3__52_ = t_2__52_ | t_2__56_;
  assign t_3__51_ = t_2__51_ | t_2__55_;
  assign t_3__50_ = t_2__50_ | t_2__54_;
  assign t_3__49_ = t_2__49_ | t_2__53_;
  assign t_3__48_ = t_2__48_ | t_2__52_;
  assign t_3__47_ = t_2__47_ | t_2__51_;
  assign t_3__46_ = t_2__46_ | t_2__50_;
  assign t_3__45_ = t_2__45_ | t_2__49_;
  assign t_3__44_ = t_2__44_ | t_2__48_;
  assign t_3__43_ = t_2__43_ | t_2__47_;
  assign t_3__42_ = t_2__42_ | t_2__46_;
  assign t_3__41_ = t_2__41_ | t_2__45_;
  assign t_3__40_ = t_2__40_ | t_2__44_;
  assign t_3__39_ = t_2__39_ | t_2__43_;
  assign t_3__38_ = t_2__38_ | t_2__42_;
  assign t_3__37_ = t_2__37_ | t_2__41_;
  assign t_3__36_ = t_2__36_ | t_2__40_;
  assign t_3__35_ = t_2__35_ | t_2__39_;
  assign t_3__34_ = t_2__34_ | t_2__38_;
  assign t_3__33_ = t_2__33_ | t_2__37_;
  assign t_3__32_ = t_2__32_ | t_2__36_;
  assign t_3__31_ = t_2__31_ | t_2__35_;
  assign t_3__30_ = t_2__30_ | t_2__34_;
  assign t_3__29_ = t_2__29_ | t_2__33_;
  assign t_3__28_ = t_2__28_ | t_2__32_;
  assign t_3__27_ = t_2__27_ | t_2__31_;
  assign t_3__26_ = t_2__26_ | t_2__30_;
  assign t_3__25_ = t_2__25_ | t_2__29_;
  assign t_3__24_ = t_2__24_ | t_2__28_;
  assign t_3__23_ = t_2__23_ | t_2__27_;
  assign t_3__22_ = t_2__22_ | t_2__26_;
  assign t_3__21_ = t_2__21_ | t_2__25_;
  assign t_3__20_ = t_2__20_ | t_2__24_;
  assign t_3__19_ = t_2__19_ | t_2__23_;
  assign t_3__18_ = t_2__18_ | t_2__22_;
  assign t_3__17_ = t_2__17_ | t_2__21_;
  assign t_3__16_ = t_2__16_ | t_2__20_;
  assign t_3__15_ = t_2__15_ | t_2__19_;
  assign t_3__14_ = t_2__14_ | t_2__18_;
  assign t_3__13_ = t_2__13_ | t_2__17_;
  assign t_3__12_ = t_2__12_ | t_2__16_;
  assign t_3__11_ = t_2__11_ | t_2__15_;
  assign t_3__10_ = t_2__10_ | t_2__14_;
  assign t_3__9_ = t_2__9_ | t_2__13_;
  assign t_3__8_ = t_2__8_ | t_2__12_;
  assign t_3__7_ = t_2__7_ | t_2__11_;
  assign t_3__6_ = t_2__6_ | t_2__10_;
  assign t_3__5_ = t_2__5_ | t_2__9_;
  assign t_3__4_ = t_2__4_ | t_2__8_;
  assign t_3__3_ = t_2__3_ | t_2__7_;
  assign t_3__2_ = t_2__2_ | t_2__6_;
  assign t_3__1_ = t_2__1_ | t_2__5_;
  assign t_3__0_ = t_2__0_ | t_2__4_;
  assign t_4__64_ = t_3__64_ | 1'b0;
  assign t_4__63_ = t_3__63_ | 1'b0;
  assign t_4__62_ = t_3__62_ | 1'b0;
  assign t_4__61_ = t_3__61_ | 1'b0;
  assign t_4__60_ = t_3__60_ | 1'b0;
  assign t_4__59_ = t_3__59_ | 1'b0;
  assign t_4__58_ = t_3__58_ | 1'b0;
  assign t_4__57_ = t_3__57_ | 1'b0;
  assign t_4__56_ = t_3__56_ | t_3__64_;
  assign t_4__55_ = t_3__55_ | t_3__63_;
  assign t_4__54_ = t_3__54_ | t_3__62_;
  assign t_4__53_ = t_3__53_ | t_3__61_;
  assign t_4__52_ = t_3__52_ | t_3__60_;
  assign t_4__51_ = t_3__51_ | t_3__59_;
  assign t_4__50_ = t_3__50_ | t_3__58_;
  assign t_4__49_ = t_3__49_ | t_3__57_;
  assign t_4__48_ = t_3__48_ | t_3__56_;
  assign t_4__47_ = t_3__47_ | t_3__55_;
  assign t_4__46_ = t_3__46_ | t_3__54_;
  assign t_4__45_ = t_3__45_ | t_3__53_;
  assign t_4__44_ = t_3__44_ | t_3__52_;
  assign t_4__43_ = t_3__43_ | t_3__51_;
  assign t_4__42_ = t_3__42_ | t_3__50_;
  assign t_4__41_ = t_3__41_ | t_3__49_;
  assign t_4__40_ = t_3__40_ | t_3__48_;
  assign t_4__39_ = t_3__39_ | t_3__47_;
  assign t_4__38_ = t_3__38_ | t_3__46_;
  assign t_4__37_ = t_3__37_ | t_3__45_;
  assign t_4__36_ = t_3__36_ | t_3__44_;
  assign t_4__35_ = t_3__35_ | t_3__43_;
  assign t_4__34_ = t_3__34_ | t_3__42_;
  assign t_4__33_ = t_3__33_ | t_3__41_;
  assign t_4__32_ = t_3__32_ | t_3__40_;
  assign t_4__31_ = t_3__31_ | t_3__39_;
  assign t_4__30_ = t_3__30_ | t_3__38_;
  assign t_4__29_ = t_3__29_ | t_3__37_;
  assign t_4__28_ = t_3__28_ | t_3__36_;
  assign t_4__27_ = t_3__27_ | t_3__35_;
  assign t_4__26_ = t_3__26_ | t_3__34_;
  assign t_4__25_ = t_3__25_ | t_3__33_;
  assign t_4__24_ = t_3__24_ | t_3__32_;
  assign t_4__23_ = t_3__23_ | t_3__31_;
  assign t_4__22_ = t_3__22_ | t_3__30_;
  assign t_4__21_ = t_3__21_ | t_3__29_;
  assign t_4__20_ = t_3__20_ | t_3__28_;
  assign t_4__19_ = t_3__19_ | t_3__27_;
  assign t_4__18_ = t_3__18_ | t_3__26_;
  assign t_4__17_ = t_3__17_ | t_3__25_;
  assign t_4__16_ = t_3__16_ | t_3__24_;
  assign t_4__15_ = t_3__15_ | t_3__23_;
  assign t_4__14_ = t_3__14_ | t_3__22_;
  assign t_4__13_ = t_3__13_ | t_3__21_;
  assign t_4__12_ = t_3__12_ | t_3__20_;
  assign t_4__11_ = t_3__11_ | t_3__19_;
  assign t_4__10_ = t_3__10_ | t_3__18_;
  assign t_4__9_ = t_3__9_ | t_3__17_;
  assign t_4__8_ = t_3__8_ | t_3__16_;
  assign t_4__7_ = t_3__7_ | t_3__15_;
  assign t_4__6_ = t_3__6_ | t_3__14_;
  assign t_4__5_ = t_3__5_ | t_3__13_;
  assign t_4__4_ = t_3__4_ | t_3__12_;
  assign t_4__3_ = t_3__3_ | t_3__11_;
  assign t_4__2_ = t_3__2_ | t_3__10_;
  assign t_4__1_ = t_3__1_ | t_3__9_;
  assign t_4__0_ = t_3__0_ | t_3__8_;
  assign t_5__64_ = t_4__64_ | 1'b0;
  assign t_5__63_ = t_4__63_ | 1'b0;
  assign t_5__62_ = t_4__62_ | 1'b0;
  assign t_5__61_ = t_4__61_ | 1'b0;
  assign t_5__60_ = t_4__60_ | 1'b0;
  assign t_5__59_ = t_4__59_ | 1'b0;
  assign t_5__58_ = t_4__58_ | 1'b0;
  assign t_5__57_ = t_4__57_ | 1'b0;
  assign t_5__56_ = t_4__56_ | 1'b0;
  assign t_5__55_ = t_4__55_ | 1'b0;
  assign t_5__54_ = t_4__54_ | 1'b0;
  assign t_5__53_ = t_4__53_ | 1'b0;
  assign t_5__52_ = t_4__52_ | 1'b0;
  assign t_5__51_ = t_4__51_ | 1'b0;
  assign t_5__50_ = t_4__50_ | 1'b0;
  assign t_5__49_ = t_4__49_ | 1'b0;
  assign t_5__48_ = t_4__48_ | t_4__64_;
  assign t_5__47_ = t_4__47_ | t_4__63_;
  assign t_5__46_ = t_4__46_ | t_4__62_;
  assign t_5__45_ = t_4__45_ | t_4__61_;
  assign t_5__44_ = t_4__44_ | t_4__60_;
  assign t_5__43_ = t_4__43_ | t_4__59_;
  assign t_5__42_ = t_4__42_ | t_4__58_;
  assign t_5__41_ = t_4__41_ | t_4__57_;
  assign t_5__40_ = t_4__40_ | t_4__56_;
  assign t_5__39_ = t_4__39_ | t_4__55_;
  assign t_5__38_ = t_4__38_ | t_4__54_;
  assign t_5__37_ = t_4__37_ | t_4__53_;
  assign t_5__36_ = t_4__36_ | t_4__52_;
  assign t_5__35_ = t_4__35_ | t_4__51_;
  assign t_5__34_ = t_4__34_ | t_4__50_;
  assign t_5__33_ = t_4__33_ | t_4__49_;
  assign t_5__32_ = t_4__32_ | t_4__48_;
  assign t_5__31_ = t_4__31_ | t_4__47_;
  assign t_5__30_ = t_4__30_ | t_4__46_;
  assign t_5__29_ = t_4__29_ | t_4__45_;
  assign t_5__28_ = t_4__28_ | t_4__44_;
  assign t_5__27_ = t_4__27_ | t_4__43_;
  assign t_5__26_ = t_4__26_ | t_4__42_;
  assign t_5__25_ = t_4__25_ | t_4__41_;
  assign t_5__24_ = t_4__24_ | t_4__40_;
  assign t_5__23_ = t_4__23_ | t_4__39_;
  assign t_5__22_ = t_4__22_ | t_4__38_;
  assign t_5__21_ = t_4__21_ | t_4__37_;
  assign t_5__20_ = t_4__20_ | t_4__36_;
  assign t_5__19_ = t_4__19_ | t_4__35_;
  assign t_5__18_ = t_4__18_ | t_4__34_;
  assign t_5__17_ = t_4__17_ | t_4__33_;
  assign t_5__16_ = t_4__16_ | t_4__32_;
  assign t_5__15_ = t_4__15_ | t_4__31_;
  assign t_5__14_ = t_4__14_ | t_4__30_;
  assign t_5__13_ = t_4__13_ | t_4__29_;
  assign t_5__12_ = t_4__12_ | t_4__28_;
  assign t_5__11_ = t_4__11_ | t_4__27_;
  assign t_5__10_ = t_4__10_ | t_4__26_;
  assign t_5__9_ = t_4__9_ | t_4__25_;
  assign t_5__8_ = t_4__8_ | t_4__24_;
  assign t_5__7_ = t_4__7_ | t_4__23_;
  assign t_5__6_ = t_4__6_ | t_4__22_;
  assign t_5__5_ = t_4__5_ | t_4__21_;
  assign t_5__4_ = t_4__4_ | t_4__20_;
  assign t_5__3_ = t_4__3_ | t_4__19_;
  assign t_5__2_ = t_4__2_ | t_4__18_;
  assign t_5__1_ = t_4__1_ | t_4__17_;
  assign t_5__0_ = t_4__0_ | t_4__16_;
  assign t_6__64_ = t_5__64_ | 1'b0;
  assign t_6__63_ = t_5__63_ | 1'b0;
  assign t_6__62_ = t_5__62_ | 1'b0;
  assign t_6__61_ = t_5__61_ | 1'b0;
  assign t_6__60_ = t_5__60_ | 1'b0;
  assign t_6__59_ = t_5__59_ | 1'b0;
  assign t_6__58_ = t_5__58_ | 1'b0;
  assign t_6__57_ = t_5__57_ | 1'b0;
  assign t_6__56_ = t_5__56_ | 1'b0;
  assign t_6__55_ = t_5__55_ | 1'b0;
  assign t_6__54_ = t_5__54_ | 1'b0;
  assign t_6__53_ = t_5__53_ | 1'b0;
  assign t_6__52_ = t_5__52_ | 1'b0;
  assign t_6__51_ = t_5__51_ | 1'b0;
  assign t_6__50_ = t_5__50_ | 1'b0;
  assign t_6__49_ = t_5__49_ | 1'b0;
  assign t_6__48_ = t_5__48_ | 1'b0;
  assign t_6__47_ = t_5__47_ | 1'b0;
  assign t_6__46_ = t_5__46_ | 1'b0;
  assign t_6__45_ = t_5__45_ | 1'b0;
  assign t_6__44_ = t_5__44_ | 1'b0;
  assign t_6__43_ = t_5__43_ | 1'b0;
  assign t_6__42_ = t_5__42_ | 1'b0;
  assign t_6__41_ = t_5__41_ | 1'b0;
  assign t_6__40_ = t_5__40_ | 1'b0;
  assign t_6__39_ = t_5__39_ | 1'b0;
  assign t_6__38_ = t_5__38_ | 1'b0;
  assign t_6__37_ = t_5__37_ | 1'b0;
  assign t_6__36_ = t_5__36_ | 1'b0;
  assign t_6__35_ = t_5__35_ | 1'b0;
  assign t_6__34_ = t_5__34_ | 1'b0;
  assign t_6__33_ = t_5__33_ | 1'b0;
  assign t_6__32_ = t_5__32_ | t_5__64_;
  assign t_6__31_ = t_5__31_ | t_5__63_;
  assign t_6__30_ = t_5__30_ | t_5__62_;
  assign t_6__29_ = t_5__29_ | t_5__61_;
  assign t_6__28_ = t_5__28_ | t_5__60_;
  assign t_6__27_ = t_5__27_ | t_5__59_;
  assign t_6__26_ = t_5__26_ | t_5__58_;
  assign t_6__25_ = t_5__25_ | t_5__57_;
  assign t_6__24_ = t_5__24_ | t_5__56_;
  assign t_6__23_ = t_5__23_ | t_5__55_;
  assign t_6__22_ = t_5__22_ | t_5__54_;
  assign t_6__21_ = t_5__21_ | t_5__53_;
  assign t_6__20_ = t_5__20_ | t_5__52_;
  assign t_6__19_ = t_5__19_ | t_5__51_;
  assign t_6__18_ = t_5__18_ | t_5__50_;
  assign t_6__17_ = t_5__17_ | t_5__49_;
  assign t_6__16_ = t_5__16_ | t_5__48_;
  assign t_6__15_ = t_5__15_ | t_5__47_;
  assign t_6__14_ = t_5__14_ | t_5__46_;
  assign t_6__13_ = t_5__13_ | t_5__45_;
  assign t_6__12_ = t_5__12_ | t_5__44_;
  assign t_6__11_ = t_5__11_ | t_5__43_;
  assign t_6__10_ = t_5__10_ | t_5__42_;
  assign t_6__9_ = t_5__9_ | t_5__41_;
  assign t_6__8_ = t_5__8_ | t_5__40_;
  assign t_6__7_ = t_5__7_ | t_5__39_;
  assign t_6__6_ = t_5__6_ | t_5__38_;
  assign t_6__5_ = t_5__5_ | t_5__37_;
  assign t_6__4_ = t_5__4_ | t_5__36_;
  assign t_6__3_ = t_5__3_ | t_5__35_;
  assign t_6__2_ = t_5__2_ | t_5__34_;
  assign t_6__1_ = t_5__1_ | t_5__33_;
  assign t_6__0_ = t_5__0_ | t_5__32_;
  assign o[0] = t_6__64_ | 1'b0;
  assign o[1] = t_6__63_ | 1'b0;
  assign o[2] = t_6__62_ | 1'b0;
  assign o[3] = t_6__61_ | 1'b0;
  assign o[4] = t_6__60_ | 1'b0;
  assign o[5] = t_6__59_ | 1'b0;
  assign o[6] = t_6__58_ | 1'b0;
  assign o[7] = t_6__57_ | 1'b0;
  assign o[8] = t_6__56_ | 1'b0;
  assign o[9] = t_6__55_ | 1'b0;
  assign o[10] = t_6__54_ | 1'b0;
  assign o[11] = t_6__53_ | 1'b0;
  assign o[12] = t_6__52_ | 1'b0;
  assign o[13] = t_6__51_ | 1'b0;
  assign o[14] = t_6__50_ | 1'b0;
  assign o[15] = t_6__49_ | 1'b0;
  assign o[16] = t_6__48_ | 1'b0;
  assign o[17] = t_6__47_ | 1'b0;
  assign o[18] = t_6__46_ | 1'b0;
  assign o[19] = t_6__45_ | 1'b0;
  assign o[20] = t_6__44_ | 1'b0;
  assign o[21] = t_6__43_ | 1'b0;
  assign o[22] = t_6__42_ | 1'b0;
  assign o[23] = t_6__41_ | 1'b0;
  assign o[24] = t_6__40_ | 1'b0;
  assign o[25] = t_6__39_ | 1'b0;
  assign o[26] = t_6__38_ | 1'b0;
  assign o[27] = t_6__37_ | 1'b0;
  assign o[28] = t_6__36_ | 1'b0;
  assign o[29] = t_6__35_ | 1'b0;
  assign o[30] = t_6__34_ | 1'b0;
  assign o[31] = t_6__33_ | 1'b0;
  assign o[32] = t_6__32_ | 1'b0;
  assign o[33] = t_6__31_ | 1'b0;
  assign o[34] = t_6__30_ | 1'b0;
  assign o[35] = t_6__29_ | 1'b0;
  assign o[36] = t_6__28_ | 1'b0;
  assign o[37] = t_6__27_ | 1'b0;
  assign o[38] = t_6__26_ | 1'b0;
  assign o[39] = t_6__25_ | 1'b0;
  assign o[40] = t_6__24_ | 1'b0;
  assign o[41] = t_6__23_ | 1'b0;
  assign o[42] = t_6__22_ | 1'b0;
  assign o[43] = t_6__21_ | 1'b0;
  assign o[44] = t_6__20_ | 1'b0;
  assign o[45] = t_6__19_ | 1'b0;
  assign o[46] = t_6__18_ | 1'b0;
  assign o[47] = t_6__17_ | 1'b0;
  assign o[48] = t_6__16_ | 1'b0;
  assign o[49] = t_6__15_ | 1'b0;
  assign o[50] = t_6__14_ | 1'b0;
  assign o[51] = t_6__13_ | 1'b0;
  assign o[52] = t_6__12_ | 1'b0;
  assign o[53] = t_6__11_ | 1'b0;
  assign o[54] = t_6__10_ | 1'b0;
  assign o[55] = t_6__9_ | 1'b0;
  assign o[56] = t_6__8_ | 1'b0;
  assign o[57] = t_6__7_ | 1'b0;
  assign o[58] = t_6__6_ | 1'b0;
  assign o[59] = t_6__5_ | 1'b0;
  assign o[60] = t_6__4_ | 1'b0;
  assign o[61] = t_6__3_ | 1'b0;
  assign o[62] = t_6__2_ | 1'b0;
  assign o[63] = t_6__1_ | 1'b0;
  assign o[64] = t_6__0_ | t_6__64_;

endmodule



module bsg_priority_encode_one_hot_out_width_p65_lo_to_hi_p1
(
  i,
  o,
  v_o
);

  input [64:0] i;
  output [64:0] o;
  output v_o;
  wire [64:0] o;
  wire v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63;
  wire [63:1] scan_lo;

  bsg_scan_width_p65_or_p1_lo_to_hi_p1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, scan_lo, o[0:0] })
  );

  assign o[64] = v_o & N0;
  assign N0 = ~scan_lo[63];
  assign o[63] = scan_lo[63] & N1;
  assign N1 = ~scan_lo[62];
  assign o[62] = scan_lo[62] & N2;
  assign N2 = ~scan_lo[61];
  assign o[61] = scan_lo[61] & N3;
  assign N3 = ~scan_lo[60];
  assign o[60] = scan_lo[60] & N4;
  assign N4 = ~scan_lo[59];
  assign o[59] = scan_lo[59] & N5;
  assign N5 = ~scan_lo[58];
  assign o[58] = scan_lo[58] & N6;
  assign N6 = ~scan_lo[57];
  assign o[57] = scan_lo[57] & N7;
  assign N7 = ~scan_lo[56];
  assign o[56] = scan_lo[56] & N8;
  assign N8 = ~scan_lo[55];
  assign o[55] = scan_lo[55] & N9;
  assign N9 = ~scan_lo[54];
  assign o[54] = scan_lo[54] & N10;
  assign N10 = ~scan_lo[53];
  assign o[53] = scan_lo[53] & N11;
  assign N11 = ~scan_lo[52];
  assign o[52] = scan_lo[52] & N12;
  assign N12 = ~scan_lo[51];
  assign o[51] = scan_lo[51] & N13;
  assign N13 = ~scan_lo[50];
  assign o[50] = scan_lo[50] & N14;
  assign N14 = ~scan_lo[49];
  assign o[49] = scan_lo[49] & N15;
  assign N15 = ~scan_lo[48];
  assign o[48] = scan_lo[48] & N16;
  assign N16 = ~scan_lo[47];
  assign o[47] = scan_lo[47] & N17;
  assign N17 = ~scan_lo[46];
  assign o[46] = scan_lo[46] & N18;
  assign N18 = ~scan_lo[45];
  assign o[45] = scan_lo[45] & N19;
  assign N19 = ~scan_lo[44];
  assign o[44] = scan_lo[44] & N20;
  assign N20 = ~scan_lo[43];
  assign o[43] = scan_lo[43] & N21;
  assign N21 = ~scan_lo[42];
  assign o[42] = scan_lo[42] & N22;
  assign N22 = ~scan_lo[41];
  assign o[41] = scan_lo[41] & N23;
  assign N23 = ~scan_lo[40];
  assign o[40] = scan_lo[40] & N24;
  assign N24 = ~scan_lo[39];
  assign o[39] = scan_lo[39] & N25;
  assign N25 = ~scan_lo[38];
  assign o[38] = scan_lo[38] & N26;
  assign N26 = ~scan_lo[37];
  assign o[37] = scan_lo[37] & N27;
  assign N27 = ~scan_lo[36];
  assign o[36] = scan_lo[36] & N28;
  assign N28 = ~scan_lo[35];
  assign o[35] = scan_lo[35] & N29;
  assign N29 = ~scan_lo[34];
  assign o[34] = scan_lo[34] & N30;
  assign N30 = ~scan_lo[33];
  assign o[33] = scan_lo[33] & N31;
  assign N31 = ~scan_lo[32];
  assign o[32] = scan_lo[32] & N32;
  assign N32 = ~scan_lo[31];
  assign o[31] = scan_lo[31] & N33;
  assign N33 = ~scan_lo[30];
  assign o[30] = scan_lo[30] & N34;
  assign N34 = ~scan_lo[29];
  assign o[29] = scan_lo[29] & N35;
  assign N35 = ~scan_lo[28];
  assign o[28] = scan_lo[28] & N36;
  assign N36 = ~scan_lo[27];
  assign o[27] = scan_lo[27] & N37;
  assign N37 = ~scan_lo[26];
  assign o[26] = scan_lo[26] & N38;
  assign N38 = ~scan_lo[25];
  assign o[25] = scan_lo[25] & N39;
  assign N39 = ~scan_lo[24];
  assign o[24] = scan_lo[24] & N40;
  assign N40 = ~scan_lo[23];
  assign o[23] = scan_lo[23] & N41;
  assign N41 = ~scan_lo[22];
  assign o[22] = scan_lo[22] & N42;
  assign N42 = ~scan_lo[21];
  assign o[21] = scan_lo[21] & N43;
  assign N43 = ~scan_lo[20];
  assign o[20] = scan_lo[20] & N44;
  assign N44 = ~scan_lo[19];
  assign o[19] = scan_lo[19] & N45;
  assign N45 = ~scan_lo[18];
  assign o[18] = scan_lo[18] & N46;
  assign N46 = ~scan_lo[17];
  assign o[17] = scan_lo[17] & N47;
  assign N47 = ~scan_lo[16];
  assign o[16] = scan_lo[16] & N48;
  assign N48 = ~scan_lo[15];
  assign o[15] = scan_lo[15] & N49;
  assign N49 = ~scan_lo[14];
  assign o[14] = scan_lo[14] & N50;
  assign N50 = ~scan_lo[13];
  assign o[13] = scan_lo[13] & N51;
  assign N51 = ~scan_lo[12];
  assign o[12] = scan_lo[12] & N52;
  assign N52 = ~scan_lo[11];
  assign o[11] = scan_lo[11] & N53;
  assign N53 = ~scan_lo[10];
  assign o[10] = scan_lo[10] & N54;
  assign N54 = ~scan_lo[9];
  assign o[9] = scan_lo[9] & N55;
  assign N55 = ~scan_lo[8];
  assign o[8] = scan_lo[8] & N56;
  assign N56 = ~scan_lo[7];
  assign o[7] = scan_lo[7] & N57;
  assign N57 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N58;
  assign N58 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N59;
  assign N59 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N60;
  assign N60 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N61;
  assign N61 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N62;
  assign N62 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N63;
  assign N63 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p65_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [64:0] i;
  output [6:0] addr_o;
  output v_o;
  wire [6:0] addr_o;
  wire v_o,v_3__120_,v_3__112_,v_3__104_,v_3__96_,v_3__88_,v_3__80_,v_3__72_,v_3__64_,
  v_3__56_,v_3__48_,v_3__40_,v_3__32_,v_3__24_,v_3__16_,v_3__8_,v_3__0_,v_2__124_,
  v_2__120_,v_2__116_,v_2__112_,v_2__108_,v_2__104_,v_2__100_,v_2__96_,v_2__92_,
  v_2__88_,v_2__84_,v_2__80_,v_2__76_,v_2__72_,v_2__68_,v_2__64_,v_2__60_,v_2__56_,
  v_2__52_,v_2__48_,v_2__44_,v_2__40_,v_2__36_,v_2__32_,v_2__28_,v_2__24_,v_2__20_,
  v_2__16_,v_2__12_,v_2__8_,v_2__4_,v_2__0_,v_1__126_,v_1__124_,v_1__122_,
  v_1__120_,v_1__118_,v_1__116_,v_1__114_,v_1__112_,v_1__110_,v_1__108_,v_1__106_,
  v_1__104_,v_1__102_,v_1__100_,v_1__98_,v_1__96_,v_1__94_,v_1__92_,v_1__90_,v_1__88_,
  v_1__86_,v_1__84_,v_1__82_,v_1__80_,v_1__78_,v_1__76_,v_1__74_,v_1__72_,v_1__70_,
  v_1__68_,v_1__66_,v_1__64_,v_1__62_,v_1__60_,v_1__58_,v_1__56_,v_1__54_,v_1__52_,
  v_1__50_,v_1__48_,v_1__46_,v_1__44_,v_1__42_,v_1__40_,v_1__38_,v_1__36_,v_1__34_,
  v_1__32_,v_1__30_,v_1__28_,v_1__26_,v_1__24_,v_1__22_,v_1__20_,v_1__18_,v_1__16_,
  v_1__14_,v_1__12_,v_1__10_,v_1__8_,v_1__6_,v_1__4_,v_1__2_,v_1__0_,addr_3__121_,
  addr_3__120_,addr_3__113_,addr_3__112_,addr_3__105_,addr_3__104_,addr_3__97_,
  addr_3__96_,addr_3__89_,addr_3__88_,addr_3__81_,addr_3__80_,addr_3__73_,addr_3__72_,
  addr_3__65_,addr_3__64_,addr_3__57_,addr_3__56_,addr_3__49_,addr_3__48_,
  addr_3__41_,addr_3__40_,addr_3__33_,addr_3__32_,addr_3__25_,addr_3__24_,addr_3__17_,
  addr_3__16_,addr_3__9_,addr_3__8_,addr_3__1_,addr_3__0_,addr_2__124_,addr_2__120_,
  addr_2__116_,addr_2__112_,addr_2__108_,addr_2__104_,addr_2__100_,addr_2__96_,
  addr_2__92_,addr_2__88_,addr_2__84_,addr_2__80_,addr_2__76_,addr_2__72_,addr_2__68_,
  addr_2__64_,addr_2__60_,addr_2__56_,addr_2__52_,addr_2__48_,addr_2__44_,
  addr_2__40_,addr_2__36_,addr_2__32_,addr_2__28_,addr_2__24_,addr_2__20_,addr_2__16_,
  addr_2__12_,addr_2__8_,addr_2__4_,addr_2__0_,v_6__0_,v_5__96_,v_5__64_,v_5__32_,
  v_5__0_,v_4__112_,v_4__96_,v_4__80_,v_4__64_,v_4__48_,v_4__32_,v_4__16_,v_4__0_,
  addr_6__68_,addr_6__67_,addr_6__66_,addr_6__65_,addr_6__64_,addr_6__4_,addr_6__3_,
  addr_6__2_,addr_6__1_,addr_6__0_,addr_5__99_,addr_5__98_,addr_5__97_,addr_5__96_,
  addr_5__67_,addr_5__66_,addr_5__65_,addr_5__64_,addr_5__35_,addr_5__34_,
  addr_5__33_,addr_5__32_,addr_5__3_,addr_5__2_,addr_5__1_,addr_5__0_,addr_4__114_,
  addr_4__113_,addr_4__112_,addr_4__98_,addr_4__97_,addr_4__96_,addr_4__82_,addr_4__81_,
  addr_4__80_,addr_4__66_,addr_4__65_,addr_4__64_,addr_4__50_,addr_4__49_,
  addr_4__48_,addr_4__34_,addr_4__33_,addr_4__32_,addr_4__18_,addr_4__17_,addr_4__16_,
  addr_4__2_,addr_4__1_,addr_4__0_;
  assign v_1__0_ = i[1] | i[0];
  assign v_1__2_ = i[3] | i[2];
  assign v_1__4_ = i[5] | i[4];
  assign v_1__6_ = i[7] | i[6];
  assign v_1__8_ = i[9] | i[8];
  assign v_1__10_ = i[11] | i[10];
  assign v_1__12_ = i[13] | i[12];
  assign v_1__14_ = i[15] | i[14];
  assign v_1__16_ = i[17] | i[16];
  assign v_1__18_ = i[19] | i[18];
  assign v_1__20_ = i[21] | i[20];
  assign v_1__22_ = i[23] | i[22];
  assign v_1__24_ = i[25] | i[24];
  assign v_1__26_ = i[27] | i[26];
  assign v_1__28_ = i[29] | i[28];
  assign v_1__30_ = i[31] | i[30];
  assign v_1__32_ = i[33] | i[32];
  assign v_1__34_ = i[35] | i[34];
  assign v_1__36_ = i[37] | i[36];
  assign v_1__38_ = i[39] | i[38];
  assign v_1__40_ = i[41] | i[40];
  assign v_1__42_ = i[43] | i[42];
  assign v_1__44_ = i[45] | i[44];
  assign v_1__46_ = i[47] | i[46];
  assign v_1__48_ = i[49] | i[48];
  assign v_1__50_ = i[51] | i[50];
  assign v_1__52_ = i[53] | i[52];
  assign v_1__54_ = i[55] | i[54];
  assign v_1__56_ = i[57] | i[56];
  assign v_1__58_ = i[59] | i[58];
  assign v_1__60_ = i[61] | i[60];
  assign v_1__62_ = i[63] | i[62];
  assign v_1__64_ = 1'b0 | i[64];
  assign v_1__66_ = 1'b0 | 1'b0;
  assign v_1__68_ = 1'b0 | 1'b0;
  assign v_1__70_ = 1'b0 | 1'b0;
  assign v_1__72_ = 1'b0 | 1'b0;
  assign v_1__74_ = 1'b0 | 1'b0;
  assign v_1__76_ = 1'b0 | 1'b0;
  assign v_1__78_ = 1'b0 | 1'b0;
  assign v_1__80_ = 1'b0 | 1'b0;
  assign v_1__82_ = 1'b0 | 1'b0;
  assign v_1__84_ = 1'b0 | 1'b0;
  assign v_1__86_ = 1'b0 | 1'b0;
  assign v_1__88_ = 1'b0 | 1'b0;
  assign v_1__90_ = 1'b0 | 1'b0;
  assign v_1__92_ = 1'b0 | 1'b0;
  assign v_1__94_ = 1'b0 | 1'b0;
  assign v_1__96_ = 1'b0 | 1'b0;
  assign v_1__98_ = 1'b0 | 1'b0;
  assign v_1__100_ = 1'b0 | 1'b0;
  assign v_1__102_ = 1'b0 | 1'b0;
  assign v_1__104_ = 1'b0 | 1'b0;
  assign v_1__106_ = 1'b0 | 1'b0;
  assign v_1__108_ = 1'b0 | 1'b0;
  assign v_1__110_ = 1'b0 | 1'b0;
  assign v_1__112_ = 1'b0 | 1'b0;
  assign v_1__114_ = 1'b0 | 1'b0;
  assign v_1__116_ = 1'b0 | 1'b0;
  assign v_1__118_ = 1'b0 | 1'b0;
  assign v_1__120_ = 1'b0 | 1'b0;
  assign v_1__122_ = 1'b0 | 1'b0;
  assign v_1__124_ = 1'b0 | 1'b0;
  assign v_1__126_ = 1'b0 | 1'b0;
  assign v_2__0_ = v_1__2_ | v_1__0_;
  assign addr_2__0_ = i[1] | i[3];
  assign v_2__4_ = v_1__6_ | v_1__4_;
  assign addr_2__4_ = i[5] | i[7];
  assign v_2__8_ = v_1__10_ | v_1__8_;
  assign addr_2__8_ = i[9] | i[11];
  assign v_2__12_ = v_1__14_ | v_1__12_;
  assign addr_2__12_ = i[13] | i[15];
  assign v_2__16_ = v_1__18_ | v_1__16_;
  assign addr_2__16_ = i[17] | i[19];
  assign v_2__20_ = v_1__22_ | v_1__20_;
  assign addr_2__20_ = i[21] | i[23];
  assign v_2__24_ = v_1__26_ | v_1__24_;
  assign addr_2__24_ = i[25] | i[27];
  assign v_2__28_ = v_1__30_ | v_1__28_;
  assign addr_2__28_ = i[29] | i[31];
  assign v_2__32_ = v_1__34_ | v_1__32_;
  assign addr_2__32_ = i[33] | i[35];
  assign v_2__36_ = v_1__38_ | v_1__36_;
  assign addr_2__36_ = i[37] | i[39];
  assign v_2__40_ = v_1__42_ | v_1__40_;
  assign addr_2__40_ = i[41] | i[43];
  assign v_2__44_ = v_1__46_ | v_1__44_;
  assign addr_2__44_ = i[45] | i[47];
  assign v_2__48_ = v_1__50_ | v_1__48_;
  assign addr_2__48_ = i[49] | i[51];
  assign v_2__52_ = v_1__54_ | v_1__52_;
  assign addr_2__52_ = i[53] | i[55];
  assign v_2__56_ = v_1__58_ | v_1__56_;
  assign addr_2__56_ = i[57] | i[59];
  assign v_2__60_ = v_1__62_ | v_1__60_;
  assign addr_2__60_ = i[61] | i[63];
  assign v_2__64_ = v_1__66_ | v_1__64_;
  assign addr_2__64_ = 1'b0 | 1'b0;
  assign v_2__68_ = v_1__70_ | v_1__68_;
  assign addr_2__68_ = 1'b0 | 1'b0;
  assign v_2__72_ = v_1__74_ | v_1__72_;
  assign addr_2__72_ = 1'b0 | 1'b0;
  assign v_2__76_ = v_1__78_ | v_1__76_;
  assign addr_2__76_ = 1'b0 | 1'b0;
  assign v_2__80_ = v_1__82_ | v_1__80_;
  assign addr_2__80_ = 1'b0 | 1'b0;
  assign v_2__84_ = v_1__86_ | v_1__84_;
  assign addr_2__84_ = 1'b0 | 1'b0;
  assign v_2__88_ = v_1__90_ | v_1__88_;
  assign addr_2__88_ = 1'b0 | 1'b0;
  assign v_2__92_ = v_1__94_ | v_1__92_;
  assign addr_2__92_ = 1'b0 | 1'b0;
  assign v_2__96_ = v_1__98_ | v_1__96_;
  assign addr_2__96_ = 1'b0 | 1'b0;
  assign v_2__100_ = v_1__102_ | v_1__100_;
  assign addr_2__100_ = 1'b0 | 1'b0;
  assign v_2__104_ = v_1__106_ | v_1__104_;
  assign addr_2__104_ = 1'b0 | 1'b0;
  assign v_2__108_ = v_1__110_ | v_1__108_;
  assign addr_2__108_ = 1'b0 | 1'b0;
  assign v_2__112_ = v_1__114_ | v_1__112_;
  assign addr_2__112_ = 1'b0 | 1'b0;
  assign v_2__116_ = v_1__118_ | v_1__116_;
  assign addr_2__116_ = 1'b0 | 1'b0;
  assign v_2__120_ = v_1__122_ | v_1__120_;
  assign addr_2__120_ = 1'b0 | 1'b0;
  assign v_2__124_ = v_1__126_ | v_1__124_;
  assign addr_2__124_ = 1'b0 | 1'b0;
  assign v_3__0_ = v_2__4_ | v_2__0_;
  assign addr_3__1_ = v_1__2_ | v_1__6_;
  assign addr_3__0_ = addr_2__0_ | addr_2__4_;
  assign v_3__8_ = v_2__12_ | v_2__8_;
  assign addr_3__9_ = v_1__10_ | v_1__14_;
  assign addr_3__8_ = addr_2__8_ | addr_2__12_;
  assign v_3__16_ = v_2__20_ | v_2__16_;
  assign addr_3__17_ = v_1__18_ | v_1__22_;
  assign addr_3__16_ = addr_2__16_ | addr_2__20_;
  assign v_3__24_ = v_2__28_ | v_2__24_;
  assign addr_3__25_ = v_1__26_ | v_1__30_;
  assign addr_3__24_ = addr_2__24_ | addr_2__28_;
  assign v_3__32_ = v_2__36_ | v_2__32_;
  assign addr_3__33_ = v_1__34_ | v_1__38_;
  assign addr_3__32_ = addr_2__32_ | addr_2__36_;
  assign v_3__40_ = v_2__44_ | v_2__40_;
  assign addr_3__41_ = v_1__42_ | v_1__46_;
  assign addr_3__40_ = addr_2__40_ | addr_2__44_;
  assign v_3__48_ = v_2__52_ | v_2__48_;
  assign addr_3__49_ = v_1__50_ | v_1__54_;
  assign addr_3__48_ = addr_2__48_ | addr_2__52_;
  assign v_3__56_ = v_2__60_ | v_2__56_;
  assign addr_3__57_ = v_1__58_ | v_1__62_;
  assign addr_3__56_ = addr_2__56_ | addr_2__60_;
  assign v_3__64_ = v_2__68_ | v_2__64_;
  assign addr_3__65_ = v_1__66_ | v_1__70_;
  assign addr_3__64_ = addr_2__64_ | addr_2__68_;
  assign v_3__72_ = v_2__76_ | v_2__72_;
  assign addr_3__73_ = v_1__74_ | v_1__78_;
  assign addr_3__72_ = addr_2__72_ | addr_2__76_;
  assign v_3__80_ = v_2__84_ | v_2__80_;
  assign addr_3__81_ = v_1__82_ | v_1__86_;
  assign addr_3__80_ = addr_2__80_ | addr_2__84_;
  assign v_3__88_ = v_2__92_ | v_2__88_;
  assign addr_3__89_ = v_1__90_ | v_1__94_;
  assign addr_3__88_ = addr_2__88_ | addr_2__92_;
  assign v_3__96_ = v_2__100_ | v_2__96_;
  assign addr_3__97_ = v_1__98_ | v_1__102_;
  assign addr_3__96_ = addr_2__96_ | addr_2__100_;
  assign v_3__104_ = v_2__108_ | v_2__104_;
  assign addr_3__105_ = v_1__106_ | v_1__110_;
  assign addr_3__104_ = addr_2__104_ | addr_2__108_;
  assign v_3__112_ = v_2__116_ | v_2__112_;
  assign addr_3__113_ = v_1__114_ | v_1__118_;
  assign addr_3__112_ = addr_2__112_ | addr_2__116_;
  assign v_3__120_ = v_2__124_ | v_2__120_;
  assign addr_3__121_ = v_1__122_ | v_1__126_;
  assign addr_3__120_ = addr_2__120_ | addr_2__124_;
  assign v_4__0_ = v_3__8_ | v_3__0_;
  assign addr_4__2_ = v_2__4_ | v_2__12_;
  assign addr_4__1_ = addr_3__1_ | addr_3__9_;
  assign addr_4__0_ = addr_3__0_ | addr_3__8_;
  assign v_4__16_ = v_3__24_ | v_3__16_;
  assign addr_4__18_ = v_2__20_ | v_2__28_;
  assign addr_4__17_ = addr_3__17_ | addr_3__25_;
  assign addr_4__16_ = addr_3__16_ | addr_3__24_;
  assign v_4__32_ = v_3__40_ | v_3__32_;
  assign addr_4__34_ = v_2__36_ | v_2__44_;
  assign addr_4__33_ = addr_3__33_ | addr_3__41_;
  assign addr_4__32_ = addr_3__32_ | addr_3__40_;
  assign v_4__48_ = v_3__56_ | v_3__48_;
  assign addr_4__50_ = v_2__52_ | v_2__60_;
  assign addr_4__49_ = addr_3__49_ | addr_3__57_;
  assign addr_4__48_ = addr_3__48_ | addr_3__56_;
  assign v_4__64_ = v_3__72_ | v_3__64_;
  assign addr_4__66_ = v_2__68_ | v_2__76_;
  assign addr_4__65_ = addr_3__65_ | addr_3__73_;
  assign addr_4__64_ = addr_3__64_ | addr_3__72_;
  assign v_4__80_ = v_3__88_ | v_3__80_;
  assign addr_4__82_ = v_2__84_ | v_2__92_;
  assign addr_4__81_ = addr_3__81_ | addr_3__89_;
  assign addr_4__80_ = addr_3__80_ | addr_3__88_;
  assign v_4__96_ = v_3__104_ | v_3__96_;
  assign addr_4__98_ = v_2__100_ | v_2__108_;
  assign addr_4__97_ = addr_3__97_ | addr_3__105_;
  assign addr_4__96_ = addr_3__96_ | addr_3__104_;
  assign v_4__112_ = v_3__120_ | v_3__112_;
  assign addr_4__114_ = v_2__116_ | v_2__124_;
  assign addr_4__113_ = addr_3__113_ | addr_3__121_;
  assign addr_4__112_ = addr_3__112_ | addr_3__120_;
  assign v_5__0_ = v_4__16_ | v_4__0_;
  assign addr_5__3_ = v_3__8_ | v_3__24_;
  assign addr_5__2_ = addr_4__2_ | addr_4__18_;
  assign addr_5__1_ = addr_4__1_ | addr_4__17_;
  assign addr_5__0_ = addr_4__0_ | addr_4__16_;
  assign v_5__32_ = v_4__48_ | v_4__32_;
  assign addr_5__35_ = v_3__40_ | v_3__56_;
  assign addr_5__34_ = addr_4__34_ | addr_4__50_;
  assign addr_5__33_ = addr_4__33_ | addr_4__49_;
  assign addr_5__32_ = addr_4__32_ | addr_4__48_;
  assign v_5__64_ = v_4__80_ | v_4__64_;
  assign addr_5__67_ = v_3__72_ | v_3__88_;
  assign addr_5__66_ = addr_4__66_ | addr_4__82_;
  assign addr_5__65_ = addr_4__65_ | addr_4__81_;
  assign addr_5__64_ = addr_4__64_ | addr_4__80_;
  assign v_5__96_ = v_4__112_ | v_4__96_;
  assign addr_5__99_ = v_3__104_ | v_3__120_;
  assign addr_5__98_ = addr_4__98_ | addr_4__114_;
  assign addr_5__97_ = addr_4__97_ | addr_4__113_;
  assign addr_5__96_ = addr_4__96_ | addr_4__112_;
  assign v_6__0_ = v_5__32_ | v_5__0_;
  assign addr_6__4_ = v_4__16_ | v_4__48_;
  assign addr_6__3_ = addr_5__3_ | addr_5__35_;
  assign addr_6__2_ = addr_5__2_ | addr_5__34_;
  assign addr_6__1_ = addr_5__1_ | addr_5__33_;
  assign addr_6__0_ = addr_5__0_ | addr_5__32_;
  assign addr_o[6] = v_5__96_ | v_5__64_;
  assign addr_6__68_ = v_4__80_ | v_4__112_;
  assign addr_6__67_ = addr_5__67_ | addr_5__99_;
  assign addr_6__66_ = addr_5__66_ | addr_5__98_;
  assign addr_6__65_ = addr_5__65_ | addr_5__97_;
  assign addr_6__64_ = addr_5__64_ | addr_5__96_;
  assign v_o = addr_o[6] | v_6__0_;
  assign addr_o[5] = v_5__32_ | v_5__96_;
  assign addr_o[4] = addr_6__4_ | addr_6__68_;
  assign addr_o[3] = addr_6__3_ | addr_6__67_;
  assign addr_o[2] = addr_6__2_ | addr_6__66_;
  assign addr_o[1] = addr_6__1_ | addr_6__65_;
  assign addr_o[0] = addr_6__0_ | addr_6__64_;

endmodule



module bsg_priority_encode_width_p65_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [64:0] i;
  output [6:0] addr_o;
  output v_o;
  wire [6:0] addr_o;
  wire v_o;
  wire [64:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p65_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_width_p65_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o)
  );


endmodule



module bsg_counting_leading_zeros_width_p64
(
  a_i,
  num_zero_o
);

  input [63:0] a_i;
  output [6:0] num_zero_o;
  wire [6:0] num_zero_o;

  bsg_priority_encode_width_p65_lo_to_hi_p1
  pe0
  (
    .i({ 1'b1, a_i[0:0], a_i[1:1], a_i[2:2], a_i[3:3], a_i[4:4], a_i[5:5], a_i[6:6], a_i[7:7], a_i[8:8], a_i[9:9], a_i[10:10], a_i[11:11], a_i[12:12], a_i[13:13], a_i[14:14], a_i[15:15], a_i[16:16], a_i[17:17], a_i[18:18], a_i[19:19], a_i[20:20], a_i[21:21], a_i[22:22], a_i[23:23], a_i[24:24], a_i[25:25], a_i[26:26], a_i[27:27], a_i[28:28], a_i[29:29], a_i[30:30], a_i[31:31], a_i[32:32], a_i[33:33], a_i[34:34], a_i[35:35], a_i[36:36], a_i[37:37], a_i[38:38], a_i[39:39], a_i[40:40], a_i[41:41], a_i[42:42], a_i[43:43], a_i[44:44], a_i[45:45], a_i[46:46], a_i[47:47], a_i[48:48], a_i[49:49], a_i[50:50], a_i[51:51], a_i[52:52], a_i[53:53], a_i[54:54], a_i[55:55], a_i[56:56], a_i[57:57], a_i[58:58], a_i[59:59], a_i[60:60], a_i[61:61], a_i[62:62], a_i[63:63] }),
    .addr_o(num_zero_o)
  );


endmodule



module iNToRawFN_intWidth64
(
  signedIn,
  in,
  isZero,
  sign,
  sExp,
  sig
);

  input [63:0] in;
  output [8:0] sExp;
  output [64:0] sig;
  input signedIn;
  output isZero;
  output sign;
  wire [8:0] sExp;
  wire [64:0] sig;
  wire isZero,sign,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66;
  wire [63:0] absIn;
  wire [6:0] num_zero_lo;
  assign sExp[7] = 1'b1;
  assign sExp[6] = 1'b0;
  assign sExp[8] = 1'b0;

  bsg_counting_leading_zeros_width_p64
  clz
  (
    .a_i(absIn),
    .num_zero_o(num_zero_lo)
  );

  assign sig = { 1'b0, absIn } << num_zero_lo[5:0];
  assign { N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3 } = 1'b0 - in;
  assign absIn = (N0)? { N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3 } : 
                 (N1)? in : 1'b0;
  assign N0 = sign;
  assign N1 = N2;
  assign sign = signedIn & in[63];
  assign N2 = ~sign;
  assign isZero = ~sig[63];
  assign sExp[5] = ~num_zero_lo[5];
  assign sExp[4] = ~num_zero_lo[4];
  assign sExp[3] = ~num_zero_lo[3];
  assign sExp[2] = ~num_zero_lo[2];
  assign sExp[1] = ~num_zero_lo[1];
  assign sExp[0] = ~num_zero_lo[0];

endmodule



module roundAnyRawFNToRecFN_inExpWidth7_inSigWidth64_outExpWidth11_outSigWidth53_options5
(
  control,
  invalidExc,
  infiniteExc,
  in_isNaN,
  in_isInf,
  in_isZero,
  in_sign,
  in_sExp,
  in_sig,
  roundingMode,
  out,
  exceptionFlags
);

  input [0:0] control;
  input [8:0] in_sExp;
  input [64:0] in_sig;
  input [2:0] roundingMode;
  output [64:0] out;
  output [4:0] exceptionFlags;
  input invalidExc;
  input infiniteExc;
  input in_isNaN;
  input in_isInf;
  input in_isZero;
  input in_sign;
  wire [64:0] out;
  wire [4:0] exceptionFlags;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,exceptionFlags_4_,exceptionFlags_3_,roundMagUp,
  isNaNOut,\genblk2.roundPosBit ,\genblk2.anyRoundExtra ,\genblk2.anyRound ,
  \genblk2.roundIncr ,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,
  N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,
  N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
  N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,
  N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,
  N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,
  N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,
  N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,
  N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,
  N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,
  N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,
  N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,
  N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,
  N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,
  N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,
  N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,
  N281,N282,N283,N284,N285,common_inexact,notNaN_isSpecialInfOut,commonCase,
  overflow_roundMagUp,pegMinNonzeroMagOut,pegMaxFiniteMagOut,notNaN_isInfOut,N286,N287,N288,
  N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,
  N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,
  N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
  N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,
  N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
  N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,
  N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,
  N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,
  N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,
  N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,
  N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,
  N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,
  N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,
  N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,
  N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,
  N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,
  N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,
  N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,
  N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,
  N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,
  N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,
  N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,
  N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,
  N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,
  N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,
  N689,N690,N691,N692,N693;
  wire [11:0] sAdjustedExp,\genblk2.sRoundedExp ;
  wire [0:0] adjustedSig;
  wire [55:0] \genblk2.roundPosMask ;
  wire [54:0] \genblk2.roundedSig ;
  wire [51:0] common_fractOut;
  assign exceptionFlags_4_ = invalidExc;
  assign exceptionFlags[4] = exceptionFlags_4_;
  assign exceptionFlags_3_ = infiniteExc;
  assign exceptionFlags[3] = exceptionFlags_3_;
  assign N343 = ~roundingMode[2];
  assign N344 = roundingMode[1] | N343;
  assign N345 = roundingMode[0] | N344;
  assign N346 = ~N345;
  assign N347 = roundingMode[1] | roundingMode[2];
  assign N348 = roundingMode[0] | N347;
  assign N349 = ~N348;
  assign N350 = ~roundingMode[1];
  assign N351 = N350 | N343;
  assign N352 = roundingMode[0] | N351;
  assign N353 = ~N352;
  assign N354 = N350 | roundingMode[2];
  assign N355 = roundingMode[0] | N354;
  assign N356 = ~N355;
  assign N357 = ~roundingMode[0];
  assign N358 = N357 | N354;
  assign N359 = ~N358;
  assign sAdjustedExp = $signed(in_sExp) + $signed({ 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 });
  assign { N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65 } = { N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64 } + 1'b1;
  assign \genblk2.sRoundedExp  = sAdjustedExp + \genblk2.roundedSig [54:53];
  assign { N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177 } = (N0)? \genblk2.roundPosMask [55:1] : 
                                                                                                                                                                                                                                                                                                                                                        (N176)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N175;
  assign \genblk2.roundedSig  = (N1)? { N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174 } : 
                                (N2)? { N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285 } : 1'b0;
  assign N1 = \genblk2.roundIncr ;
  assign N2 = N9;
  assign common_fractOut = (N3)? \genblk2.roundedSig [52:1] : 
                           (N4)? \genblk2.roundedSig [51:0] : 1'b0;
  assign N3 = 1'b0;
  assign N4 = N373;
  assign out[64] = (N5)? 1'b0 : 
                   (N6)? in_sign : 1'b0;
  assign N5 = isNaNOut;
  assign N6 = N657;
  assign N289 = (N7)? common_fractOut[51] : 
                (N288)? 1'b0 : 1'b0;
  assign N7 = N287;
  assign { N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292 } = (N8)? common_fractOut[50:0] : 
                                                                                                                                                                                                                                                                                                                                (N291)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = N290;
  assign roundMagUp = N360 | N362;
  assign N360 = N356 & in_sign;
  assign N362 = N359 & N361;
  assign N361 = ~in_sign;
  assign isNaNOut = exceptionFlags_4_ | N364;
  assign N364 = N363 & in_isNaN;
  assign N363 = ~exceptionFlags_3_;
  assign adjustedSig[0] = N372 | in_sig[0];
  assign N372 = N371 | in_sig[1];
  assign N371 = N370 | in_sig[2];
  assign N370 = N369 | in_sig[3];
  assign N369 = N368 | in_sig[4];
  assign N368 = N367 | in_sig[5];
  assign N367 = N366 | in_sig[6];
  assign N366 = N365 | in_sig[7];
  assign N365 = in_sig[9] | in_sig[8];
  assign \genblk2.roundPosMask [55] = N373 & 1'b0;
  assign N373 = ~1'b0;
  assign \genblk2.roundPosMask [54] = N373 & 1'b0;
  assign \genblk2.roundPosMask [53] = N373 & 1'b0;
  assign \genblk2.roundPosMask [52] = N373 & 1'b0;
  assign \genblk2.roundPosMask [51] = N373 & 1'b0;
  assign \genblk2.roundPosMask [50] = N373 & 1'b0;
  assign \genblk2.roundPosMask [49] = N373 & 1'b0;
  assign \genblk2.roundPosMask [48] = N373 & 1'b0;
  assign \genblk2.roundPosMask [47] = N373 & 1'b0;
  assign \genblk2.roundPosMask [46] = N373 & 1'b0;
  assign \genblk2.roundPosMask [45] = N373 & 1'b0;
  assign \genblk2.roundPosMask [44] = N373 & 1'b0;
  assign \genblk2.roundPosMask [43] = N373 & 1'b0;
  assign \genblk2.roundPosMask [42] = N373 & 1'b0;
  assign \genblk2.roundPosMask [41] = N373 & 1'b0;
  assign \genblk2.roundPosMask [40] = N373 & 1'b0;
  assign \genblk2.roundPosMask [39] = N373 & 1'b0;
  assign \genblk2.roundPosMask [38] = N373 & 1'b0;
  assign \genblk2.roundPosMask [37] = N373 & 1'b0;
  assign \genblk2.roundPosMask [36] = N373 & 1'b0;
  assign \genblk2.roundPosMask [35] = N373 & 1'b0;
  assign \genblk2.roundPosMask [34] = N373 & 1'b0;
  assign \genblk2.roundPosMask [33] = N373 & 1'b0;
  assign \genblk2.roundPosMask [32] = N373 & 1'b0;
  assign \genblk2.roundPosMask [31] = N373 & 1'b0;
  assign \genblk2.roundPosMask [30] = N373 & 1'b0;
  assign \genblk2.roundPosMask [29] = N373 & 1'b0;
  assign \genblk2.roundPosMask [28] = N373 & 1'b0;
  assign \genblk2.roundPosMask [27] = N373 & 1'b0;
  assign \genblk2.roundPosMask [26] = N373 & 1'b0;
  assign \genblk2.roundPosMask [25] = N373 & 1'b0;
  assign \genblk2.roundPosMask [24] = N373 & 1'b0;
  assign \genblk2.roundPosMask [23] = N373 & 1'b0;
  assign \genblk2.roundPosMask [22] = N373 & 1'b0;
  assign \genblk2.roundPosMask [21] = N373 & 1'b0;
  assign \genblk2.roundPosMask [20] = N373 & 1'b0;
  assign \genblk2.roundPosMask [19] = N373 & 1'b0;
  assign \genblk2.roundPosMask [18] = N373 & 1'b0;
  assign \genblk2.roundPosMask [17] = N373 & 1'b0;
  assign \genblk2.roundPosMask [16] = N373 & 1'b0;
  assign \genblk2.roundPosMask [15] = N373 & 1'b0;
  assign \genblk2.roundPosMask [14] = N373 & 1'b0;
  assign \genblk2.roundPosMask [13] = N373 & 1'b0;
  assign \genblk2.roundPosMask [12] = N373 & 1'b0;
  assign \genblk2.roundPosMask [11] = N373 & 1'b0;
  assign \genblk2.roundPosMask [10] = N373 & 1'b0;
  assign \genblk2.roundPosMask [9] = N373 & 1'b0;
  assign \genblk2.roundPosMask [8] = N373 & 1'b0;
  assign \genblk2.roundPosMask [7] = N373 & 1'b0;
  assign \genblk2.roundPosMask [6] = N373 & 1'b0;
  assign \genblk2.roundPosMask [5] = N373 & 1'b0;
  assign \genblk2.roundPosMask [4] = N373 & 1'b0;
  assign \genblk2.roundPosMask [3] = N373 & 1'b0;
  assign \genblk2.roundPosMask [2] = N373 & 1'b0;
  assign \genblk2.roundPosMask [1] = N373 & 1'b1;
  assign \genblk2.roundPosMask [0] = N374 & 1'b1;
  assign N374 = ~1'b1;
  assign \genblk2.roundPosBit  = N479 | N485;
  assign N479 = N477 | N478;
  assign N477 = N475 | N476;
  assign N475 = N473 | N474;
  assign N473 = N471 | N472;
  assign N471 = N469 | N470;
  assign N469 = N467 | N468;
  assign N467 = N465 | N466;
  assign N465 = N463 | N464;
  assign N463 = N461 | N462;
  assign N461 = N459 | N460;
  assign N459 = N457 | N458;
  assign N457 = N455 | N456;
  assign N455 = N453 | N454;
  assign N453 = N451 | N452;
  assign N451 = N449 | N450;
  assign N449 = N447 | N448;
  assign N447 = N445 | N446;
  assign N445 = N443 | N444;
  assign N443 = N441 | N442;
  assign N441 = N439 | N440;
  assign N439 = N437 | N438;
  assign N437 = N435 | N436;
  assign N435 = N433 | N434;
  assign N433 = N431 | N432;
  assign N431 = N429 | N430;
  assign N429 = N427 | N428;
  assign N427 = N425 | N426;
  assign N425 = N423 | N424;
  assign N423 = N421 | N422;
  assign N421 = N419 | N420;
  assign N419 = N417 | N418;
  assign N417 = N415 | N416;
  assign N415 = N413 | N414;
  assign N413 = N411 | N412;
  assign N411 = N409 | N410;
  assign N409 = N407 | N408;
  assign N407 = N405 | N406;
  assign N405 = N403 | N404;
  assign N403 = N401 | N402;
  assign N401 = N399 | N400;
  assign N399 = N397 | N398;
  assign N397 = N395 | N396;
  assign N395 = N393 | N394;
  assign N393 = N391 | N392;
  assign N391 = N389 | N390;
  assign N389 = N387 | N388;
  assign N387 = N385 | N386;
  assign N385 = N383 | N384;
  assign N383 = N381 | N382;
  assign N381 = N379 | N380;
  assign N379 = N377 | N378;
  assign N377 = N375 | N376;
  assign N375 = in_sig[64] & \genblk2.roundPosMask [55];
  assign N376 = in_sig[63] & \genblk2.roundPosMask [54];
  assign N378 = in_sig[62] & \genblk2.roundPosMask [53];
  assign N380 = in_sig[61] & \genblk2.roundPosMask [52];
  assign N382 = in_sig[60] & \genblk2.roundPosMask [51];
  assign N384 = in_sig[59] & \genblk2.roundPosMask [50];
  assign N386 = in_sig[58] & \genblk2.roundPosMask [49];
  assign N388 = in_sig[57] & \genblk2.roundPosMask [48];
  assign N390 = in_sig[56] & \genblk2.roundPosMask [47];
  assign N392 = in_sig[55] & \genblk2.roundPosMask [46];
  assign N394 = in_sig[54] & \genblk2.roundPosMask [45];
  assign N396 = in_sig[53] & \genblk2.roundPosMask [44];
  assign N398 = in_sig[52] & \genblk2.roundPosMask [43];
  assign N400 = in_sig[51] & \genblk2.roundPosMask [42];
  assign N402 = in_sig[50] & \genblk2.roundPosMask [41];
  assign N404 = in_sig[49] & \genblk2.roundPosMask [40];
  assign N406 = in_sig[48] & \genblk2.roundPosMask [39];
  assign N408 = in_sig[47] & \genblk2.roundPosMask [38];
  assign N410 = in_sig[46] & \genblk2.roundPosMask [37];
  assign N412 = in_sig[45] & \genblk2.roundPosMask [36];
  assign N414 = in_sig[44] & \genblk2.roundPosMask [35];
  assign N416 = in_sig[43] & \genblk2.roundPosMask [34];
  assign N418 = in_sig[42] & \genblk2.roundPosMask [33];
  assign N420 = in_sig[41] & \genblk2.roundPosMask [32];
  assign N422 = in_sig[40] & \genblk2.roundPosMask [31];
  assign N424 = in_sig[39] & \genblk2.roundPosMask [30];
  assign N426 = in_sig[38] & \genblk2.roundPosMask [29];
  assign N428 = in_sig[37] & \genblk2.roundPosMask [28];
  assign N430 = in_sig[36] & \genblk2.roundPosMask [27];
  assign N432 = in_sig[35] & \genblk2.roundPosMask [26];
  assign N434 = in_sig[34] & \genblk2.roundPosMask [25];
  assign N436 = in_sig[33] & \genblk2.roundPosMask [24];
  assign N438 = in_sig[32] & \genblk2.roundPosMask [23];
  assign N440 = in_sig[31] & \genblk2.roundPosMask [22];
  assign N442 = in_sig[30] & \genblk2.roundPosMask [21];
  assign N444 = in_sig[29] & \genblk2.roundPosMask [20];
  assign N446 = in_sig[28] & \genblk2.roundPosMask [19];
  assign N448 = in_sig[27] & \genblk2.roundPosMask [18];
  assign N450 = in_sig[26] & \genblk2.roundPosMask [17];
  assign N452 = in_sig[25] & \genblk2.roundPosMask [16];
  assign N454 = in_sig[24] & \genblk2.roundPosMask [15];
  assign N456 = in_sig[23] & \genblk2.roundPosMask [14];
  assign N458 = in_sig[22] & \genblk2.roundPosMask [13];
  assign N460 = in_sig[21] & \genblk2.roundPosMask [12];
  assign N462 = in_sig[20] & \genblk2.roundPosMask [11];
  assign N464 = in_sig[19] & \genblk2.roundPosMask [10];
  assign N466 = in_sig[18] & \genblk2.roundPosMask [9];
  assign N468 = in_sig[17] & \genblk2.roundPosMask [8];
  assign N470 = in_sig[16] & \genblk2.roundPosMask [7];
  assign N472 = in_sig[15] & \genblk2.roundPosMask [6];
  assign N474 = in_sig[14] & \genblk2.roundPosMask [5];
  assign N476 = in_sig[13] & \genblk2.roundPosMask [4];
  assign N478 = in_sig[12] & \genblk2.roundPosMask [3];
  assign N485 = N484 & N373;
  assign N484 = N482 | N483;
  assign N482 = N480 | N481;
  assign N480 = in_sig[11] & \genblk2.roundPosMask [2];
  assign N481 = in_sig[10] & \genblk2.roundPosMask [1];
  assign N483 = adjustedSig[0] & \genblk2.roundPosMask [0];
  assign \genblk2.anyRoundExtra  = N590 | N596;
  assign N590 = N588 | N589;
  assign N588 = N586 | N587;
  assign N586 = N584 | N585;
  assign N584 = N582 | N583;
  assign N582 = N580 | N581;
  assign N580 = N578 | N579;
  assign N578 = N576 | N577;
  assign N576 = N574 | N575;
  assign N574 = N572 | N573;
  assign N572 = N570 | N571;
  assign N570 = N568 | N569;
  assign N568 = N566 | N567;
  assign N566 = N564 | N565;
  assign N564 = N562 | N563;
  assign N562 = N560 | N561;
  assign N560 = N558 | N559;
  assign N558 = N556 | N557;
  assign N556 = N554 | N555;
  assign N554 = N552 | N553;
  assign N552 = N550 | N551;
  assign N550 = N548 | N549;
  assign N548 = N546 | N547;
  assign N546 = N544 | N545;
  assign N544 = N542 | N543;
  assign N542 = N540 | N541;
  assign N540 = N538 | N539;
  assign N538 = N536 | N537;
  assign N536 = N534 | N535;
  assign N534 = N532 | N533;
  assign N532 = N530 | N531;
  assign N530 = N528 | N529;
  assign N528 = N526 | N527;
  assign N526 = N524 | N525;
  assign N524 = N522 | N523;
  assign N522 = N520 | N521;
  assign N520 = N518 | N519;
  assign N518 = N516 | N517;
  assign N516 = N514 | N515;
  assign N514 = N512 | N513;
  assign N512 = N510 | N511;
  assign N510 = N508 | N509;
  assign N508 = N506 | N507;
  assign N506 = N504 | N505;
  assign N504 = N502 | N503;
  assign N502 = N500 | N501;
  assign N500 = N498 | N499;
  assign N498 = N496 | N497;
  assign N496 = N494 | N495;
  assign N494 = N492 | N493;
  assign N492 = N490 | N491;
  assign N490 = N488 | N489;
  assign N488 = N486 | N487;
  assign N486 = in_sig[64] & 1'b0;
  assign N487 = in_sig[63] & 1'b0;
  assign N489 = in_sig[62] & 1'b0;
  assign N491 = in_sig[61] & 1'b0;
  assign N493 = in_sig[60] & 1'b0;
  assign N495 = in_sig[59] & 1'b0;
  assign N497 = in_sig[58] & 1'b0;
  assign N499 = in_sig[57] & 1'b0;
  assign N501 = in_sig[56] & 1'b0;
  assign N503 = in_sig[55] & 1'b0;
  assign N505 = in_sig[54] & 1'b0;
  assign N507 = in_sig[53] & 1'b0;
  assign N509 = in_sig[52] & 1'b0;
  assign N511 = in_sig[51] & 1'b0;
  assign N513 = in_sig[50] & 1'b0;
  assign N515 = in_sig[49] & 1'b0;
  assign N517 = in_sig[48] & 1'b0;
  assign N519 = in_sig[47] & 1'b0;
  assign N521 = in_sig[46] & 1'b0;
  assign N523 = in_sig[45] & 1'b0;
  assign N525 = in_sig[44] & 1'b0;
  assign N527 = in_sig[43] & 1'b0;
  assign N529 = in_sig[42] & 1'b0;
  assign N531 = in_sig[41] & 1'b0;
  assign N533 = in_sig[40] & 1'b0;
  assign N535 = in_sig[39] & 1'b0;
  assign N537 = in_sig[38] & 1'b0;
  assign N539 = in_sig[37] & 1'b0;
  assign N541 = in_sig[36] & 1'b0;
  assign N543 = in_sig[35] & 1'b0;
  assign N545 = in_sig[34] & 1'b0;
  assign N547 = in_sig[33] & 1'b0;
  assign N549 = in_sig[32] & 1'b0;
  assign N551 = in_sig[31] & 1'b0;
  assign N553 = in_sig[30] & 1'b0;
  assign N555 = in_sig[29] & 1'b0;
  assign N557 = in_sig[28] & 1'b0;
  assign N559 = in_sig[27] & 1'b0;
  assign N561 = in_sig[26] & 1'b0;
  assign N563 = in_sig[25] & 1'b0;
  assign N565 = in_sig[24] & 1'b0;
  assign N567 = in_sig[23] & 1'b0;
  assign N569 = in_sig[22] & 1'b0;
  assign N571 = in_sig[21] & 1'b0;
  assign N573 = in_sig[20] & 1'b0;
  assign N575 = in_sig[19] & 1'b0;
  assign N577 = in_sig[18] & 1'b0;
  assign N579 = in_sig[17] & 1'b0;
  assign N581 = in_sig[16] & 1'b0;
  assign N583 = in_sig[15] & 1'b0;
  assign N585 = in_sig[14] & 1'b0;
  assign N587 = in_sig[13] & 1'b0;
  assign N589 = in_sig[12] & 1'b0;
  assign N596 = N595 & N373;
  assign N595 = N593 | N594;
  assign N593 = N591 | N592;
  assign N591 = in_sig[11] & 1'b0;
  assign N592 = in_sig[10] & 1'b0;
  assign N594 = adjustedSig[0] & 1'b1;
  assign \genblk2.anyRound  = \genblk2.roundPosBit  | \genblk2.anyRoundExtra ;
  assign \genblk2.roundIncr  = N598 | N599;
  assign N598 = N597 & \genblk2.roundPosBit ;
  assign N597 = N349 | N346;
  assign N599 = roundMagUp & \genblk2.anyRound ;
  assign N9 = ~\genblk2.roundIncr ;
  assign N10 = N600 & N601;
  assign N600 = N349 & \genblk2.roundPosBit ;
  assign N601 = ~\genblk2.anyRoundExtra ;
  assign N11 = in_sig[64] | 1'b0;
  assign N12 = in_sig[63] | 1'b0;
  assign N13 = in_sig[62] | 1'b0;
  assign N14 = in_sig[61] | 1'b0;
  assign N15 = in_sig[60] | 1'b0;
  assign N16 = in_sig[59] | 1'b0;
  assign N17 = in_sig[58] | 1'b0;
  assign N18 = in_sig[57] | 1'b0;
  assign N19 = in_sig[56] | 1'b0;
  assign N20 = in_sig[55] | 1'b0;
  assign N21 = in_sig[54] | 1'b0;
  assign N22 = in_sig[53] | 1'b0;
  assign N23 = in_sig[52] | 1'b0;
  assign N24 = in_sig[51] | 1'b0;
  assign N25 = in_sig[50] | 1'b0;
  assign N26 = in_sig[49] | 1'b0;
  assign N27 = in_sig[48] | 1'b0;
  assign N28 = in_sig[47] | 1'b0;
  assign N29 = in_sig[46] | 1'b0;
  assign N30 = in_sig[45] | 1'b0;
  assign N31 = in_sig[44] | 1'b0;
  assign N32 = in_sig[43] | 1'b0;
  assign N33 = in_sig[42] | 1'b0;
  assign N34 = in_sig[41] | 1'b0;
  assign N35 = in_sig[40] | 1'b0;
  assign N36 = in_sig[39] | 1'b0;
  assign N37 = in_sig[38] | 1'b0;
  assign N38 = in_sig[37] | 1'b0;
  assign N39 = in_sig[36] | 1'b0;
  assign N40 = in_sig[35] | 1'b0;
  assign N41 = in_sig[34] | 1'b0;
  assign N42 = in_sig[33] | 1'b0;
  assign N43 = in_sig[32] | 1'b0;
  assign N44 = in_sig[31] | 1'b0;
  assign N45 = in_sig[30] | 1'b0;
  assign N46 = in_sig[29] | 1'b0;
  assign N47 = in_sig[28] | 1'b0;
  assign N48 = in_sig[27] | 1'b0;
  assign N49 = in_sig[26] | 1'b0;
  assign N50 = in_sig[25] | 1'b0;
  assign N51 = in_sig[24] | 1'b0;
  assign N52 = in_sig[23] | 1'b0;
  assign N53 = in_sig[22] | 1'b0;
  assign N54 = in_sig[21] | 1'b0;
  assign N55 = in_sig[20] | 1'b0;
  assign N56 = in_sig[19] | 1'b0;
  assign N57 = in_sig[18] | 1'b0;
  assign N58 = in_sig[17] | 1'b0;
  assign N59 = in_sig[16] | 1'b0;
  assign N60 = in_sig[15] | 1'b0;
  assign N61 = in_sig[14] | 1'b0;
  assign N62 = in_sig[13] | 1'b0;
  assign N63 = in_sig[12] | 1'b0;
  assign N64 = in_sig[11] | 1'b0;
  assign N120 = N119 & N373;
  assign N121 = N118 & N373;
  assign N122 = N117 & N373;
  assign N123 = N116 & N373;
  assign N124 = N115 & N373;
  assign N125 = N114 & N373;
  assign N126 = N113 & N373;
  assign N127 = N112 & N373;
  assign N128 = N111 & N373;
  assign N129 = N110 & N373;
  assign N130 = N109 & N373;
  assign N131 = N108 & N373;
  assign N132 = N107 & N373;
  assign N133 = N106 & N373;
  assign N134 = N105 & N373;
  assign N135 = N104 & N373;
  assign N136 = N103 & N373;
  assign N137 = N102 & N373;
  assign N138 = N101 & N373;
  assign N139 = N100 & N373;
  assign N140 = N99 & N373;
  assign N141 = N98 & N373;
  assign N142 = N97 & N373;
  assign N143 = N96 & N373;
  assign N144 = N95 & N373;
  assign N145 = N94 & N373;
  assign N146 = N93 & N373;
  assign N147 = N92 & N373;
  assign N148 = N91 & N373;
  assign N149 = N90 & N373;
  assign N150 = N89 & N373;
  assign N151 = N88 & N373;
  assign N152 = N87 & N373;
  assign N153 = N86 & N373;
  assign N154 = N85 & N373;
  assign N155 = N84 & N373;
  assign N156 = N83 & N373;
  assign N157 = N82 & N373;
  assign N158 = N81 & N373;
  assign N159 = N80 & N373;
  assign N160 = N79 & N373;
  assign N161 = N78 & N373;
  assign N162 = N77 & N373;
  assign N163 = N76 & N373;
  assign N164 = N75 & N373;
  assign N165 = N74 & N373;
  assign N166 = N73 & N373;
  assign N167 = N72 & N373;
  assign N168 = N71 & N373;
  assign N169 = N70 & N373;
  assign N170 = N69 & N373;
  assign N171 = N68 & N373;
  assign N172 = N67 & N373;
  assign N173 = N66 & N373;
  assign N174 = N65 & N602;
  assign N602 = ~N10;
  assign N175 = N353 & \genblk2.anyRound ;
  assign N176 = ~N175;
  assign N232 = N603 | N230;
  assign N603 = in_sig[64] & N373;
  assign N233 = N604 | N229;
  assign N604 = in_sig[63] & N373;
  assign N234 = N605 | N228;
  assign N605 = in_sig[62] & N373;
  assign N235 = N606 | N227;
  assign N606 = in_sig[61] & N373;
  assign N236 = N607 | N226;
  assign N607 = in_sig[60] & N373;
  assign N237 = N608 | N225;
  assign N608 = in_sig[59] & N373;
  assign N238 = N609 | N224;
  assign N609 = in_sig[58] & N373;
  assign N239 = N610 | N223;
  assign N610 = in_sig[57] & N373;
  assign N240 = N611 | N222;
  assign N611 = in_sig[56] & N373;
  assign N241 = N612 | N221;
  assign N612 = in_sig[55] & N373;
  assign N242 = N613 | N220;
  assign N613 = in_sig[54] & N373;
  assign N243 = N614 | N219;
  assign N614 = in_sig[53] & N373;
  assign N244 = N615 | N218;
  assign N615 = in_sig[52] & N373;
  assign N245 = N616 | N217;
  assign N616 = in_sig[51] & N373;
  assign N246 = N617 | N216;
  assign N617 = in_sig[50] & N373;
  assign N247 = N618 | N215;
  assign N618 = in_sig[49] & N373;
  assign N248 = N619 | N214;
  assign N619 = in_sig[48] & N373;
  assign N249 = N620 | N213;
  assign N620 = in_sig[47] & N373;
  assign N250 = N621 | N212;
  assign N621 = in_sig[46] & N373;
  assign N251 = N622 | N211;
  assign N622 = in_sig[45] & N373;
  assign N252 = N623 | N210;
  assign N623 = in_sig[44] & N373;
  assign N253 = N624 | N209;
  assign N624 = in_sig[43] & N373;
  assign N254 = N625 | N208;
  assign N625 = in_sig[42] & N373;
  assign N255 = N626 | N207;
  assign N626 = in_sig[41] & N373;
  assign N256 = N627 | N206;
  assign N627 = in_sig[40] & N373;
  assign N257 = N628 | N205;
  assign N628 = in_sig[39] & N373;
  assign N258 = N629 | N204;
  assign N629 = in_sig[38] & N373;
  assign N259 = N630 | N203;
  assign N630 = in_sig[37] & N373;
  assign N260 = N631 | N202;
  assign N631 = in_sig[36] & N373;
  assign N261 = N632 | N201;
  assign N632 = in_sig[35] & N373;
  assign N262 = N633 | N200;
  assign N633 = in_sig[34] & N373;
  assign N263 = N634 | N199;
  assign N634 = in_sig[33] & N373;
  assign N264 = N635 | N198;
  assign N635 = in_sig[32] & N373;
  assign N265 = N636 | N197;
  assign N636 = in_sig[31] & N373;
  assign N266 = N637 | N196;
  assign N637 = in_sig[30] & N373;
  assign N267 = N638 | N195;
  assign N638 = in_sig[29] & N373;
  assign N268 = N639 | N194;
  assign N639 = in_sig[28] & N373;
  assign N269 = N640 | N193;
  assign N640 = in_sig[27] & N373;
  assign N270 = N641 | N192;
  assign N641 = in_sig[26] & N373;
  assign N271 = N642 | N191;
  assign N642 = in_sig[25] & N373;
  assign N272 = N643 | N190;
  assign N643 = in_sig[24] & N373;
  assign N273 = N644 | N189;
  assign N644 = in_sig[23] & N373;
  assign N274 = N645 | N188;
  assign N645 = in_sig[22] & N373;
  assign N275 = N646 | N187;
  assign N646 = in_sig[21] & N373;
  assign N276 = N647 | N186;
  assign N647 = in_sig[20] & N373;
  assign N277 = N648 | N185;
  assign N648 = in_sig[19] & N373;
  assign N278 = N649 | N184;
  assign N649 = in_sig[18] & N373;
  assign N279 = N650 | N183;
  assign N650 = in_sig[17] & N373;
  assign N280 = N651 | N182;
  assign N651 = in_sig[16] & N373;
  assign N281 = N652 | N181;
  assign N652 = in_sig[15] & N373;
  assign N282 = N653 | N180;
  assign N653 = in_sig[14] & N373;
  assign N283 = N654 | N179;
  assign N654 = in_sig[13] & N373;
  assign N284 = N655 | N178;
  assign N655 = in_sig[12] & N373;
  assign N285 = N656 | N177;
  assign N656 = in_sig[11] & N373;
  assign common_inexact = 1'b0 | \genblk2.anyRound ;
  assign notNaN_isSpecialInfOut = exceptionFlags_3_ | in_isInf;
  assign commonCase = N659 & N660;
  assign N659 = N657 & N658;
  assign N657 = ~isNaNOut;
  assign N658 = ~notNaN_isSpecialInfOut;
  assign N660 = ~in_isZero;
  assign exceptionFlags[2] = commonCase & 1'b0;
  assign exceptionFlags[1] = commonCase & 1'b0;
  assign exceptionFlags[0] = exceptionFlags[2] | N661;
  assign N661 = commonCase & common_inexact;
  assign overflow_roundMagUp = N662 | roundMagUp;
  assign N662 = N349 | N346;
  assign pegMinNonzeroMagOut = N663 & N664;
  assign N663 = commonCase & 1'b0;
  assign N664 = roundMagUp | N353;
  assign pegMaxFiniteMagOut = exceptionFlags[2] & N665;
  assign N665 = ~overflow_roundMagUp;
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | N666;
  assign N666 = exceptionFlags[2] & overflow_roundMagUp;
  assign N286 = in_isZero | 1'b0;
  assign out[63] = N672 | isNaNOut;
  assign N672 = N671 | notNaN_isInfOut;
  assign N671 = N670 | pegMaxFiniteMagOut;
  assign N670 = N668 & N669;
  assign N668 = \genblk2.sRoundedExp [11] & N667;
  assign N667 = ~N286;
  assign N669 = ~pegMinNonzeroMagOut;
  assign out[62] = N677 | isNaNOut;
  assign N677 = N676 | notNaN_isInfOut;
  assign N676 = N674 & N675;
  assign N674 = N673 & N669;
  assign N673 = \genblk2.sRoundedExp [10] & N667;
  assign N675 = ~pegMaxFiniteMagOut;
  assign out[61] = N682 | isNaNOut;
  assign N682 = N681 | pegMaxFiniteMagOut;
  assign N681 = N680 | pegMinNonzeroMagOut;
  assign N680 = N678 & N679;
  assign N678 = \genblk2.sRoundedExp [9] & N667;
  assign N679 = ~notNaN_isInfOut;
  assign out[60] = N683 | pegMaxFiniteMagOut;
  assign N683 = \genblk2.sRoundedExp [8] | pegMinNonzeroMagOut;
  assign out[59] = N684 | pegMaxFiniteMagOut;
  assign N684 = \genblk2.sRoundedExp [7] | pegMinNonzeroMagOut;
  assign out[58] = N685 | pegMaxFiniteMagOut;
  assign N685 = \genblk2.sRoundedExp [6] | pegMinNonzeroMagOut;
  assign out[57] = N686 | pegMaxFiniteMagOut;
  assign N686 = \genblk2.sRoundedExp [5] & N669;
  assign out[56] = N687 | pegMaxFiniteMagOut;
  assign N687 = \genblk2.sRoundedExp [4] & N669;
  assign out[55] = N688 | pegMaxFiniteMagOut;
  assign N688 = \genblk2.sRoundedExp [3] | pegMinNonzeroMagOut;
  assign out[54] = N689 | pegMaxFiniteMagOut;
  assign N689 = \genblk2.sRoundedExp [2] | pegMinNonzeroMagOut;
  assign out[53] = N690 | pegMaxFiniteMagOut;
  assign N690 = \genblk2.sRoundedExp [1] | pegMinNonzeroMagOut;
  assign out[52] = N691 | pegMaxFiniteMagOut;
  assign N691 = \genblk2.sRoundedExp [0] & N669;
  assign N287 = N660 & N373;
  assign N288 = ~N287;
  assign N290 = N692 & N373;
  assign N692 = N657 & N660;
  assign N291 = ~N290;
  assign out[51] = N693 | pegMaxFiniteMagOut;
  assign N693 = isNaNOut | N289;
  assign out[50] = N342 | pegMaxFiniteMagOut;
  assign out[49] = N341 | pegMaxFiniteMagOut;
  assign out[48] = N340 | pegMaxFiniteMagOut;
  assign out[47] = N339 | pegMaxFiniteMagOut;
  assign out[46] = N338 | pegMaxFiniteMagOut;
  assign out[45] = N337 | pegMaxFiniteMagOut;
  assign out[44] = N336 | pegMaxFiniteMagOut;
  assign out[43] = N335 | pegMaxFiniteMagOut;
  assign out[42] = N334 | pegMaxFiniteMagOut;
  assign out[41] = N333 | pegMaxFiniteMagOut;
  assign out[40] = N332 | pegMaxFiniteMagOut;
  assign out[39] = N331 | pegMaxFiniteMagOut;
  assign out[38] = N330 | pegMaxFiniteMagOut;
  assign out[37] = N329 | pegMaxFiniteMagOut;
  assign out[36] = N328 | pegMaxFiniteMagOut;
  assign out[35] = N327 | pegMaxFiniteMagOut;
  assign out[34] = N326 | pegMaxFiniteMagOut;
  assign out[33] = N325 | pegMaxFiniteMagOut;
  assign out[32] = N324 | pegMaxFiniteMagOut;
  assign out[31] = N323 | pegMaxFiniteMagOut;
  assign out[30] = N322 | pegMaxFiniteMagOut;
  assign out[29] = N321 | pegMaxFiniteMagOut;
  assign out[28] = N320 | pegMaxFiniteMagOut;
  assign out[27] = N319 | pegMaxFiniteMagOut;
  assign out[26] = N318 | pegMaxFiniteMagOut;
  assign out[25] = N317 | pegMaxFiniteMagOut;
  assign out[24] = N316 | pegMaxFiniteMagOut;
  assign out[23] = N315 | pegMaxFiniteMagOut;
  assign out[22] = N314 | pegMaxFiniteMagOut;
  assign out[21] = N313 | pegMaxFiniteMagOut;
  assign out[20] = N312 | pegMaxFiniteMagOut;
  assign out[19] = N311 | pegMaxFiniteMagOut;
  assign out[18] = N310 | pegMaxFiniteMagOut;
  assign out[17] = N309 | pegMaxFiniteMagOut;
  assign out[16] = N308 | pegMaxFiniteMagOut;
  assign out[15] = N307 | pegMaxFiniteMagOut;
  assign out[14] = N306 | pegMaxFiniteMagOut;
  assign out[13] = N305 | pegMaxFiniteMagOut;
  assign out[12] = N304 | pegMaxFiniteMagOut;
  assign out[11] = N303 | pegMaxFiniteMagOut;
  assign out[10] = N302 | pegMaxFiniteMagOut;
  assign out[9] = N301 | pegMaxFiniteMagOut;
  assign out[8] = N300 | pegMaxFiniteMagOut;
  assign out[7] = N299 | pegMaxFiniteMagOut;
  assign out[6] = N298 | pegMaxFiniteMagOut;
  assign out[5] = N297 | pegMaxFiniteMagOut;
  assign out[4] = N296 | pegMaxFiniteMagOut;
  assign out[3] = N295 | pegMaxFiniteMagOut;
  assign out[2] = N294 | pegMaxFiniteMagOut;
  assign out[1] = N293 | pegMaxFiniteMagOut;
  assign out[0] = N292 | pegMaxFiniteMagOut;

endmodule



module iNToRecFN_intWidth64_expWidth11_sigWidth53
(
  control,
  signedIn,
  in,
  roundingMode,
  out,
  exceptionFlags
);

  input [0:0] control;
  input [63:0] in;
  input [2:0] roundingMode;
  output [64:0] out;
  output [4:0] exceptionFlags;
  input signedIn;
  wire [64:0] out,sig;
  wire [4:0] exceptionFlags;
  wire isZero,sign;
  wire [8:0] sExp;

  iNToRawFN_intWidth64
  iNToRawFN
  (
    .signedIn(signedIn),
    .in(in),
    .isZero(isZero),
    .sign(sign),
    .sExp(sExp),
    .sig(sig)
  );


  roundAnyRawFNToRecFN_inExpWidth7_inSigWidth64_outExpWidth11_outSigWidth53_options5
  roundRawToOut
  (
    .control(control[0]),
    .invalidExc(1'b0),
    .infiniteExc(1'b0),
    .in_isNaN(1'b0),
    .in_isInf(1'b0),
    .in_isZero(isZero),
    .in_sign(sign),
    .in_sExp(sExp),
    .in_sig(sig),
    .roundingMode(roundingMode),
    .out(out),
    .exceptionFlags(exceptionFlags)
  );


endmodule



module iNFromException_width64
(
  signedOut,
  isNaN,
  sign,
  out
);

  output [63:0] out;
  input signedOut;
  input isNaN;
  input sign;
  wire [63:0] out;
  wire out_62_,N0;
  assign out[0] = out_62_;
  assign out[1] = out_62_;
  assign out[2] = out_62_;
  assign out[3] = out_62_;
  assign out[4] = out_62_;
  assign out[5] = out_62_;
  assign out[6] = out_62_;
  assign out[7] = out_62_;
  assign out[8] = out_62_;
  assign out[9] = out_62_;
  assign out[10] = out_62_;
  assign out[11] = out_62_;
  assign out[12] = out_62_;
  assign out[13] = out_62_;
  assign out[14] = out_62_;
  assign out[15] = out_62_;
  assign out[16] = out_62_;
  assign out[17] = out_62_;
  assign out[18] = out_62_;
  assign out[19] = out_62_;
  assign out[20] = out_62_;
  assign out[21] = out_62_;
  assign out[22] = out_62_;
  assign out[23] = out_62_;
  assign out[24] = out_62_;
  assign out[25] = out_62_;
  assign out[26] = out_62_;
  assign out[27] = out_62_;
  assign out[28] = out_62_;
  assign out[29] = out_62_;
  assign out[30] = out_62_;
  assign out[31] = out_62_;
  assign out[32] = out_62_;
  assign out[33] = out_62_;
  assign out[34] = out_62_;
  assign out[35] = out_62_;
  assign out[36] = out_62_;
  assign out[37] = out_62_;
  assign out[38] = out_62_;
  assign out[39] = out_62_;
  assign out[40] = out_62_;
  assign out[41] = out_62_;
  assign out[42] = out_62_;
  assign out[43] = out_62_;
  assign out[44] = out_62_;
  assign out[45] = out_62_;
  assign out[46] = out_62_;
  assign out[47] = out_62_;
  assign out[48] = out_62_;
  assign out[49] = out_62_;
  assign out[50] = out_62_;
  assign out[51] = out_62_;
  assign out[52] = out_62_;
  assign out[53] = out_62_;
  assign out[54] = out_62_;
  assign out[55] = out_62_;
  assign out[56] = out_62_;
  assign out[57] = out_62_;
  assign out[58] = out_62_;
  assign out[59] = out_62_;
  assign out[60] = out_62_;
  assign out[61] = out_62_;
  assign out[62] = out_62_;
  assign out_62_ = isNaN | N0;
  assign N0 = ~sign;
  assign out[63] = signedOut ^ out_62_;

endmodule



module recFNToIN_expWidth11_sigWidth53_intWidth64
(
  control,
  in,
  roundingMode,
  signedOut,
  out,
  intExceptionFlags
);

  input [0:0] control;
  input [64:0] in;
  input [2:0] roundingMode;
  output [63:0] out;
  output [2:0] intExceptionFlags;
  input signedOut;
  wire [63:0] out,complUnroundedInt,roundedInt,excOut;
  wire [2:0] intExceptionFlags;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,isNaN,isInf,isZero,sign,magJustBelowOne,
  N12,N13,N14,N15,N16,N17,N18,common_inexact,N19,roundIncr_near_even,
  roundIncr_near_maxMag,roundIncr,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,
  N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,
  N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,
  N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,
  N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,
  N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,
  N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,
  N144,N145,N146,N147,N148,N149,N150,N151,N152,roundCarryBut2,N153,N154,N155,N156,
  N157,N158,N159,N160,N161,N162,N163,N164,common_overflow,N165,N166,N167,N168,N169,
  N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,
  N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,
  N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,
  N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,
  N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,
  N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,
  N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,
  N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,
  N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,
  N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,
  N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,
  N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,
  N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,
  N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,
  N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,
  N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425;
  wire [12:0] sExp;
  wire [53:0] sig;
  wire [115:0] shiftedSig;
  wire [0:0] alignedSig;

  recFNToRawFN_expWidth11_sigWidth53
  recFNToRawFN
  (
    .in(in),
    .isNaN(isNaN),
    .isInf(isInf),
    .isZero(isZero),
    .sign(sign),
    .sExp(sExp),
    .sig(sig)
  );


  iNFromException_width64
  iNFromException
  (
    .signedOut(signedOut),
    .isNaN(isNaN),
    .sign(sign),
    .out(excOut)
  );

  assign N168 = ~sExp[5];
  assign N169 = ~sExp[4];
  assign N170 = ~sExp[3];
  assign N171 = ~sExp[2];
  assign N172 = ~sExp[1];
  assign N173 = ~sExp[0];
  assign N174 = sExp[9] | sExp[10];
  assign N175 = sExp[8] | N174;
  assign N176 = sExp[7] | N175;
  assign N177 = sExp[6] | N176;
  assign N178 = N168 | N177;
  assign N179 = N169 | N178;
  assign N180 = N170 | N179;
  assign N181 = N171 | N180;
  assign N182 = N172 | N181;
  assign N183 = N173 | N182;
  assign N184 = ~N183;
  assign N185 = sExp[9] | sExp[10];
  assign N186 = sExp[8] | N185;
  assign N187 = sExp[7] | N186;
  assign N188 = sExp[6] | N187;
  assign N189 = N168 | N188;
  assign N190 = N169 | N189;
  assign N191 = N170 | N190;
  assign N192 = N171 | N191;
  assign N193 = N172 | N192;
  assign N194 = sExp[0] | N193;
  assign N195 = ~N194;
  assign N196 = roundingMode[1] | roundingMode[2];
  assign N197 = roundingMode[0] | N196;
  assign N198 = ~N197;
  assign N199 = ~roundingMode[2];
  assign N200 = roundingMode[1] | N199;
  assign N201 = roundingMode[0] | N200;
  assign N202 = ~N201;
  assign N203 = ~roundingMode[1];
  assign N204 = N203 | roundingMode[2];
  assign N205 = roundingMode[0] | N204;
  assign N206 = ~N205;
  assign N207 = N203 | N199;
  assign N208 = roundingMode[0] | N207;
  assign N209 = ~N208;
  assign N210 = ~roundingMode[0];
  assign N211 = N210 | N204;
  assign N212 = ~N211;
  assign shiftedSig = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sExp[11:11], sig[51:0] } << { N17, N16, N15, N14, N13, N12 };
  assign { N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88 } = complUnroundedInt + 1'b1;
  assign { N17, N16, N15, N14, N13, N12 } = (N0)? sExp[5:0] : 
                                            (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = sExp[11];
  assign N1 = N213;
  assign common_inexact = (N0)? N18 : 
                          (N1)? N19 : 1'b0;
  assign complUnroundedInt = (N2)? { N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85 } : 
                             (N3)? shiftedSig[115:52] : 1'b0;
  assign N2 = N21;
  assign N3 = N20;
  assign { roundedInt[63:1], N152 } = (N4)? { N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88 } : 
                                      (N87)? complUnroundedInt : 1'b0;
  assign N4 = N86;
  assign N159 = (N5)? N157 : 
                (N6)? N158 : 1'b0;
  assign N5 = N156;
  assign N6 = N155;
  assign N161 = (N7)? N159 : 
                (N8)? N160 : 1'b0;
  assign N7 = N154;
  assign N8 = N153;
  assign N164 = (N9)? 1'b1 : 
                (N10)? N161 : 1'b0;
  assign N9 = N162;
  assign N10 = N163;
  assign common_overflow = (N0)? N164 : 
                           (N1)? N165 : 1'b0;
  assign out = (N11)? excOut : 
               (N167)? roundedInt : 1'b0;
  assign N11 = N166;
  assign magJustBelowOne = N213 & N223;
  assign N213 = ~sExp[11];
  assign N223 = N222 & sExp[0];
  assign N222 = N221 & sExp[1];
  assign N221 = N220 & sExp[2];
  assign N220 = N219 & sExp[3];
  assign N219 = N218 & sExp[4];
  assign N218 = N217 & sExp[5];
  assign N217 = N216 & sExp[6];
  assign N216 = N215 & sExp[7];
  assign N215 = N214 & sExp[8];
  assign N214 = sExp[10] & sExp[9];
  assign alignedSig[0] = N272 | shiftedSig[0];
  assign N272 = N271 | shiftedSig[1];
  assign N271 = N270 | shiftedSig[2];
  assign N270 = N269 | shiftedSig[3];
  assign N269 = N268 | shiftedSig[4];
  assign N268 = N267 | shiftedSig[5];
  assign N267 = N266 | shiftedSig[6];
  assign N266 = N265 | shiftedSig[7];
  assign N265 = N264 | shiftedSig[8];
  assign N264 = N263 | shiftedSig[9];
  assign N263 = N262 | shiftedSig[10];
  assign N262 = N261 | shiftedSig[11];
  assign N261 = N260 | shiftedSig[12];
  assign N260 = N259 | shiftedSig[13];
  assign N259 = N258 | shiftedSig[14];
  assign N258 = N257 | shiftedSig[15];
  assign N257 = N256 | shiftedSig[16];
  assign N256 = N255 | shiftedSig[17];
  assign N255 = N254 | shiftedSig[18];
  assign N254 = N253 | shiftedSig[19];
  assign N253 = N252 | shiftedSig[20];
  assign N252 = N251 | shiftedSig[21];
  assign N251 = N250 | shiftedSig[22];
  assign N250 = N249 | shiftedSig[23];
  assign N249 = N248 | shiftedSig[24];
  assign N248 = N247 | shiftedSig[25];
  assign N247 = N246 | shiftedSig[26];
  assign N246 = N245 | shiftedSig[27];
  assign N245 = N244 | shiftedSig[28];
  assign N244 = N243 | shiftedSig[29];
  assign N243 = N242 | shiftedSig[30];
  assign N242 = N241 | shiftedSig[31];
  assign N241 = N240 | shiftedSig[32];
  assign N240 = N239 | shiftedSig[33];
  assign N239 = N238 | shiftedSig[34];
  assign N238 = N237 | shiftedSig[35];
  assign N237 = N236 | shiftedSig[36];
  assign N236 = N235 | shiftedSig[37];
  assign N235 = N234 | shiftedSig[38];
  assign N234 = N233 | shiftedSig[39];
  assign N233 = N232 | shiftedSig[40];
  assign N232 = N231 | shiftedSig[41];
  assign N231 = N230 | shiftedSig[42];
  assign N230 = N229 | shiftedSig[43];
  assign N229 = N228 | shiftedSig[44];
  assign N228 = N227 | shiftedSig[45];
  assign N227 = N226 | shiftedSig[46];
  assign N226 = N225 | shiftedSig[47];
  assign N225 = N224 | shiftedSig[48];
  assign N224 = shiftedSig[50] | shiftedSig[49];
  assign N18 = shiftedSig[51] | alignedSig[0];
  assign N19 = ~isZero;
  assign roundIncr_near_even = N276 | N278;
  assign N276 = sExp[11] & N275;
  assign N275 = N273 | N274;
  assign N273 = shiftedSig[52] & shiftedSig[51];
  assign N274 = shiftedSig[51] & alignedSig[0];
  assign N278 = magJustBelowOne & N277;
  assign N277 = shiftedSig[51] | alignedSig[0];
  assign roundIncr_near_maxMag = N279 | magJustBelowOne;
  assign N279 = sExp[11] & shiftedSig[51];
  assign roundIncr = N286 | N289;
  assign N286 = N282 | N285;
  assign N282 = N280 | N281;
  assign N280 = N198 & roundIncr_near_even;
  assign N281 = N202 & roundIncr_near_maxMag;
  assign N285 = N283 & N284;
  assign N283 = N206 | N209;
  assign N284 = sign & common_inexact;
  assign N289 = N212 & N288;
  assign N288 = N287 & common_inexact;
  assign N287 = ~sign;
  assign N20 = ~sign;
  assign N21 = sign;
  assign N22 = ~shiftedSig[115];
  assign N23 = ~shiftedSig[114];
  assign N24 = ~shiftedSig[113];
  assign N25 = ~shiftedSig[112];
  assign N26 = ~shiftedSig[111];
  assign N27 = ~shiftedSig[110];
  assign N28 = ~shiftedSig[109];
  assign N29 = ~shiftedSig[108];
  assign N30 = ~shiftedSig[107];
  assign N31 = ~shiftedSig[106];
  assign N32 = ~shiftedSig[105];
  assign N33 = ~shiftedSig[104];
  assign N34 = ~shiftedSig[103];
  assign N35 = ~shiftedSig[102];
  assign N36 = ~shiftedSig[101];
  assign N37 = ~shiftedSig[100];
  assign N38 = ~shiftedSig[99];
  assign N39 = ~shiftedSig[98];
  assign N40 = ~shiftedSig[97];
  assign N41 = ~shiftedSig[96];
  assign N42 = ~shiftedSig[95];
  assign N43 = ~shiftedSig[94];
  assign N44 = ~shiftedSig[93];
  assign N45 = ~shiftedSig[92];
  assign N46 = ~shiftedSig[91];
  assign N47 = ~shiftedSig[90];
  assign N48 = ~shiftedSig[89];
  assign N49 = ~shiftedSig[88];
  assign N50 = ~shiftedSig[87];
  assign N51 = ~shiftedSig[86];
  assign N52 = ~shiftedSig[85];
  assign N53 = ~shiftedSig[84];
  assign N54 = ~shiftedSig[83];
  assign N55 = ~shiftedSig[82];
  assign N56 = ~shiftedSig[81];
  assign N57 = ~shiftedSig[80];
  assign N58 = ~shiftedSig[79];
  assign N59 = ~shiftedSig[78];
  assign N60 = ~shiftedSig[77];
  assign N61 = ~shiftedSig[76];
  assign N62 = ~shiftedSig[75];
  assign N63 = ~shiftedSig[74];
  assign N64 = ~shiftedSig[73];
  assign N65 = ~shiftedSig[72];
  assign N66 = ~shiftedSig[71];
  assign N67 = ~shiftedSig[70];
  assign N68 = ~shiftedSig[69];
  assign N69 = ~shiftedSig[68];
  assign N70 = ~shiftedSig[67];
  assign N71 = ~shiftedSig[66];
  assign N72 = ~shiftedSig[65];
  assign N73 = ~shiftedSig[64];
  assign N74 = ~shiftedSig[63];
  assign N75 = ~shiftedSig[62];
  assign N76 = ~shiftedSig[61];
  assign N77 = ~shiftedSig[60];
  assign N78 = ~shiftedSig[59];
  assign N79 = ~shiftedSig[58];
  assign N80 = ~shiftedSig[57];
  assign N81 = ~shiftedSig[56];
  assign N82 = ~shiftedSig[55];
  assign N83 = ~shiftedSig[54];
  assign N84 = ~shiftedSig[53];
  assign N85 = ~shiftedSig[52];
  assign N86 = roundIncr ^ sign;
  assign N87 = ~N86;
  assign roundedInt[0] = N152 | N290;
  assign N290 = N209 & common_inexact;
  assign roundCarryBut2 = N351 & roundIncr;
  assign N351 = N350 & shiftedSig[52];
  assign N350 = N349 & shiftedSig[53];
  assign N349 = N348 & shiftedSig[54];
  assign N348 = N347 & shiftedSig[55];
  assign N347 = N346 & shiftedSig[56];
  assign N346 = N345 & shiftedSig[57];
  assign N345 = N344 & shiftedSig[58];
  assign N344 = N343 & shiftedSig[59];
  assign N343 = N342 & shiftedSig[60];
  assign N342 = N341 & shiftedSig[61];
  assign N341 = N340 & shiftedSig[62];
  assign N340 = N339 & shiftedSig[63];
  assign N339 = N338 & shiftedSig[64];
  assign N338 = N337 & shiftedSig[65];
  assign N337 = N336 & shiftedSig[66];
  assign N336 = N335 & shiftedSig[67];
  assign N335 = N334 & shiftedSig[68];
  assign N334 = N333 & shiftedSig[69];
  assign N333 = N332 & shiftedSig[70];
  assign N332 = N331 & shiftedSig[71];
  assign N331 = N330 & shiftedSig[72];
  assign N330 = N329 & shiftedSig[73];
  assign N329 = N328 & shiftedSig[74];
  assign N328 = N327 & shiftedSig[75];
  assign N327 = N326 & shiftedSig[76];
  assign N326 = N325 & shiftedSig[77];
  assign N325 = N324 & shiftedSig[78];
  assign N324 = N323 & shiftedSig[79];
  assign N323 = N322 & shiftedSig[80];
  assign N322 = N321 & shiftedSig[81];
  assign N321 = N320 & shiftedSig[82];
  assign N320 = N319 & shiftedSig[83];
  assign N319 = N318 & shiftedSig[84];
  assign N318 = N317 & shiftedSig[85];
  assign N317 = N316 & shiftedSig[86];
  assign N316 = N315 & shiftedSig[87];
  assign N315 = N314 & shiftedSig[88];
  assign N314 = N313 & shiftedSig[89];
  assign N313 = N312 & shiftedSig[90];
  assign N312 = N311 & shiftedSig[91];
  assign N311 = N310 & shiftedSig[92];
  assign N310 = N309 & shiftedSig[93];
  assign N309 = N308 & shiftedSig[94];
  assign N308 = N307 & shiftedSig[95];
  assign N307 = N306 & shiftedSig[96];
  assign N306 = N305 & shiftedSig[97];
  assign N305 = N304 & shiftedSig[98];
  assign N304 = N303 & shiftedSig[99];
  assign N303 = N302 & shiftedSig[100];
  assign N302 = N301 & shiftedSig[101];
  assign N301 = N300 & shiftedSig[102];
  assign N300 = N299 & shiftedSig[103];
  assign N299 = N298 & shiftedSig[104];
  assign N298 = N297 & shiftedSig[105];
  assign N297 = N296 & shiftedSig[106];
  assign N296 = N295 & shiftedSig[107];
  assign N295 = N294 & shiftedSig[108];
  assign N294 = N293 & shiftedSig[109];
  assign N293 = N292 & shiftedSig[110];
  assign N292 = N291 & shiftedSig[111];
  assign N291 = shiftedSig[113] & shiftedSig[112];
  assign N153 = ~signedOut;
  assign N154 = signedOut;
  assign N155 = ~sign;
  assign N156 = sign;
  assign N157 = N184 & N414;
  assign N414 = N413 | roundIncr;
  assign N413 = N412 | shiftedSig[52];
  assign N412 = N411 | shiftedSig[53];
  assign N411 = N410 | shiftedSig[54];
  assign N410 = N409 | shiftedSig[55];
  assign N409 = N408 | shiftedSig[56];
  assign N408 = N407 | shiftedSig[57];
  assign N407 = N406 | shiftedSig[58];
  assign N406 = N405 | shiftedSig[59];
  assign N405 = N404 | shiftedSig[60];
  assign N404 = N403 | shiftedSig[61];
  assign N403 = N402 | shiftedSig[62];
  assign N402 = N401 | shiftedSig[63];
  assign N401 = N400 | shiftedSig[64];
  assign N400 = N399 | shiftedSig[65];
  assign N399 = N398 | shiftedSig[66];
  assign N398 = N397 | shiftedSig[67];
  assign N397 = N396 | shiftedSig[68];
  assign N396 = N395 | shiftedSig[69];
  assign N395 = N394 | shiftedSig[70];
  assign N394 = N393 | shiftedSig[71];
  assign N393 = N392 | shiftedSig[72];
  assign N392 = N391 | shiftedSig[73];
  assign N391 = N390 | shiftedSig[74];
  assign N390 = N389 | shiftedSig[75];
  assign N389 = N388 | shiftedSig[76];
  assign N388 = N387 | shiftedSig[77];
  assign N387 = N386 | shiftedSig[78];
  assign N386 = N385 | shiftedSig[79];
  assign N385 = N384 | shiftedSig[80];
  assign N384 = N383 | shiftedSig[81];
  assign N383 = N382 | shiftedSig[82];
  assign N382 = N381 | shiftedSig[83];
  assign N381 = N380 | shiftedSig[84];
  assign N380 = N379 | shiftedSig[85];
  assign N379 = N378 | shiftedSig[86];
  assign N378 = N377 | shiftedSig[87];
  assign N377 = N376 | shiftedSig[88];
  assign N376 = N375 | shiftedSig[89];
  assign N375 = N374 | shiftedSig[90];
  assign N374 = N373 | shiftedSig[91];
  assign N373 = N372 | shiftedSig[92];
  assign N372 = N371 | shiftedSig[93];
  assign N371 = N370 | shiftedSig[94];
  assign N370 = N369 | shiftedSig[95];
  assign N369 = N368 | shiftedSig[96];
  assign N368 = N367 | shiftedSig[97];
  assign N367 = N366 | shiftedSig[98];
  assign N366 = N365 | shiftedSig[99];
  assign N365 = N364 | shiftedSig[100];
  assign N364 = N363 | shiftedSig[101];
  assign N363 = N362 | shiftedSig[102];
  assign N362 = N361 | shiftedSig[103];
  assign N361 = N360 | shiftedSig[104];
  assign N360 = N359 | shiftedSig[105];
  assign N359 = N358 | shiftedSig[106];
  assign N358 = N357 | shiftedSig[107];
  assign N357 = N356 | shiftedSig[108];
  assign N356 = N355 | shiftedSig[109];
  assign N355 = N354 | shiftedSig[110];
  assign N354 = N353 | shiftedSig[111];
  assign N353 = N352 | shiftedSig[112];
  assign N352 = shiftedSig[114] | shiftedSig[113];
  assign N158 = N184 | N415;
  assign N415 = N195 & roundCarryBut2;
  assign N160 = sign | N417;
  assign N417 = N416 & roundCarryBut2;
  assign N416 = N184 & shiftedSig[114];
  assign N162 = N420 | sExp[6];
  assign N420 = N419 | sExp[7];
  assign N419 = N418 | sExp[8];
  assign N418 = sExp[10] | sExp[9];
  assign N163 = ~N162;
  assign N165 = N422 & roundIncr;
  assign N422 = N421 & sign;
  assign N421 = ~signedOut;
  assign intExceptionFlags[2] = isNaN | isInf;
  assign intExceptionFlags[1] = N423 & common_overflow;
  assign N423 = ~intExceptionFlags[2];
  assign intExceptionFlags[0] = N425 & common_inexact;
  assign N425 = N423 & N424;
  assign N424 = ~common_overflow;
  assign N166 = intExceptionFlags[2] | common_overflow;
  assign N167 = ~N166;

endmodule



module iNFromException_width32
(
  signedOut,
  isNaN,
  sign,
  out
);

  output [31:0] out;
  input signedOut;
  input isNaN;
  input sign;
  wire [31:0] out;
  wire out_30_,N0;
  assign out[0] = out_30_;
  assign out[1] = out_30_;
  assign out[2] = out_30_;
  assign out[3] = out_30_;
  assign out[4] = out_30_;
  assign out[5] = out_30_;
  assign out[6] = out_30_;
  assign out[7] = out_30_;
  assign out[8] = out_30_;
  assign out[9] = out_30_;
  assign out[10] = out_30_;
  assign out[11] = out_30_;
  assign out[12] = out_30_;
  assign out[13] = out_30_;
  assign out[14] = out_30_;
  assign out[15] = out_30_;
  assign out[16] = out_30_;
  assign out[17] = out_30_;
  assign out[18] = out_30_;
  assign out[19] = out_30_;
  assign out[20] = out_30_;
  assign out[21] = out_30_;
  assign out[22] = out_30_;
  assign out[23] = out_30_;
  assign out[24] = out_30_;
  assign out[25] = out_30_;
  assign out[26] = out_30_;
  assign out[27] = out_30_;
  assign out[28] = out_30_;
  assign out[29] = out_30_;
  assign out[30] = out_30_;
  assign out_30_ = isNaN | N0;
  assign N0 = ~sign;
  assign out[31] = signedOut ^ out_30_;

endmodule



module recFNToIN_expWidth11_sigWidth53_intWidth32
(
  control,
  in,
  roundingMode,
  signedOut,
  out,
  intExceptionFlags
);

  input [0:0] control;
  input [64:0] in;
  input [2:0] roundingMode;
  output [31:0] out;
  output [2:0] intExceptionFlags;
  input signedOut;
  wire [31:0] out,complUnroundedInt,roundedInt,excOut;
  wire [2:0] intExceptionFlags;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,isNaN,isInf,isZero,sign,magJustBelowOne,
  N12,N13,N14,N15,N16,N17,common_inexact,N18,roundIncr_near_even,
  roundIncr_near_maxMag,roundIncr,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,
  N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,
  N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,
  N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,roundCarryBut2,N88,N89,N90,N91,
  N92,N93,N94,N95,N96,N97,N98,N99,common_overflow,N100,N101,N102,N103,N104,N105,
  N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,
  N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,
  N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,
  N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,
  N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,
  N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,
  N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,
  N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,
  N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,
  N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,
  N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,
  N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296;
  wire [12:0] sExp;
  wire [53:0] sig;
  wire [83:0] shiftedSig;
  wire [0:0] alignedSig;

  recFNToRawFN_expWidth11_sigWidth53
  recFNToRawFN
  (
    .in(in),
    .isNaN(isNaN),
    .isInf(isInf),
    .isZero(isZero),
    .sign(sign),
    .sExp(sExp),
    .sig(sig)
  );


  iNFromException_width32
  iNFromException
  (
    .signedOut(signedOut),
    .isNaN(isNaN),
    .sign(sign),
    .out(excOut)
  );

  assign N103 = ~sExp[4];
  assign N104 = ~sExp[3];
  assign N105 = ~sExp[2];
  assign N106 = ~sExp[1];
  assign N107 = ~sExp[0];
  assign N108 = sExp[9] | sExp[10];
  assign N109 = sExp[8] | N108;
  assign N110 = sExp[7] | N109;
  assign N111 = sExp[6] | N110;
  assign N112 = sExp[5] | N111;
  assign N113 = N103 | N112;
  assign N114 = N104 | N113;
  assign N115 = N105 | N114;
  assign N116 = N106 | N115;
  assign N117 = N107 | N116;
  assign N118 = ~N117;
  assign N119 = sExp[9] | sExp[10];
  assign N120 = sExp[8] | N119;
  assign N121 = sExp[7] | N120;
  assign N122 = sExp[6] | N121;
  assign N123 = sExp[5] | N122;
  assign N124 = N103 | N123;
  assign N125 = N104 | N124;
  assign N126 = N105 | N125;
  assign N127 = N106 | N126;
  assign N128 = sExp[0] | N127;
  assign N129 = ~N128;
  assign N130 = roundingMode[1] | roundingMode[2];
  assign N131 = roundingMode[0] | N130;
  assign N132 = ~N131;
  assign N133 = ~roundingMode[2];
  assign N134 = roundingMode[1] | N133;
  assign N135 = roundingMode[0] | N134;
  assign N136 = ~N135;
  assign N137 = ~roundingMode[1];
  assign N138 = N137 | roundingMode[2];
  assign N139 = roundingMode[0] | N138;
  assign N140 = ~N139;
  assign N141 = N137 | N133;
  assign N142 = roundingMode[0] | N141;
  assign N143 = ~N142;
  assign N144 = ~roundingMode[0];
  assign N145 = N144 | N138;
  assign N146 = ~N145;
  assign shiftedSig = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sExp[11:11], sig[51:0] } << { N16, N15, N14, N13, N12 };
  assign { N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55 } = complUnroundedInt + 1'b1;
  assign { N16, N15, N14, N13, N12 } = (N0)? sExp[4:0] : 
                                       (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = sExp[11];
  assign N1 = N147;
  assign common_inexact = (N0)? N17 : 
                          (N1)? N18 : 1'b0;
  assign complUnroundedInt = (N2)? { N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52 } : 
                             (N3)? shiftedSig[83:52] : 1'b0;
  assign N2 = N20;
  assign N3 = N19;
  assign { roundedInt[31:1], N87 } = (N4)? { N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55 } : 
                                     (N54)? complUnroundedInt : 1'b0;
  assign N4 = N53;
  assign N94 = (N5)? N92 : 
               (N6)? N93 : 1'b0;
  assign N5 = N91;
  assign N6 = N90;
  assign N96 = (N7)? N94 : 
               (N8)? N95 : 1'b0;
  assign N7 = N89;
  assign N8 = N88;
  assign N99 = (N9)? 1'b1 : 
               (N10)? N96 : 1'b0;
  assign N9 = N97;
  assign N10 = N98;
  assign common_overflow = (N0)? N99 : 
                           (N1)? N100 : 1'b0;
  assign out = (N11)? excOut : 
               (N102)? roundedInt : 1'b0;
  assign N11 = N101;
  assign magJustBelowOne = N147 & N157;
  assign N147 = ~sExp[11];
  assign N157 = N156 & sExp[0];
  assign N156 = N155 & sExp[1];
  assign N155 = N154 & sExp[2];
  assign N154 = N153 & sExp[3];
  assign N153 = N152 & sExp[4];
  assign N152 = N151 & sExp[5];
  assign N151 = N150 & sExp[6];
  assign N150 = N149 & sExp[7];
  assign N149 = N148 & sExp[8];
  assign N148 = sExp[10] & sExp[9];
  assign alignedSig[0] = N206 | shiftedSig[0];
  assign N206 = N205 | shiftedSig[1];
  assign N205 = N204 | shiftedSig[2];
  assign N204 = N203 | shiftedSig[3];
  assign N203 = N202 | shiftedSig[4];
  assign N202 = N201 | shiftedSig[5];
  assign N201 = N200 | shiftedSig[6];
  assign N200 = N199 | shiftedSig[7];
  assign N199 = N198 | shiftedSig[8];
  assign N198 = N197 | shiftedSig[9];
  assign N197 = N196 | shiftedSig[10];
  assign N196 = N195 | shiftedSig[11];
  assign N195 = N194 | shiftedSig[12];
  assign N194 = N193 | shiftedSig[13];
  assign N193 = N192 | shiftedSig[14];
  assign N192 = N191 | shiftedSig[15];
  assign N191 = N190 | shiftedSig[16];
  assign N190 = N189 | shiftedSig[17];
  assign N189 = N188 | shiftedSig[18];
  assign N188 = N187 | shiftedSig[19];
  assign N187 = N186 | shiftedSig[20];
  assign N186 = N185 | shiftedSig[21];
  assign N185 = N184 | shiftedSig[22];
  assign N184 = N183 | shiftedSig[23];
  assign N183 = N182 | shiftedSig[24];
  assign N182 = N181 | shiftedSig[25];
  assign N181 = N180 | shiftedSig[26];
  assign N180 = N179 | shiftedSig[27];
  assign N179 = N178 | shiftedSig[28];
  assign N178 = N177 | shiftedSig[29];
  assign N177 = N176 | shiftedSig[30];
  assign N176 = N175 | shiftedSig[31];
  assign N175 = N174 | shiftedSig[32];
  assign N174 = N173 | shiftedSig[33];
  assign N173 = N172 | shiftedSig[34];
  assign N172 = N171 | shiftedSig[35];
  assign N171 = N170 | shiftedSig[36];
  assign N170 = N169 | shiftedSig[37];
  assign N169 = N168 | shiftedSig[38];
  assign N168 = N167 | shiftedSig[39];
  assign N167 = N166 | shiftedSig[40];
  assign N166 = N165 | shiftedSig[41];
  assign N165 = N164 | shiftedSig[42];
  assign N164 = N163 | shiftedSig[43];
  assign N163 = N162 | shiftedSig[44];
  assign N162 = N161 | shiftedSig[45];
  assign N161 = N160 | shiftedSig[46];
  assign N160 = N159 | shiftedSig[47];
  assign N159 = N158 | shiftedSig[48];
  assign N158 = shiftedSig[50] | shiftedSig[49];
  assign N17 = shiftedSig[51] | alignedSig[0];
  assign N18 = ~isZero;
  assign roundIncr_near_even = N210 | N212;
  assign N210 = sExp[11] & N209;
  assign N209 = N207 | N208;
  assign N207 = shiftedSig[52] & shiftedSig[51];
  assign N208 = shiftedSig[51] & alignedSig[0];
  assign N212 = magJustBelowOne & N211;
  assign N211 = shiftedSig[51] | alignedSig[0];
  assign roundIncr_near_maxMag = N213 | magJustBelowOne;
  assign N213 = sExp[11] & shiftedSig[51];
  assign roundIncr = N220 | N223;
  assign N220 = N216 | N219;
  assign N216 = N214 | N215;
  assign N214 = N132 & roundIncr_near_even;
  assign N215 = N136 & roundIncr_near_maxMag;
  assign N219 = N217 & N218;
  assign N217 = N140 | N143;
  assign N218 = sign & common_inexact;
  assign N223 = N146 & N222;
  assign N222 = N221 & common_inexact;
  assign N221 = ~sign;
  assign N19 = ~sign;
  assign N20 = sign;
  assign N21 = ~shiftedSig[83];
  assign N22 = ~shiftedSig[82];
  assign N23 = ~shiftedSig[81];
  assign N24 = ~shiftedSig[80];
  assign N25 = ~shiftedSig[79];
  assign N26 = ~shiftedSig[78];
  assign N27 = ~shiftedSig[77];
  assign N28 = ~shiftedSig[76];
  assign N29 = ~shiftedSig[75];
  assign N30 = ~shiftedSig[74];
  assign N31 = ~shiftedSig[73];
  assign N32 = ~shiftedSig[72];
  assign N33 = ~shiftedSig[71];
  assign N34 = ~shiftedSig[70];
  assign N35 = ~shiftedSig[69];
  assign N36 = ~shiftedSig[68];
  assign N37 = ~shiftedSig[67];
  assign N38 = ~shiftedSig[66];
  assign N39 = ~shiftedSig[65];
  assign N40 = ~shiftedSig[64];
  assign N41 = ~shiftedSig[63];
  assign N42 = ~shiftedSig[62];
  assign N43 = ~shiftedSig[61];
  assign N44 = ~shiftedSig[60];
  assign N45 = ~shiftedSig[59];
  assign N46 = ~shiftedSig[58];
  assign N47 = ~shiftedSig[57];
  assign N48 = ~shiftedSig[56];
  assign N49 = ~shiftedSig[55];
  assign N50 = ~shiftedSig[54];
  assign N51 = ~shiftedSig[53];
  assign N52 = ~shiftedSig[52];
  assign N53 = roundIncr ^ sign;
  assign N54 = ~N53;
  assign roundedInt[0] = N87 | N224;
  assign N224 = N143 & common_inexact;
  assign roundCarryBut2 = N253 & roundIncr;
  assign N253 = N252 & shiftedSig[52];
  assign N252 = N251 & shiftedSig[53];
  assign N251 = N250 & shiftedSig[54];
  assign N250 = N249 & shiftedSig[55];
  assign N249 = N248 & shiftedSig[56];
  assign N248 = N247 & shiftedSig[57];
  assign N247 = N246 & shiftedSig[58];
  assign N246 = N245 & shiftedSig[59];
  assign N245 = N244 & shiftedSig[60];
  assign N244 = N243 & shiftedSig[61];
  assign N243 = N242 & shiftedSig[62];
  assign N242 = N241 & shiftedSig[63];
  assign N241 = N240 & shiftedSig[64];
  assign N240 = N239 & shiftedSig[65];
  assign N239 = N238 & shiftedSig[66];
  assign N238 = N237 & shiftedSig[67];
  assign N237 = N236 & shiftedSig[68];
  assign N236 = N235 & shiftedSig[69];
  assign N235 = N234 & shiftedSig[70];
  assign N234 = N233 & shiftedSig[71];
  assign N233 = N232 & shiftedSig[72];
  assign N232 = N231 & shiftedSig[73];
  assign N231 = N230 & shiftedSig[74];
  assign N230 = N229 & shiftedSig[75];
  assign N229 = N228 & shiftedSig[76];
  assign N228 = N227 & shiftedSig[77];
  assign N227 = N226 & shiftedSig[78];
  assign N226 = N225 & shiftedSig[79];
  assign N225 = shiftedSig[81] & shiftedSig[80];
  assign N88 = ~signedOut;
  assign N89 = signedOut;
  assign N90 = ~sign;
  assign N91 = sign;
  assign N92 = N118 & N284;
  assign N284 = N283 | roundIncr;
  assign N283 = N282 | shiftedSig[52];
  assign N282 = N281 | shiftedSig[53];
  assign N281 = N280 | shiftedSig[54];
  assign N280 = N279 | shiftedSig[55];
  assign N279 = N278 | shiftedSig[56];
  assign N278 = N277 | shiftedSig[57];
  assign N277 = N276 | shiftedSig[58];
  assign N276 = N275 | shiftedSig[59];
  assign N275 = N274 | shiftedSig[60];
  assign N274 = N273 | shiftedSig[61];
  assign N273 = N272 | shiftedSig[62];
  assign N272 = N271 | shiftedSig[63];
  assign N271 = N270 | shiftedSig[64];
  assign N270 = N269 | shiftedSig[65];
  assign N269 = N268 | shiftedSig[66];
  assign N268 = N267 | shiftedSig[67];
  assign N267 = N266 | shiftedSig[68];
  assign N266 = N265 | shiftedSig[69];
  assign N265 = N264 | shiftedSig[70];
  assign N264 = N263 | shiftedSig[71];
  assign N263 = N262 | shiftedSig[72];
  assign N262 = N261 | shiftedSig[73];
  assign N261 = N260 | shiftedSig[74];
  assign N260 = N259 | shiftedSig[75];
  assign N259 = N258 | shiftedSig[76];
  assign N258 = N257 | shiftedSig[77];
  assign N257 = N256 | shiftedSig[78];
  assign N256 = N255 | shiftedSig[79];
  assign N255 = N254 | shiftedSig[80];
  assign N254 = shiftedSig[82] | shiftedSig[81];
  assign N93 = N118 | N285;
  assign N285 = N129 & roundCarryBut2;
  assign N95 = sign | N287;
  assign N287 = N286 & roundCarryBut2;
  assign N286 = N118 & shiftedSig[82];
  assign N97 = N291 | sExp[5];
  assign N291 = N290 | sExp[6];
  assign N290 = N289 | sExp[7];
  assign N289 = N288 | sExp[8];
  assign N288 = sExp[10] | sExp[9];
  assign N98 = ~N97;
  assign N100 = N293 & roundIncr;
  assign N293 = N292 & sign;
  assign N292 = ~signedOut;
  assign intExceptionFlags[2] = isNaN | isInf;
  assign intExceptionFlags[1] = N294 & common_overflow;
  assign N294 = ~intExceptionFlags[2];
  assign intExceptionFlags[0] = N296 & common_inexact;
  assign N296 = N294 & N295;
  assign N295 = ~common_overflow;
  assign N101 = intExceptionFlags[2] | common_overflow;
  assign N102 = ~N101;

endmodule



module compareRecFN_expWidth11_sigWidth53
(
  a,
  b,
  signaling,
  lt,
  eq,
  gt,
  unordered,
  exceptionFlags
);

  input [64:0] a;
  input [64:0] b;
  output [4:0] exceptionFlags;
  input signaling;
  output lt;
  output eq;
  output gt;
  output unordered;
  wire [4:0] exceptionFlags;
  wire lt,eq,gt,unordered,N0,isNaNA,isInfA,isZeroA,signA,isSigNaNA,isNaNB,isInfB,
  isZeroB,signB,isSigNaNB,ordered,bothInfs,bothZeros,eqHiExps,N1,eqExps,N2,N3,N4,
  common_ltMags,N5,common_eqMags,ordered_lt,N6,ordered_eq,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31;
  wire [12:0] sExpA,sExpB;
  wire [53:0] sigA,sigB;
  assign exceptionFlags[0] = 1'b0;
  assign exceptionFlags[1] = 1'b0;
  assign exceptionFlags[2] = 1'b0;
  assign exceptionFlags[3] = 1'b0;

  recFNToRawFN_expWidth11_sigWidth53
  recFNToRawFN_a
  (
    .in(a),
    .isNaN(isNaNA),
    .isInf(isInfA),
    .isZero(isZeroA),
    .sign(signA),
    .sExp(sExpA),
    .sig(sigA)
  );


  isSigNaNRecFN_expWidth11_sigWidth53
  isSigNaN_a
  (
    .in(a),
    .isSigNaN(isSigNaNA)
  );


  recFNToRawFN_expWidth11_sigWidth53
  recFNToRawFN_b
  (
    .in(b),
    .isNaN(isNaNB),
    .isInf(isInfB),
    .isZero(isZeroB),
    .sign(signB),
    .sExp(sExpB),
    .sig(sigB)
  );


  isSigNaNRecFN_expWidth11_sigWidth53
  isSigNaN_b
  (
    .in(b),
    .isSigNaN(isSigNaNB)
  );

  assign eqHiExps = $signed({ 1'b0, sExpA[12:9] }) == $signed({ 1'b0, sExpB[12:9] });
  assign N1 = sExpA[8:0] == sExpB[8:0];
  assign N2 = $signed({ 1'b0, sExpA[12:9] }) < $signed({ 1'b0, sExpB[12:9] });
  assign N3 = sExpA[8:0] < sExpB[8:0];
  assign N4 = sigA < sigB;
  assign N5 = sigA == sigB;
  assign N0 = signA ^ signB;
  assign N6 = ~N0;
  assign ordered = N7 & N8;
  assign N7 = ~isNaNA;
  assign N8 = ~isNaNB;
  assign bothInfs = isInfA & isInfB;
  assign bothZeros = isZeroA & isZeroB;
  assign eqExps = eqHiExps & N1;
  assign common_ltMags = N10 | N11;
  assign N10 = N2 | N9;
  assign N9 = eqHiExps & N3;
  assign N11 = eqExps & N4;
  assign common_eqMags = eqExps & N5;
  assign ordered_lt = N12 & N23;
  assign N12 = ~bothZeros;
  assign N23 = N14 | N22;
  assign N14 = signA & N13;
  assign N13 = ~signB;
  assign N22 = N15 & N21;
  assign N15 = ~bothInfs;
  assign N21 = N19 | N20;
  assign N19 = N17 & N18;
  assign N17 = signA & N16;
  assign N16 = ~common_ltMags;
  assign N18 = ~common_eqMags;
  assign N20 = N13 & common_ltMags;
  assign ordered_eq = bothZeros | N25;
  assign N25 = N6 & N24;
  assign N24 = bothInfs | common_eqMags;
  assign exceptionFlags[4] = N26 | N28;
  assign N26 = isSigNaNA | isSigNaNB;
  assign N28 = signaling & N27;
  assign N27 = ~ordered;
  assign lt = ordered & ordered_lt;
  assign eq = ordered & ordered_eq;
  assign gt = N30 & N31;
  assign N30 = ordered & N29;
  assign N29 = ~ordered_lt;
  assign N31 = ~ordered_eq;
  assign unordered = ~ordered;

endmodule



module bsg_scan_width_p24_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [23:0] i;
  output [23:0] o;
  wire [23:0] o;
  wire t_4__23_,t_4__22_,t_4__21_,t_4__20_,t_4__19_,t_4__18_,t_4__17_,t_4__16_,
  t_4__15_,t_4__14_,t_4__13_,t_4__12_,t_4__11_,t_4__10_,t_4__9_,t_4__8_,t_4__7_,t_4__6_,
  t_4__5_,t_4__4_,t_4__3_,t_4__2_,t_4__1_,t_4__0_,t_3__23_,t_3__22_,t_3__21_,
  t_3__20_,t_3__19_,t_3__18_,t_3__17_,t_3__16_,t_3__15_,t_3__14_,t_3__13_,t_3__12_,
  t_3__11_,t_3__10_,t_3__9_,t_3__8_,t_3__7_,t_3__6_,t_3__5_,t_3__4_,t_3__3_,t_3__2_,
  t_3__1_,t_3__0_,t_2__23_,t_2__22_,t_2__21_,t_2__20_,t_2__19_,t_2__18_,t_2__17_,
  t_2__16_,t_2__15_,t_2__14_,t_2__13_,t_2__12_,t_2__11_,t_2__10_,t_2__9_,t_2__8_,
  t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__23_,t_1__22_,
  t_1__21_,t_1__20_,t_1__19_,t_1__18_,t_1__17_,t_1__16_,t_1__15_,t_1__14_,t_1__13_,
  t_1__12_,t_1__11_,t_1__10_,t_1__9_,t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,t_1__3_,
  t_1__2_,t_1__1_,t_1__0_;
  assign t_1__23_ = i[0] | 1'b0;
  assign t_1__22_ = i[1] | i[0];
  assign t_1__21_ = i[2] | i[1];
  assign t_1__20_ = i[3] | i[2];
  assign t_1__19_ = i[4] | i[3];
  assign t_1__18_ = i[5] | i[4];
  assign t_1__17_ = i[6] | i[5];
  assign t_1__16_ = i[7] | i[6];
  assign t_1__15_ = i[8] | i[7];
  assign t_1__14_ = i[9] | i[8];
  assign t_1__13_ = i[10] | i[9];
  assign t_1__12_ = i[11] | i[10];
  assign t_1__11_ = i[12] | i[11];
  assign t_1__10_ = i[13] | i[12];
  assign t_1__9_ = i[14] | i[13];
  assign t_1__8_ = i[15] | i[14];
  assign t_1__7_ = i[16] | i[15];
  assign t_1__6_ = i[17] | i[16];
  assign t_1__5_ = i[18] | i[17];
  assign t_1__4_ = i[19] | i[18];
  assign t_1__3_ = i[20] | i[19];
  assign t_1__2_ = i[21] | i[20];
  assign t_1__1_ = i[22] | i[21];
  assign t_1__0_ = i[23] | i[22];
  assign t_2__23_ = t_1__23_ | 1'b0;
  assign t_2__22_ = t_1__22_ | 1'b0;
  assign t_2__21_ = t_1__21_ | t_1__23_;
  assign t_2__20_ = t_1__20_ | t_1__22_;
  assign t_2__19_ = t_1__19_ | t_1__21_;
  assign t_2__18_ = t_1__18_ | t_1__20_;
  assign t_2__17_ = t_1__17_ | t_1__19_;
  assign t_2__16_ = t_1__16_ | t_1__18_;
  assign t_2__15_ = t_1__15_ | t_1__17_;
  assign t_2__14_ = t_1__14_ | t_1__16_;
  assign t_2__13_ = t_1__13_ | t_1__15_;
  assign t_2__12_ = t_1__12_ | t_1__14_;
  assign t_2__11_ = t_1__11_ | t_1__13_;
  assign t_2__10_ = t_1__10_ | t_1__12_;
  assign t_2__9_ = t_1__9_ | t_1__11_;
  assign t_2__8_ = t_1__8_ | t_1__10_;
  assign t_2__7_ = t_1__7_ | t_1__9_;
  assign t_2__6_ = t_1__6_ | t_1__8_;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign t_3__23_ = t_2__23_ | 1'b0;
  assign t_3__22_ = t_2__22_ | 1'b0;
  assign t_3__21_ = t_2__21_ | 1'b0;
  assign t_3__20_ = t_2__20_ | 1'b0;
  assign t_3__19_ = t_2__19_ | t_2__23_;
  assign t_3__18_ = t_2__18_ | t_2__22_;
  assign t_3__17_ = t_2__17_ | t_2__21_;
  assign t_3__16_ = t_2__16_ | t_2__20_;
  assign t_3__15_ = t_2__15_ | t_2__19_;
  assign t_3__14_ = t_2__14_ | t_2__18_;
  assign t_3__13_ = t_2__13_ | t_2__17_;
  assign t_3__12_ = t_2__12_ | t_2__16_;
  assign t_3__11_ = t_2__11_ | t_2__15_;
  assign t_3__10_ = t_2__10_ | t_2__14_;
  assign t_3__9_ = t_2__9_ | t_2__13_;
  assign t_3__8_ = t_2__8_ | t_2__12_;
  assign t_3__7_ = t_2__7_ | t_2__11_;
  assign t_3__6_ = t_2__6_ | t_2__10_;
  assign t_3__5_ = t_2__5_ | t_2__9_;
  assign t_3__4_ = t_2__4_ | t_2__8_;
  assign t_3__3_ = t_2__3_ | t_2__7_;
  assign t_3__2_ = t_2__2_ | t_2__6_;
  assign t_3__1_ = t_2__1_ | t_2__5_;
  assign t_3__0_ = t_2__0_ | t_2__4_;
  assign t_4__23_ = t_3__23_ | 1'b0;
  assign t_4__22_ = t_3__22_ | 1'b0;
  assign t_4__21_ = t_3__21_ | 1'b0;
  assign t_4__20_ = t_3__20_ | 1'b0;
  assign t_4__19_ = t_3__19_ | 1'b0;
  assign t_4__18_ = t_3__18_ | 1'b0;
  assign t_4__17_ = t_3__17_ | 1'b0;
  assign t_4__16_ = t_3__16_ | 1'b0;
  assign t_4__15_ = t_3__15_ | t_3__23_;
  assign t_4__14_ = t_3__14_ | t_3__22_;
  assign t_4__13_ = t_3__13_ | t_3__21_;
  assign t_4__12_ = t_3__12_ | t_3__20_;
  assign t_4__11_ = t_3__11_ | t_3__19_;
  assign t_4__10_ = t_3__10_ | t_3__18_;
  assign t_4__9_ = t_3__9_ | t_3__17_;
  assign t_4__8_ = t_3__8_ | t_3__16_;
  assign t_4__7_ = t_3__7_ | t_3__15_;
  assign t_4__6_ = t_3__6_ | t_3__14_;
  assign t_4__5_ = t_3__5_ | t_3__13_;
  assign t_4__4_ = t_3__4_ | t_3__12_;
  assign t_4__3_ = t_3__3_ | t_3__11_;
  assign t_4__2_ = t_3__2_ | t_3__10_;
  assign t_4__1_ = t_3__1_ | t_3__9_;
  assign t_4__0_ = t_3__0_ | t_3__8_;
  assign o[0] = t_4__23_ | 1'b0;
  assign o[1] = t_4__22_ | 1'b0;
  assign o[2] = t_4__21_ | 1'b0;
  assign o[3] = t_4__20_ | 1'b0;
  assign o[4] = t_4__19_ | 1'b0;
  assign o[5] = t_4__18_ | 1'b0;
  assign o[6] = t_4__17_ | 1'b0;
  assign o[7] = t_4__16_ | 1'b0;
  assign o[8] = t_4__15_ | 1'b0;
  assign o[9] = t_4__14_ | 1'b0;
  assign o[10] = t_4__13_ | 1'b0;
  assign o[11] = t_4__12_ | 1'b0;
  assign o[12] = t_4__11_ | 1'b0;
  assign o[13] = t_4__10_ | 1'b0;
  assign o[14] = t_4__9_ | 1'b0;
  assign o[15] = t_4__8_ | 1'b0;
  assign o[16] = t_4__7_ | t_4__23_;
  assign o[17] = t_4__6_ | t_4__22_;
  assign o[18] = t_4__5_ | t_4__21_;
  assign o[19] = t_4__4_ | t_4__20_;
  assign o[20] = t_4__3_ | t_4__19_;
  assign o[21] = t_4__2_ | t_4__18_;
  assign o[22] = t_4__1_ | t_4__17_;
  assign o[23] = t_4__0_ | t_4__16_;

endmodule



module bsg_priority_encode_one_hot_out_width_p24_lo_to_hi_p1
(
  i,
  o,
  v_o
);

  input [23:0] i;
  output [23:0] o;
  output v_o;
  wire [23:0] o;
  wire v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22;
  wire [22:1] scan_lo;

  bsg_scan_width_p24_or_p1_lo_to_hi_p1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, scan_lo, o[0:0] })
  );

  assign o[23] = v_o & N0;
  assign N0 = ~scan_lo[22];
  assign o[22] = scan_lo[22] & N1;
  assign N1 = ~scan_lo[21];
  assign o[21] = scan_lo[21] & N2;
  assign N2 = ~scan_lo[20];
  assign o[20] = scan_lo[20] & N3;
  assign N3 = ~scan_lo[19];
  assign o[19] = scan_lo[19] & N4;
  assign N4 = ~scan_lo[18];
  assign o[18] = scan_lo[18] & N5;
  assign N5 = ~scan_lo[17];
  assign o[17] = scan_lo[17] & N6;
  assign N6 = ~scan_lo[16];
  assign o[16] = scan_lo[16] & N7;
  assign N7 = ~scan_lo[15];
  assign o[15] = scan_lo[15] & N8;
  assign N8 = ~scan_lo[14];
  assign o[14] = scan_lo[14] & N9;
  assign N9 = ~scan_lo[13];
  assign o[13] = scan_lo[13] & N10;
  assign N10 = ~scan_lo[12];
  assign o[12] = scan_lo[12] & N11;
  assign N11 = ~scan_lo[11];
  assign o[11] = scan_lo[11] & N12;
  assign N12 = ~scan_lo[10];
  assign o[10] = scan_lo[10] & N13;
  assign N13 = ~scan_lo[9];
  assign o[9] = scan_lo[9] & N14;
  assign N14 = ~scan_lo[8];
  assign o[8] = scan_lo[8] & N15;
  assign N15 = ~scan_lo[7];
  assign o[7] = scan_lo[7] & N16;
  assign N16 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N17;
  assign N17 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N18;
  assign N18 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N19;
  assign N19 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N20;
  assign N20 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N21;
  assign N21 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N22;
  assign N22 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p24_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [23:0] i;
  output [4:0] addr_o;
  output v_o;
  wire [4:0] addr_o;
  wire v_o,v_4__0_,v_3__24_,v_3__16_,v_3__8_,v_3__0_,v_2__28_,v_2__24_,v_2__20_,
  v_2__16_,v_2__12_,v_2__8_,v_2__4_,v_2__0_,v_1__30_,v_1__28_,v_1__26_,v_1__24_,v_1__22_,
  v_1__20_,v_1__18_,v_1__16_,v_1__14_,v_1__12_,v_1__10_,v_1__8_,v_1__6_,v_1__4_,
  v_1__2_,v_1__0_,addr_4__18_,addr_4__17_,addr_4__16_,addr_4__2_,addr_4__1_,
  addr_4__0_,addr_3__25_,addr_3__24_,addr_3__17_,addr_3__16_,addr_3__9_,addr_3__8_,
  addr_3__1_,addr_3__0_,addr_2__28_,addr_2__24_,addr_2__20_,addr_2__16_,addr_2__12_,
  addr_2__8_,addr_2__4_,addr_2__0_;
  assign v_1__0_ = i[1] | i[0];
  assign v_1__2_ = i[3] | i[2];
  assign v_1__4_ = i[5] | i[4];
  assign v_1__6_ = i[7] | i[6];
  assign v_1__8_ = i[9] | i[8];
  assign v_1__10_ = i[11] | i[10];
  assign v_1__12_ = i[13] | i[12];
  assign v_1__14_ = i[15] | i[14];
  assign v_1__16_ = i[17] | i[16];
  assign v_1__18_ = i[19] | i[18];
  assign v_1__20_ = i[21] | i[20];
  assign v_1__22_ = i[23] | i[22];
  assign v_1__24_ = 1'b0 | 1'b0;
  assign v_1__26_ = 1'b0 | 1'b0;
  assign v_1__28_ = 1'b0 | 1'b0;
  assign v_1__30_ = 1'b0 | 1'b0;
  assign v_2__0_ = v_1__2_ | v_1__0_;
  assign addr_2__0_ = i[1] | i[3];
  assign v_2__4_ = v_1__6_ | v_1__4_;
  assign addr_2__4_ = i[5] | i[7];
  assign v_2__8_ = v_1__10_ | v_1__8_;
  assign addr_2__8_ = i[9] | i[11];
  assign v_2__12_ = v_1__14_ | v_1__12_;
  assign addr_2__12_ = i[13] | i[15];
  assign v_2__16_ = v_1__18_ | v_1__16_;
  assign addr_2__16_ = i[17] | i[19];
  assign v_2__20_ = v_1__22_ | v_1__20_;
  assign addr_2__20_ = i[21] | i[23];
  assign v_2__24_ = v_1__26_ | v_1__24_;
  assign addr_2__24_ = 1'b0 | 1'b0;
  assign v_2__28_ = v_1__30_ | v_1__28_;
  assign addr_2__28_ = 1'b0 | 1'b0;
  assign v_3__0_ = v_2__4_ | v_2__0_;
  assign addr_3__1_ = v_1__2_ | v_1__6_;
  assign addr_3__0_ = addr_2__0_ | addr_2__4_;
  assign v_3__8_ = v_2__12_ | v_2__8_;
  assign addr_3__9_ = v_1__10_ | v_1__14_;
  assign addr_3__8_ = addr_2__8_ | addr_2__12_;
  assign v_3__16_ = v_2__20_ | v_2__16_;
  assign addr_3__17_ = v_1__18_ | v_1__22_;
  assign addr_3__16_ = addr_2__16_ | addr_2__20_;
  assign v_3__24_ = v_2__28_ | v_2__24_;
  assign addr_3__25_ = v_1__26_ | v_1__30_;
  assign addr_3__24_ = addr_2__24_ | addr_2__28_;
  assign v_4__0_ = v_3__8_ | v_3__0_;
  assign addr_4__2_ = v_2__4_ | v_2__12_;
  assign addr_4__1_ = addr_3__1_ | addr_3__9_;
  assign addr_4__0_ = addr_3__0_ | addr_3__8_;
  assign addr_o[4] = v_3__24_ | v_3__16_;
  assign addr_4__18_ = v_2__20_ | v_2__28_;
  assign addr_4__17_ = addr_3__17_ | addr_3__25_;
  assign addr_4__16_ = addr_3__16_ | addr_3__24_;
  assign v_o = addr_o[4] | v_4__0_;
  assign addr_o[3] = v_3__8_ | v_3__24_;
  assign addr_o[2] = addr_4__2_ | addr_4__18_;
  assign addr_o[1] = addr_4__1_ | addr_4__17_;
  assign addr_o[0] = addr_4__0_ | addr_4__16_;

endmodule



module bsg_priority_encode_width_p24_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [23:0] i;
  output [4:0] addr_o;
  output v_o;
  wire [4:0] addr_o;
  wire v_o;
  wire [23:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p24_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_width_p24_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o)
  );


endmodule



module bsg_counting_leading_zeros_width_p23
(
  a_i,
  num_zero_o
);

  input [22:0] a_i;
  output [4:0] num_zero_o;
  wire [4:0] num_zero_o;

  bsg_priority_encode_width_p24_lo_to_hi_p1
  pe0
  (
    .i({ 1'b1, a_i[0:0], a_i[1:1], a_i[2:2], a_i[3:3], a_i[4:4], a_i[5:5], a_i[6:6], a_i[7:7], a_i[8:8], a_i[9:9], a_i[10:10], a_i[11:11], a_i[12:12], a_i[13:13], a_i[14:14], a_i[15:15], a_i[16:16], a_i[17:17], a_i[18:18], a_i[19:19], a_i[20:20], a_i[21:21], a_i[22:22] }),
    .addr_o(num_zero_o)
  );


endmodule



module fNToRecFN_expWidth8_sigWidth24
(
  in,
  out
);

  input [31:0] in;
  output [32:0] out;
  wire [32:0] out;
  wire N0,N1,N2,out_32_,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,isZero,isSpecial,
  N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,
  N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50;
  wire [4:0] normDist;
  wire [22:1] subnormFract;
  wire [8:6] adjustedExp;
  assign out_32_ = in[31];
  assign out[32] = out_32_;

  bsg_counting_leading_zeros_width_p23
  clz
  (
    .a_i(in[22:0]),
    .num_zero_o(normDist)
  );

  assign isSpecial = adjustedExp[8:7] == { 1'b1, 1'b1 };
  assign subnormFract = in[21:0] << normDist;
  assign N20 = in[21] | in[22];
  assign N21 = in[20] | N20;
  assign N22 = in[19] | N21;
  assign N23 = in[18] | N22;
  assign N24 = in[17] | N23;
  assign N25 = in[16] | N24;
  assign N26 = in[15] | N25;
  assign N27 = in[14] | N26;
  assign N28 = in[13] | N27;
  assign N29 = in[12] | N28;
  assign N30 = in[11] | N29;
  assign N31 = in[10] | N30;
  assign N32 = in[9] | N31;
  assign N33 = in[8] | N32;
  assign N34 = in[7] | N33;
  assign N35 = in[6] | N34;
  assign N36 = in[5] | N35;
  assign N37 = in[4] | N36;
  assign N38 = in[3] | N37;
  assign N39 = in[2] | N38;
  assign N40 = in[1] | N39;
  assign N41 = in[0] | N40;
  assign N42 = ~N41;
  assign N43 = in[29] | in[30];
  assign N44 = in[28] | N43;
  assign N45 = in[27] | N44;
  assign N46 = in[26] | N45;
  assign N47 = in[25] | N46;
  assign N48 = in[24] | N47;
  assign N49 = in[23] | N48;
  assign N50 = ~N49;
  assign { adjustedExp, out[28:23] } = { N50, N15, N14, N13, N12, N11, N10, N9, N8 } + { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N50, N49 };
  assign { N15, N14, N13, N12, N11, N10, N9, N8 } = (N0)? { 1'b1, 1'b1, 1'b1, N3, N4, N5, N6, N7 } : 
                                                    (N1)? in[30:23] : 1'b0;
  assign N0 = N50;
  assign N1 = N49;
  assign out[31:29] = (N2)? { 1'b1, 1'b1, N41 } : 
                      (N19)? { 1'b0, 1'b0, 1'b0 } : 
                      (N17)? adjustedExp : 1'b0;
  assign N2 = isSpecial;
  assign out[22:0] = (N0)? { subnormFract, 1'b0 } : 
                     (N1)? in[22:0] : 1'b0;
  assign N3 = ~normDist[4];
  assign N4 = ~normDist[3];
  assign N5 = ~normDist[2];
  assign N6 = ~normDist[1];
  assign N7 = ~normDist[0];
  assign isZero = N50 & N42;
  assign N16 = isZero | isSpecial;
  assign N17 = ~N16;
  assign N18 = ~isSpecial;
  assign N19 = isZero & N18;

endmodule



module bsg_scan_width_p53_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [52:0] i;
  output [52:0] o;
  wire [52:0] o;
  wire t_5__52_,t_5__51_,t_5__50_,t_5__49_,t_5__48_,t_5__47_,t_5__46_,t_5__45_,
  t_5__44_,t_5__43_,t_5__42_,t_5__41_,t_5__40_,t_5__39_,t_5__38_,t_5__37_,t_5__36_,
  t_5__35_,t_5__34_,t_5__33_,t_5__32_,t_5__31_,t_5__30_,t_5__29_,t_5__28_,t_5__27_,
  t_5__26_,t_5__25_,t_5__24_,t_5__23_,t_5__22_,t_5__21_,t_5__20_,t_5__19_,t_5__18_,
  t_5__17_,t_5__16_,t_5__15_,t_5__14_,t_5__13_,t_5__12_,t_5__11_,t_5__10_,t_5__9_,
  t_5__8_,t_5__7_,t_5__6_,t_5__5_,t_5__4_,t_5__3_,t_5__2_,t_5__1_,t_5__0_,t_4__52_,
  t_4__51_,t_4__50_,t_4__49_,t_4__48_,t_4__47_,t_4__46_,t_4__45_,t_4__44_,t_4__43_,
  t_4__42_,t_4__41_,t_4__40_,t_4__39_,t_4__38_,t_4__37_,t_4__36_,t_4__35_,t_4__34_,
  t_4__33_,t_4__32_,t_4__31_,t_4__30_,t_4__29_,t_4__28_,t_4__27_,t_4__26_,t_4__25_,
  t_4__24_,t_4__23_,t_4__22_,t_4__21_,t_4__20_,t_4__19_,t_4__18_,t_4__17_,t_4__16_,
  t_4__15_,t_4__14_,t_4__13_,t_4__12_,t_4__11_,t_4__10_,t_4__9_,t_4__8_,t_4__7_,
  t_4__6_,t_4__5_,t_4__4_,t_4__3_,t_4__2_,t_4__1_,t_4__0_,t_3__52_,t_3__51_,
  t_3__50_,t_3__49_,t_3__48_,t_3__47_,t_3__46_,t_3__45_,t_3__44_,t_3__43_,t_3__42_,
  t_3__41_,t_3__40_,t_3__39_,t_3__38_,t_3__37_,t_3__36_,t_3__35_,t_3__34_,t_3__33_,
  t_3__32_,t_3__31_,t_3__30_,t_3__29_,t_3__28_,t_3__27_,t_3__26_,t_3__25_,t_3__24_,
  t_3__23_,t_3__22_,t_3__21_,t_3__20_,t_3__19_,t_3__18_,t_3__17_,t_3__16_,t_3__15_,
  t_3__14_,t_3__13_,t_3__12_,t_3__11_,t_3__10_,t_3__9_,t_3__8_,t_3__7_,t_3__6_,
  t_3__5_,t_3__4_,t_3__3_,t_3__2_,t_3__1_,t_3__0_,t_2__52_,t_2__51_,t_2__50_,t_2__49_,
  t_2__48_,t_2__47_,t_2__46_,t_2__45_,t_2__44_,t_2__43_,t_2__42_,t_2__41_,t_2__40_,
  t_2__39_,t_2__38_,t_2__37_,t_2__36_,t_2__35_,t_2__34_,t_2__33_,t_2__32_,t_2__31_,
  t_2__30_,t_2__29_,t_2__28_,t_2__27_,t_2__26_,t_2__25_,t_2__24_,t_2__23_,t_2__22_,
  t_2__21_,t_2__20_,t_2__19_,t_2__18_,t_2__17_,t_2__16_,t_2__15_,t_2__14_,
  t_2__13_,t_2__12_,t_2__11_,t_2__10_,t_2__9_,t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,
  t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__52_,t_1__51_,t_1__50_,t_1__49_,t_1__48_,
  t_1__47_,t_1__46_,t_1__45_,t_1__44_,t_1__43_,t_1__42_,t_1__41_,t_1__40_,t_1__39_,
  t_1__38_,t_1__37_,t_1__36_,t_1__35_,t_1__34_,t_1__33_,t_1__32_,t_1__31_,t_1__30_,
  t_1__29_,t_1__28_,t_1__27_,t_1__26_,t_1__25_,t_1__24_,t_1__23_,t_1__22_,t_1__21_,
  t_1__20_,t_1__19_,t_1__18_,t_1__17_,t_1__16_,t_1__15_,t_1__14_,t_1__13_,t_1__12_,
  t_1__11_,t_1__10_,t_1__9_,t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,
  t_1__1_,t_1__0_;
  assign t_1__52_ = i[0] | 1'b0;
  assign t_1__51_ = i[1] | i[0];
  assign t_1__50_ = i[2] | i[1];
  assign t_1__49_ = i[3] | i[2];
  assign t_1__48_ = i[4] | i[3];
  assign t_1__47_ = i[5] | i[4];
  assign t_1__46_ = i[6] | i[5];
  assign t_1__45_ = i[7] | i[6];
  assign t_1__44_ = i[8] | i[7];
  assign t_1__43_ = i[9] | i[8];
  assign t_1__42_ = i[10] | i[9];
  assign t_1__41_ = i[11] | i[10];
  assign t_1__40_ = i[12] | i[11];
  assign t_1__39_ = i[13] | i[12];
  assign t_1__38_ = i[14] | i[13];
  assign t_1__37_ = i[15] | i[14];
  assign t_1__36_ = i[16] | i[15];
  assign t_1__35_ = i[17] | i[16];
  assign t_1__34_ = i[18] | i[17];
  assign t_1__33_ = i[19] | i[18];
  assign t_1__32_ = i[20] | i[19];
  assign t_1__31_ = i[21] | i[20];
  assign t_1__30_ = i[22] | i[21];
  assign t_1__29_ = i[23] | i[22];
  assign t_1__28_ = i[24] | i[23];
  assign t_1__27_ = i[25] | i[24];
  assign t_1__26_ = i[26] | i[25];
  assign t_1__25_ = i[27] | i[26];
  assign t_1__24_ = i[28] | i[27];
  assign t_1__23_ = i[29] | i[28];
  assign t_1__22_ = i[30] | i[29];
  assign t_1__21_ = i[31] | i[30];
  assign t_1__20_ = i[32] | i[31];
  assign t_1__19_ = i[33] | i[32];
  assign t_1__18_ = i[34] | i[33];
  assign t_1__17_ = i[35] | i[34];
  assign t_1__16_ = i[36] | i[35];
  assign t_1__15_ = i[37] | i[36];
  assign t_1__14_ = i[38] | i[37];
  assign t_1__13_ = i[39] | i[38];
  assign t_1__12_ = i[40] | i[39];
  assign t_1__11_ = i[41] | i[40];
  assign t_1__10_ = i[42] | i[41];
  assign t_1__9_ = i[43] | i[42];
  assign t_1__8_ = i[44] | i[43];
  assign t_1__7_ = i[45] | i[44];
  assign t_1__6_ = i[46] | i[45];
  assign t_1__5_ = i[47] | i[46];
  assign t_1__4_ = i[48] | i[47];
  assign t_1__3_ = i[49] | i[48];
  assign t_1__2_ = i[50] | i[49];
  assign t_1__1_ = i[51] | i[50];
  assign t_1__0_ = i[52] | i[51];
  assign t_2__52_ = t_1__52_ | 1'b0;
  assign t_2__51_ = t_1__51_ | 1'b0;
  assign t_2__50_ = t_1__50_ | t_1__52_;
  assign t_2__49_ = t_1__49_ | t_1__51_;
  assign t_2__48_ = t_1__48_ | t_1__50_;
  assign t_2__47_ = t_1__47_ | t_1__49_;
  assign t_2__46_ = t_1__46_ | t_1__48_;
  assign t_2__45_ = t_1__45_ | t_1__47_;
  assign t_2__44_ = t_1__44_ | t_1__46_;
  assign t_2__43_ = t_1__43_ | t_1__45_;
  assign t_2__42_ = t_1__42_ | t_1__44_;
  assign t_2__41_ = t_1__41_ | t_1__43_;
  assign t_2__40_ = t_1__40_ | t_1__42_;
  assign t_2__39_ = t_1__39_ | t_1__41_;
  assign t_2__38_ = t_1__38_ | t_1__40_;
  assign t_2__37_ = t_1__37_ | t_1__39_;
  assign t_2__36_ = t_1__36_ | t_1__38_;
  assign t_2__35_ = t_1__35_ | t_1__37_;
  assign t_2__34_ = t_1__34_ | t_1__36_;
  assign t_2__33_ = t_1__33_ | t_1__35_;
  assign t_2__32_ = t_1__32_ | t_1__34_;
  assign t_2__31_ = t_1__31_ | t_1__33_;
  assign t_2__30_ = t_1__30_ | t_1__32_;
  assign t_2__29_ = t_1__29_ | t_1__31_;
  assign t_2__28_ = t_1__28_ | t_1__30_;
  assign t_2__27_ = t_1__27_ | t_1__29_;
  assign t_2__26_ = t_1__26_ | t_1__28_;
  assign t_2__25_ = t_1__25_ | t_1__27_;
  assign t_2__24_ = t_1__24_ | t_1__26_;
  assign t_2__23_ = t_1__23_ | t_1__25_;
  assign t_2__22_ = t_1__22_ | t_1__24_;
  assign t_2__21_ = t_1__21_ | t_1__23_;
  assign t_2__20_ = t_1__20_ | t_1__22_;
  assign t_2__19_ = t_1__19_ | t_1__21_;
  assign t_2__18_ = t_1__18_ | t_1__20_;
  assign t_2__17_ = t_1__17_ | t_1__19_;
  assign t_2__16_ = t_1__16_ | t_1__18_;
  assign t_2__15_ = t_1__15_ | t_1__17_;
  assign t_2__14_ = t_1__14_ | t_1__16_;
  assign t_2__13_ = t_1__13_ | t_1__15_;
  assign t_2__12_ = t_1__12_ | t_1__14_;
  assign t_2__11_ = t_1__11_ | t_1__13_;
  assign t_2__10_ = t_1__10_ | t_1__12_;
  assign t_2__9_ = t_1__9_ | t_1__11_;
  assign t_2__8_ = t_1__8_ | t_1__10_;
  assign t_2__7_ = t_1__7_ | t_1__9_;
  assign t_2__6_ = t_1__6_ | t_1__8_;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign t_3__52_ = t_2__52_ | 1'b0;
  assign t_3__51_ = t_2__51_ | 1'b0;
  assign t_3__50_ = t_2__50_ | 1'b0;
  assign t_3__49_ = t_2__49_ | 1'b0;
  assign t_3__48_ = t_2__48_ | t_2__52_;
  assign t_3__47_ = t_2__47_ | t_2__51_;
  assign t_3__46_ = t_2__46_ | t_2__50_;
  assign t_3__45_ = t_2__45_ | t_2__49_;
  assign t_3__44_ = t_2__44_ | t_2__48_;
  assign t_3__43_ = t_2__43_ | t_2__47_;
  assign t_3__42_ = t_2__42_ | t_2__46_;
  assign t_3__41_ = t_2__41_ | t_2__45_;
  assign t_3__40_ = t_2__40_ | t_2__44_;
  assign t_3__39_ = t_2__39_ | t_2__43_;
  assign t_3__38_ = t_2__38_ | t_2__42_;
  assign t_3__37_ = t_2__37_ | t_2__41_;
  assign t_3__36_ = t_2__36_ | t_2__40_;
  assign t_3__35_ = t_2__35_ | t_2__39_;
  assign t_3__34_ = t_2__34_ | t_2__38_;
  assign t_3__33_ = t_2__33_ | t_2__37_;
  assign t_3__32_ = t_2__32_ | t_2__36_;
  assign t_3__31_ = t_2__31_ | t_2__35_;
  assign t_3__30_ = t_2__30_ | t_2__34_;
  assign t_3__29_ = t_2__29_ | t_2__33_;
  assign t_3__28_ = t_2__28_ | t_2__32_;
  assign t_3__27_ = t_2__27_ | t_2__31_;
  assign t_3__26_ = t_2__26_ | t_2__30_;
  assign t_3__25_ = t_2__25_ | t_2__29_;
  assign t_3__24_ = t_2__24_ | t_2__28_;
  assign t_3__23_ = t_2__23_ | t_2__27_;
  assign t_3__22_ = t_2__22_ | t_2__26_;
  assign t_3__21_ = t_2__21_ | t_2__25_;
  assign t_3__20_ = t_2__20_ | t_2__24_;
  assign t_3__19_ = t_2__19_ | t_2__23_;
  assign t_3__18_ = t_2__18_ | t_2__22_;
  assign t_3__17_ = t_2__17_ | t_2__21_;
  assign t_3__16_ = t_2__16_ | t_2__20_;
  assign t_3__15_ = t_2__15_ | t_2__19_;
  assign t_3__14_ = t_2__14_ | t_2__18_;
  assign t_3__13_ = t_2__13_ | t_2__17_;
  assign t_3__12_ = t_2__12_ | t_2__16_;
  assign t_3__11_ = t_2__11_ | t_2__15_;
  assign t_3__10_ = t_2__10_ | t_2__14_;
  assign t_3__9_ = t_2__9_ | t_2__13_;
  assign t_3__8_ = t_2__8_ | t_2__12_;
  assign t_3__7_ = t_2__7_ | t_2__11_;
  assign t_3__6_ = t_2__6_ | t_2__10_;
  assign t_3__5_ = t_2__5_ | t_2__9_;
  assign t_3__4_ = t_2__4_ | t_2__8_;
  assign t_3__3_ = t_2__3_ | t_2__7_;
  assign t_3__2_ = t_2__2_ | t_2__6_;
  assign t_3__1_ = t_2__1_ | t_2__5_;
  assign t_3__0_ = t_2__0_ | t_2__4_;
  assign t_4__52_ = t_3__52_ | 1'b0;
  assign t_4__51_ = t_3__51_ | 1'b0;
  assign t_4__50_ = t_3__50_ | 1'b0;
  assign t_4__49_ = t_3__49_ | 1'b0;
  assign t_4__48_ = t_3__48_ | 1'b0;
  assign t_4__47_ = t_3__47_ | 1'b0;
  assign t_4__46_ = t_3__46_ | 1'b0;
  assign t_4__45_ = t_3__45_ | 1'b0;
  assign t_4__44_ = t_3__44_ | t_3__52_;
  assign t_4__43_ = t_3__43_ | t_3__51_;
  assign t_4__42_ = t_3__42_ | t_3__50_;
  assign t_4__41_ = t_3__41_ | t_3__49_;
  assign t_4__40_ = t_3__40_ | t_3__48_;
  assign t_4__39_ = t_3__39_ | t_3__47_;
  assign t_4__38_ = t_3__38_ | t_3__46_;
  assign t_4__37_ = t_3__37_ | t_3__45_;
  assign t_4__36_ = t_3__36_ | t_3__44_;
  assign t_4__35_ = t_3__35_ | t_3__43_;
  assign t_4__34_ = t_3__34_ | t_3__42_;
  assign t_4__33_ = t_3__33_ | t_3__41_;
  assign t_4__32_ = t_3__32_ | t_3__40_;
  assign t_4__31_ = t_3__31_ | t_3__39_;
  assign t_4__30_ = t_3__30_ | t_3__38_;
  assign t_4__29_ = t_3__29_ | t_3__37_;
  assign t_4__28_ = t_3__28_ | t_3__36_;
  assign t_4__27_ = t_3__27_ | t_3__35_;
  assign t_4__26_ = t_3__26_ | t_3__34_;
  assign t_4__25_ = t_3__25_ | t_3__33_;
  assign t_4__24_ = t_3__24_ | t_3__32_;
  assign t_4__23_ = t_3__23_ | t_3__31_;
  assign t_4__22_ = t_3__22_ | t_3__30_;
  assign t_4__21_ = t_3__21_ | t_3__29_;
  assign t_4__20_ = t_3__20_ | t_3__28_;
  assign t_4__19_ = t_3__19_ | t_3__27_;
  assign t_4__18_ = t_3__18_ | t_3__26_;
  assign t_4__17_ = t_3__17_ | t_3__25_;
  assign t_4__16_ = t_3__16_ | t_3__24_;
  assign t_4__15_ = t_3__15_ | t_3__23_;
  assign t_4__14_ = t_3__14_ | t_3__22_;
  assign t_4__13_ = t_3__13_ | t_3__21_;
  assign t_4__12_ = t_3__12_ | t_3__20_;
  assign t_4__11_ = t_3__11_ | t_3__19_;
  assign t_4__10_ = t_3__10_ | t_3__18_;
  assign t_4__9_ = t_3__9_ | t_3__17_;
  assign t_4__8_ = t_3__8_ | t_3__16_;
  assign t_4__7_ = t_3__7_ | t_3__15_;
  assign t_4__6_ = t_3__6_ | t_3__14_;
  assign t_4__5_ = t_3__5_ | t_3__13_;
  assign t_4__4_ = t_3__4_ | t_3__12_;
  assign t_4__3_ = t_3__3_ | t_3__11_;
  assign t_4__2_ = t_3__2_ | t_3__10_;
  assign t_4__1_ = t_3__1_ | t_3__9_;
  assign t_4__0_ = t_3__0_ | t_3__8_;
  assign t_5__52_ = t_4__52_ | 1'b0;
  assign t_5__51_ = t_4__51_ | 1'b0;
  assign t_5__50_ = t_4__50_ | 1'b0;
  assign t_5__49_ = t_4__49_ | 1'b0;
  assign t_5__48_ = t_4__48_ | 1'b0;
  assign t_5__47_ = t_4__47_ | 1'b0;
  assign t_5__46_ = t_4__46_ | 1'b0;
  assign t_5__45_ = t_4__45_ | 1'b0;
  assign t_5__44_ = t_4__44_ | 1'b0;
  assign t_5__43_ = t_4__43_ | 1'b0;
  assign t_5__42_ = t_4__42_ | 1'b0;
  assign t_5__41_ = t_4__41_ | 1'b0;
  assign t_5__40_ = t_4__40_ | 1'b0;
  assign t_5__39_ = t_4__39_ | 1'b0;
  assign t_5__38_ = t_4__38_ | 1'b0;
  assign t_5__37_ = t_4__37_ | 1'b0;
  assign t_5__36_ = t_4__36_ | t_4__52_;
  assign t_5__35_ = t_4__35_ | t_4__51_;
  assign t_5__34_ = t_4__34_ | t_4__50_;
  assign t_5__33_ = t_4__33_ | t_4__49_;
  assign t_5__32_ = t_4__32_ | t_4__48_;
  assign t_5__31_ = t_4__31_ | t_4__47_;
  assign t_5__30_ = t_4__30_ | t_4__46_;
  assign t_5__29_ = t_4__29_ | t_4__45_;
  assign t_5__28_ = t_4__28_ | t_4__44_;
  assign t_5__27_ = t_4__27_ | t_4__43_;
  assign t_5__26_ = t_4__26_ | t_4__42_;
  assign t_5__25_ = t_4__25_ | t_4__41_;
  assign t_5__24_ = t_4__24_ | t_4__40_;
  assign t_5__23_ = t_4__23_ | t_4__39_;
  assign t_5__22_ = t_4__22_ | t_4__38_;
  assign t_5__21_ = t_4__21_ | t_4__37_;
  assign t_5__20_ = t_4__20_ | t_4__36_;
  assign t_5__19_ = t_4__19_ | t_4__35_;
  assign t_5__18_ = t_4__18_ | t_4__34_;
  assign t_5__17_ = t_4__17_ | t_4__33_;
  assign t_5__16_ = t_4__16_ | t_4__32_;
  assign t_5__15_ = t_4__15_ | t_4__31_;
  assign t_5__14_ = t_4__14_ | t_4__30_;
  assign t_5__13_ = t_4__13_ | t_4__29_;
  assign t_5__12_ = t_4__12_ | t_4__28_;
  assign t_5__11_ = t_4__11_ | t_4__27_;
  assign t_5__10_ = t_4__10_ | t_4__26_;
  assign t_5__9_ = t_4__9_ | t_4__25_;
  assign t_5__8_ = t_4__8_ | t_4__24_;
  assign t_5__7_ = t_4__7_ | t_4__23_;
  assign t_5__6_ = t_4__6_ | t_4__22_;
  assign t_5__5_ = t_4__5_ | t_4__21_;
  assign t_5__4_ = t_4__4_ | t_4__20_;
  assign t_5__3_ = t_4__3_ | t_4__19_;
  assign t_5__2_ = t_4__2_ | t_4__18_;
  assign t_5__1_ = t_4__1_ | t_4__17_;
  assign t_5__0_ = t_4__0_ | t_4__16_;
  assign o[0] = t_5__52_ | 1'b0;
  assign o[1] = t_5__51_ | 1'b0;
  assign o[2] = t_5__50_ | 1'b0;
  assign o[3] = t_5__49_ | 1'b0;
  assign o[4] = t_5__48_ | 1'b0;
  assign o[5] = t_5__47_ | 1'b0;
  assign o[6] = t_5__46_ | 1'b0;
  assign o[7] = t_5__45_ | 1'b0;
  assign o[8] = t_5__44_ | 1'b0;
  assign o[9] = t_5__43_ | 1'b0;
  assign o[10] = t_5__42_ | 1'b0;
  assign o[11] = t_5__41_ | 1'b0;
  assign o[12] = t_5__40_ | 1'b0;
  assign o[13] = t_5__39_ | 1'b0;
  assign o[14] = t_5__38_ | 1'b0;
  assign o[15] = t_5__37_ | 1'b0;
  assign o[16] = t_5__36_ | 1'b0;
  assign o[17] = t_5__35_ | 1'b0;
  assign o[18] = t_5__34_ | 1'b0;
  assign o[19] = t_5__33_ | 1'b0;
  assign o[20] = t_5__32_ | 1'b0;
  assign o[21] = t_5__31_ | 1'b0;
  assign o[22] = t_5__30_ | 1'b0;
  assign o[23] = t_5__29_ | 1'b0;
  assign o[24] = t_5__28_ | 1'b0;
  assign o[25] = t_5__27_ | 1'b0;
  assign o[26] = t_5__26_ | 1'b0;
  assign o[27] = t_5__25_ | 1'b0;
  assign o[28] = t_5__24_ | 1'b0;
  assign o[29] = t_5__23_ | 1'b0;
  assign o[30] = t_5__22_ | 1'b0;
  assign o[31] = t_5__21_ | 1'b0;
  assign o[32] = t_5__20_ | t_5__52_;
  assign o[33] = t_5__19_ | t_5__51_;
  assign o[34] = t_5__18_ | t_5__50_;
  assign o[35] = t_5__17_ | t_5__49_;
  assign o[36] = t_5__16_ | t_5__48_;
  assign o[37] = t_5__15_ | t_5__47_;
  assign o[38] = t_5__14_ | t_5__46_;
  assign o[39] = t_5__13_ | t_5__45_;
  assign o[40] = t_5__12_ | t_5__44_;
  assign o[41] = t_5__11_ | t_5__43_;
  assign o[42] = t_5__10_ | t_5__42_;
  assign o[43] = t_5__9_ | t_5__41_;
  assign o[44] = t_5__8_ | t_5__40_;
  assign o[45] = t_5__7_ | t_5__39_;
  assign o[46] = t_5__6_ | t_5__38_;
  assign o[47] = t_5__5_ | t_5__37_;
  assign o[48] = t_5__4_ | t_5__36_;
  assign o[49] = t_5__3_ | t_5__35_;
  assign o[50] = t_5__2_ | t_5__34_;
  assign o[51] = t_5__1_ | t_5__33_;
  assign o[52] = t_5__0_ | t_5__32_;

endmodule



module bsg_priority_encode_one_hot_out_width_p53_lo_to_hi_p1
(
  i,
  o,
  v_o
);

  input [52:0] i;
  output [52:0] o;
  output v_o;
  wire [52:0] o;
  wire v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51;
  wire [51:1] scan_lo;

  bsg_scan_width_p53_or_p1_lo_to_hi_p1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, scan_lo, o[0:0] })
  );

  assign o[52] = v_o & N0;
  assign N0 = ~scan_lo[51];
  assign o[51] = scan_lo[51] & N1;
  assign N1 = ~scan_lo[50];
  assign o[50] = scan_lo[50] & N2;
  assign N2 = ~scan_lo[49];
  assign o[49] = scan_lo[49] & N3;
  assign N3 = ~scan_lo[48];
  assign o[48] = scan_lo[48] & N4;
  assign N4 = ~scan_lo[47];
  assign o[47] = scan_lo[47] & N5;
  assign N5 = ~scan_lo[46];
  assign o[46] = scan_lo[46] & N6;
  assign N6 = ~scan_lo[45];
  assign o[45] = scan_lo[45] & N7;
  assign N7 = ~scan_lo[44];
  assign o[44] = scan_lo[44] & N8;
  assign N8 = ~scan_lo[43];
  assign o[43] = scan_lo[43] & N9;
  assign N9 = ~scan_lo[42];
  assign o[42] = scan_lo[42] & N10;
  assign N10 = ~scan_lo[41];
  assign o[41] = scan_lo[41] & N11;
  assign N11 = ~scan_lo[40];
  assign o[40] = scan_lo[40] & N12;
  assign N12 = ~scan_lo[39];
  assign o[39] = scan_lo[39] & N13;
  assign N13 = ~scan_lo[38];
  assign o[38] = scan_lo[38] & N14;
  assign N14 = ~scan_lo[37];
  assign o[37] = scan_lo[37] & N15;
  assign N15 = ~scan_lo[36];
  assign o[36] = scan_lo[36] & N16;
  assign N16 = ~scan_lo[35];
  assign o[35] = scan_lo[35] & N17;
  assign N17 = ~scan_lo[34];
  assign o[34] = scan_lo[34] & N18;
  assign N18 = ~scan_lo[33];
  assign o[33] = scan_lo[33] & N19;
  assign N19 = ~scan_lo[32];
  assign o[32] = scan_lo[32] & N20;
  assign N20 = ~scan_lo[31];
  assign o[31] = scan_lo[31] & N21;
  assign N21 = ~scan_lo[30];
  assign o[30] = scan_lo[30] & N22;
  assign N22 = ~scan_lo[29];
  assign o[29] = scan_lo[29] & N23;
  assign N23 = ~scan_lo[28];
  assign o[28] = scan_lo[28] & N24;
  assign N24 = ~scan_lo[27];
  assign o[27] = scan_lo[27] & N25;
  assign N25 = ~scan_lo[26];
  assign o[26] = scan_lo[26] & N26;
  assign N26 = ~scan_lo[25];
  assign o[25] = scan_lo[25] & N27;
  assign N27 = ~scan_lo[24];
  assign o[24] = scan_lo[24] & N28;
  assign N28 = ~scan_lo[23];
  assign o[23] = scan_lo[23] & N29;
  assign N29 = ~scan_lo[22];
  assign o[22] = scan_lo[22] & N30;
  assign N30 = ~scan_lo[21];
  assign o[21] = scan_lo[21] & N31;
  assign N31 = ~scan_lo[20];
  assign o[20] = scan_lo[20] & N32;
  assign N32 = ~scan_lo[19];
  assign o[19] = scan_lo[19] & N33;
  assign N33 = ~scan_lo[18];
  assign o[18] = scan_lo[18] & N34;
  assign N34 = ~scan_lo[17];
  assign o[17] = scan_lo[17] & N35;
  assign N35 = ~scan_lo[16];
  assign o[16] = scan_lo[16] & N36;
  assign N36 = ~scan_lo[15];
  assign o[15] = scan_lo[15] & N37;
  assign N37 = ~scan_lo[14];
  assign o[14] = scan_lo[14] & N38;
  assign N38 = ~scan_lo[13];
  assign o[13] = scan_lo[13] & N39;
  assign N39 = ~scan_lo[12];
  assign o[12] = scan_lo[12] & N40;
  assign N40 = ~scan_lo[11];
  assign o[11] = scan_lo[11] & N41;
  assign N41 = ~scan_lo[10];
  assign o[10] = scan_lo[10] & N42;
  assign N42 = ~scan_lo[9];
  assign o[9] = scan_lo[9] & N43;
  assign N43 = ~scan_lo[8];
  assign o[8] = scan_lo[8] & N44;
  assign N44 = ~scan_lo[7];
  assign o[7] = scan_lo[7] & N45;
  assign N45 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N46;
  assign N46 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N47;
  assign N47 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N48;
  assign N48 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N49;
  assign N49 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N50;
  assign N50 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N51;
  assign N51 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p53_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [52:0] i;
  output [5:0] addr_o;
  output v_o;
  wire [5:0] addr_o;
  wire v_o,v_5__0_,v_4__48_,v_4__32_,v_4__16_,v_4__0_,v_3__56_,v_3__48_,v_3__40_,
  v_3__32_,v_3__24_,v_3__16_,v_3__8_,v_3__0_,v_2__60_,v_2__56_,v_2__52_,v_2__48_,
  v_2__44_,v_2__40_,v_2__36_,v_2__32_,v_2__28_,v_2__24_,v_2__20_,v_2__16_,v_2__12_,
  v_2__8_,v_2__4_,v_2__0_,v_1__62_,v_1__60_,v_1__58_,v_1__56_,v_1__54_,v_1__52_,
  v_1__50_,v_1__48_,v_1__46_,v_1__44_,v_1__42_,v_1__40_,v_1__38_,v_1__36_,v_1__34_,
  v_1__32_,v_1__30_,v_1__28_,v_1__26_,v_1__24_,v_1__22_,v_1__20_,v_1__18_,v_1__16_,
  v_1__14_,v_1__12_,v_1__10_,v_1__8_,v_1__6_,v_1__4_,v_1__2_,v_1__0_,addr_5__35_,
  addr_5__34_,addr_5__33_,addr_5__32_,addr_5__3_,addr_5__2_,addr_5__1_,addr_5__0_,
  addr_4__50_,addr_4__49_,addr_4__48_,addr_4__34_,addr_4__33_,addr_4__32_,addr_4__18_,
  addr_4__17_,addr_4__16_,addr_4__2_,addr_4__1_,addr_4__0_,addr_3__57_,addr_3__56_,
  addr_3__49_,addr_3__48_,addr_3__41_,addr_3__40_,addr_3__33_,addr_3__32_,
  addr_3__25_,addr_3__24_,addr_3__17_,addr_3__16_,addr_3__9_,addr_3__8_,addr_3__1_,
  addr_3__0_,addr_2__60_,addr_2__56_,addr_2__52_,addr_2__48_,addr_2__44_,addr_2__40_,
  addr_2__36_,addr_2__32_,addr_2__28_,addr_2__24_,addr_2__20_,addr_2__16_,addr_2__12_,
  addr_2__8_,addr_2__4_,addr_2__0_;
  assign v_1__0_ = i[1] | i[0];
  assign v_1__2_ = i[3] | i[2];
  assign v_1__4_ = i[5] | i[4];
  assign v_1__6_ = i[7] | i[6];
  assign v_1__8_ = i[9] | i[8];
  assign v_1__10_ = i[11] | i[10];
  assign v_1__12_ = i[13] | i[12];
  assign v_1__14_ = i[15] | i[14];
  assign v_1__16_ = i[17] | i[16];
  assign v_1__18_ = i[19] | i[18];
  assign v_1__20_ = i[21] | i[20];
  assign v_1__22_ = i[23] | i[22];
  assign v_1__24_ = i[25] | i[24];
  assign v_1__26_ = i[27] | i[26];
  assign v_1__28_ = i[29] | i[28];
  assign v_1__30_ = i[31] | i[30];
  assign v_1__32_ = i[33] | i[32];
  assign v_1__34_ = i[35] | i[34];
  assign v_1__36_ = i[37] | i[36];
  assign v_1__38_ = i[39] | i[38];
  assign v_1__40_ = i[41] | i[40];
  assign v_1__42_ = i[43] | i[42];
  assign v_1__44_ = i[45] | i[44];
  assign v_1__46_ = i[47] | i[46];
  assign v_1__48_ = i[49] | i[48];
  assign v_1__50_ = i[51] | i[50];
  assign v_1__52_ = 1'b0 | i[52];
  assign v_1__54_ = 1'b0 | 1'b0;
  assign v_1__56_ = 1'b0 | 1'b0;
  assign v_1__58_ = 1'b0 | 1'b0;
  assign v_1__60_ = 1'b0 | 1'b0;
  assign v_1__62_ = 1'b0 | 1'b0;
  assign v_2__0_ = v_1__2_ | v_1__0_;
  assign addr_2__0_ = i[1] | i[3];
  assign v_2__4_ = v_1__6_ | v_1__4_;
  assign addr_2__4_ = i[5] | i[7];
  assign v_2__8_ = v_1__10_ | v_1__8_;
  assign addr_2__8_ = i[9] | i[11];
  assign v_2__12_ = v_1__14_ | v_1__12_;
  assign addr_2__12_ = i[13] | i[15];
  assign v_2__16_ = v_1__18_ | v_1__16_;
  assign addr_2__16_ = i[17] | i[19];
  assign v_2__20_ = v_1__22_ | v_1__20_;
  assign addr_2__20_ = i[21] | i[23];
  assign v_2__24_ = v_1__26_ | v_1__24_;
  assign addr_2__24_ = i[25] | i[27];
  assign v_2__28_ = v_1__30_ | v_1__28_;
  assign addr_2__28_ = i[29] | i[31];
  assign v_2__32_ = v_1__34_ | v_1__32_;
  assign addr_2__32_ = i[33] | i[35];
  assign v_2__36_ = v_1__38_ | v_1__36_;
  assign addr_2__36_ = i[37] | i[39];
  assign v_2__40_ = v_1__42_ | v_1__40_;
  assign addr_2__40_ = i[41] | i[43];
  assign v_2__44_ = v_1__46_ | v_1__44_;
  assign addr_2__44_ = i[45] | i[47];
  assign v_2__48_ = v_1__50_ | v_1__48_;
  assign addr_2__48_ = i[49] | i[51];
  assign v_2__52_ = v_1__54_ | v_1__52_;
  assign addr_2__52_ = 1'b0 | 1'b0;
  assign v_2__56_ = v_1__58_ | v_1__56_;
  assign addr_2__56_ = 1'b0 | 1'b0;
  assign v_2__60_ = v_1__62_ | v_1__60_;
  assign addr_2__60_ = 1'b0 | 1'b0;
  assign v_3__0_ = v_2__4_ | v_2__0_;
  assign addr_3__1_ = v_1__2_ | v_1__6_;
  assign addr_3__0_ = addr_2__0_ | addr_2__4_;
  assign v_3__8_ = v_2__12_ | v_2__8_;
  assign addr_3__9_ = v_1__10_ | v_1__14_;
  assign addr_3__8_ = addr_2__8_ | addr_2__12_;
  assign v_3__16_ = v_2__20_ | v_2__16_;
  assign addr_3__17_ = v_1__18_ | v_1__22_;
  assign addr_3__16_ = addr_2__16_ | addr_2__20_;
  assign v_3__24_ = v_2__28_ | v_2__24_;
  assign addr_3__25_ = v_1__26_ | v_1__30_;
  assign addr_3__24_ = addr_2__24_ | addr_2__28_;
  assign v_3__32_ = v_2__36_ | v_2__32_;
  assign addr_3__33_ = v_1__34_ | v_1__38_;
  assign addr_3__32_ = addr_2__32_ | addr_2__36_;
  assign v_3__40_ = v_2__44_ | v_2__40_;
  assign addr_3__41_ = v_1__42_ | v_1__46_;
  assign addr_3__40_ = addr_2__40_ | addr_2__44_;
  assign v_3__48_ = v_2__52_ | v_2__48_;
  assign addr_3__49_ = v_1__50_ | v_1__54_;
  assign addr_3__48_ = addr_2__48_ | addr_2__52_;
  assign v_3__56_ = v_2__60_ | v_2__56_;
  assign addr_3__57_ = v_1__58_ | v_1__62_;
  assign addr_3__56_ = addr_2__56_ | addr_2__60_;
  assign v_4__0_ = v_3__8_ | v_3__0_;
  assign addr_4__2_ = v_2__4_ | v_2__12_;
  assign addr_4__1_ = addr_3__1_ | addr_3__9_;
  assign addr_4__0_ = addr_3__0_ | addr_3__8_;
  assign v_4__16_ = v_3__24_ | v_3__16_;
  assign addr_4__18_ = v_2__20_ | v_2__28_;
  assign addr_4__17_ = addr_3__17_ | addr_3__25_;
  assign addr_4__16_ = addr_3__16_ | addr_3__24_;
  assign v_4__32_ = v_3__40_ | v_3__32_;
  assign addr_4__34_ = v_2__36_ | v_2__44_;
  assign addr_4__33_ = addr_3__33_ | addr_3__41_;
  assign addr_4__32_ = addr_3__32_ | addr_3__40_;
  assign v_4__48_ = v_3__56_ | v_3__48_;
  assign addr_4__50_ = v_2__52_ | v_2__60_;
  assign addr_4__49_ = addr_3__49_ | addr_3__57_;
  assign addr_4__48_ = addr_3__48_ | addr_3__56_;
  assign v_5__0_ = v_4__16_ | v_4__0_;
  assign addr_5__3_ = v_3__8_ | v_3__24_;
  assign addr_5__2_ = addr_4__2_ | addr_4__18_;
  assign addr_5__1_ = addr_4__1_ | addr_4__17_;
  assign addr_5__0_ = addr_4__0_ | addr_4__16_;
  assign addr_o[5] = v_4__48_ | v_4__32_;
  assign addr_5__35_ = v_3__40_ | v_3__56_;
  assign addr_5__34_ = addr_4__34_ | addr_4__50_;
  assign addr_5__33_ = addr_4__33_ | addr_4__49_;
  assign addr_5__32_ = addr_4__32_ | addr_4__48_;
  assign v_o = addr_o[5] | v_5__0_;
  assign addr_o[4] = v_4__16_ | v_4__48_;
  assign addr_o[3] = addr_5__3_ | addr_5__35_;
  assign addr_o[2] = addr_5__2_ | addr_5__34_;
  assign addr_o[1] = addr_5__1_ | addr_5__33_;
  assign addr_o[0] = addr_5__0_ | addr_5__32_;

endmodule



module bsg_priority_encode_width_p53_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [52:0] i;
  output [5:0] addr_o;
  output v_o;
  wire [5:0] addr_o;
  wire v_o;
  wire [52:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p53_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_width_p53_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o)
  );


endmodule



module bsg_counting_leading_zeros_width_p52
(
  a_i,
  num_zero_o
);

  input [51:0] a_i;
  output [5:0] num_zero_o;
  wire [5:0] num_zero_o;

  bsg_priority_encode_width_p53_lo_to_hi_p1
  pe0
  (
    .i({ 1'b1, a_i[0:0], a_i[1:1], a_i[2:2], a_i[3:3], a_i[4:4], a_i[5:5], a_i[6:6], a_i[7:7], a_i[8:8], a_i[9:9], a_i[10:10], a_i[11:11], a_i[12:12], a_i[13:13], a_i[14:14], a_i[15:15], a_i[16:16], a_i[17:17], a_i[18:18], a_i[19:19], a_i[20:20], a_i[21:21], a_i[22:22], a_i[23:23], a_i[24:24], a_i[25:25], a_i[26:26], a_i[27:27], a_i[28:28], a_i[29:29], a_i[30:30], a_i[31:31], a_i[32:32], a_i[33:33], a_i[34:34], a_i[35:35], a_i[36:36], a_i[37:37], a_i[38:38], a_i[39:39], a_i[40:40], a_i[41:41], a_i[42:42], a_i[43:43], a_i[44:44], a_i[45:45], a_i[46:46], a_i[47:47], a_i[48:48], a_i[49:49], a_i[50:50], a_i[51:51] }),
    .addr_o(num_zero_o)
  );


endmodule



module fNToRecFN_expWidth11_sigWidth53
(
  in,
  out
);

  input [63:0] in;
  output [64:0] out;
  wire [64:0] out;
  wire N0,N1,N2,out_64_,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  isZero,isSpecial,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,
  N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,
  N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,
  N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86;
  wire [5:0] normDist;
  wire [51:1] subnormFract;
  wire [11:9] adjustedExp;
  assign out_64_ = in[63];
  assign out[64] = out_64_;

  bsg_counting_leading_zeros_width_p52
  clz
  (
    .a_i(in[51:0]),
    .num_zero_o(normDist)
  );

  assign isSpecial = adjustedExp[11:10] == { 1'b1, 1'b1 };
  assign subnormFract = in[50:0] << normDist;
  assign N24 = in[50] | in[51];
  assign N25 = in[49] | N24;
  assign N26 = in[48] | N25;
  assign N27 = in[47] | N26;
  assign N28 = in[46] | N27;
  assign N29 = in[45] | N28;
  assign N30 = in[44] | N29;
  assign N31 = in[43] | N30;
  assign N32 = in[42] | N31;
  assign N33 = in[41] | N32;
  assign N34 = in[40] | N33;
  assign N35 = in[39] | N34;
  assign N36 = in[38] | N35;
  assign N37 = in[37] | N36;
  assign N38 = in[36] | N37;
  assign N39 = in[35] | N38;
  assign N40 = in[34] | N39;
  assign N41 = in[33] | N40;
  assign N42 = in[32] | N41;
  assign N43 = in[31] | N42;
  assign N44 = in[30] | N43;
  assign N45 = in[29] | N44;
  assign N46 = in[28] | N45;
  assign N47 = in[27] | N46;
  assign N48 = in[26] | N47;
  assign N49 = in[25] | N48;
  assign N50 = in[24] | N49;
  assign N51 = in[23] | N50;
  assign N52 = in[22] | N51;
  assign N53 = in[21] | N52;
  assign N54 = in[20] | N53;
  assign N55 = in[19] | N54;
  assign N56 = in[18] | N55;
  assign N57 = in[17] | N56;
  assign N58 = in[16] | N57;
  assign N59 = in[15] | N58;
  assign N60 = in[14] | N59;
  assign N61 = in[13] | N60;
  assign N62 = in[12] | N61;
  assign N63 = in[11] | N62;
  assign N64 = in[10] | N63;
  assign N65 = in[9] | N64;
  assign N66 = in[8] | N65;
  assign N67 = in[7] | N66;
  assign N68 = in[6] | N67;
  assign N69 = in[5] | N68;
  assign N70 = in[4] | N69;
  assign N71 = in[3] | N70;
  assign N72 = in[2] | N71;
  assign N73 = in[1] | N72;
  assign N74 = in[0] | N73;
  assign N75 = ~N74;
  assign N76 = in[61] | in[62];
  assign N77 = in[60] | N76;
  assign N78 = in[59] | N77;
  assign N79 = in[58] | N78;
  assign N80 = in[57] | N79;
  assign N81 = in[56] | N80;
  assign N82 = in[55] | N81;
  assign N83 = in[54] | N82;
  assign N84 = in[53] | N83;
  assign N85 = in[52] | N84;
  assign N86 = ~N85;
  assign { adjustedExp, out[60:52] } = { N86, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9 } + { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N86, N85 };
  assign { N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9 } = (N0)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, N3, N4, N5, N6, N7, N8 } : 
                                                                    (N1)? in[62:52] : 1'b0;
  assign N0 = N86;
  assign N1 = N85;
  assign out[63:61] = (N2)? { 1'b1, 1'b1, N74 } : 
                      (N23)? { 1'b0, 1'b0, 1'b0 } : 
                      (N21)? adjustedExp : 1'b0;
  assign N2 = isSpecial;
  assign out[51:0] = (N0)? { subnormFract, 1'b0 } : 
                     (N1)? in[51:0] : 1'b0;
  assign N3 = ~normDist[5];
  assign N4 = ~normDist[4];
  assign N5 = ~normDist[3];
  assign N6 = ~normDist[2];
  assign N7 = ~normDist[1];
  assign N8 = ~normDist[0];
  assign isZero = N86 & N75;
  assign N20 = isZero | isSpecial;
  assign N21 = ~N20;
  assign N22 = ~isSpecial;
  assign N23 = isZero & N22;

endmodule



module bp_be_fp_box_00
(
  ieee_i,
  tag_i,
  reg_o
);

  input [63:0] ieee_i;
  input [0:0] tag_i;
  output [65:0] reg_o;
  wire [65:0] reg_o;
  wire N0,N1,N2,N3,N4,special,N5,sp2dp_rec_exp__11_,sp2dp_rec_exp__10_,
  sp2dp_rec_exp__9_,nanbox_v_li,encode_as_sp,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39;
  wire [32:0] in_sp_rec_li;
  wire [64:0] in_dp_rec_li;
  wire [11:0] adjusted_exp;

  fNToRecFN_expWidth8_sigWidth24
  in32_rec
  (
    .in(ieee_i[31:0]),
    .out(in_sp_rec_li)
  );


  fNToRecFN_expWidth11_sigWidth53
  in64_rec
  (
    .in(ieee_i),
    .out(in_dp_rec_li)
  );

  assign N4 = in_sp_rec_li[31:29] >= { 1'b1, 1'b1, 1'b0 };
  assign N7 = in_sp_rec_li[30] | in_sp_rec_li[31];
  assign N8 = in_sp_rec_li[29] | N7;
  assign N9 = ~N8;
  assign adjusted_exp = in_sp_rec_li[31:23] + { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign { sp2dp_rec_exp__11_, sp2dp_rec_exp__10_, sp2dp_rec_exp__9_ } = (N0)? in_sp_rec_li[31:29] : 
                                                                         (N1)? adjusted_exp[11:9] : 1'b0;
  assign N0 = special;
  assign N1 = N5;
  assign reg_o[64:0] = (N2)? { in_sp_rec_li[32:32], sp2dp_rec_exp__11_, sp2dp_rec_exp__10_, sp2dp_rec_exp__9_, adjusted_exp[8:0], in_sp_rec_li[22:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N3)? in_dp_rec_li : 1'b0;
  assign N2 = reg_o[65];
  assign N3 = N6;
  assign special = N9 | N4;
  assign N5 = ~special;
  assign nanbox_v_li = N39 & ieee_i[32];
  assign N39 = N38 & ieee_i[33];
  assign N38 = N37 & ieee_i[34];
  assign N37 = N36 & ieee_i[35];
  assign N36 = N35 & ieee_i[36];
  assign N35 = N34 & ieee_i[37];
  assign N34 = N33 & ieee_i[38];
  assign N33 = N32 & ieee_i[39];
  assign N32 = N31 & ieee_i[40];
  assign N31 = N30 & ieee_i[41];
  assign N30 = N29 & ieee_i[42];
  assign N29 = N28 & ieee_i[43];
  assign N28 = N27 & ieee_i[44];
  assign N27 = N26 & ieee_i[45];
  assign N26 = N25 & ieee_i[46];
  assign N25 = N24 & ieee_i[47];
  assign N24 = N23 & ieee_i[48];
  assign N23 = N22 & ieee_i[49];
  assign N22 = N21 & ieee_i[50];
  assign N21 = N20 & ieee_i[51];
  assign N20 = N19 & ieee_i[52];
  assign N19 = N18 & ieee_i[53];
  assign N18 = N17 & ieee_i[54];
  assign N17 = N16 & ieee_i[55];
  assign N16 = N15 & ieee_i[56];
  assign N15 = N14 & ieee_i[57];
  assign N14 = N13 & ieee_i[58];
  assign N13 = N12 & ieee_i[59];
  assign N12 = N11 & ieee_i[60];
  assign N11 = N10 & ieee_i[61];
  assign N10 = ieee_i[63] & ieee_i[62];
  assign encode_as_sp = nanbox_v_li | tag_i[0];
  assign N6 = ~encode_as_sp;
  assign reg_o[65] = encode_as_sp;

endmodule



module reverse_width54
(
  in,
  out
);

  input [53:0] in;
  output [53:0] out;
  wire [53:0] out;
  assign out[53] = in[0];
  assign out[52] = in[1];
  assign out[51] = in[2];
  assign out[50] = in[3];
  assign out[49] = in[4];
  assign out[48] = in[5];
  assign out[47] = in[6];
  assign out[46] = in[7];
  assign out[45] = in[8];
  assign out[44] = in[9];
  assign out[43] = in[10];
  assign out[42] = in[11];
  assign out[41] = in[12];
  assign out[40] = in[13];
  assign out[39] = in[14];
  assign out[38] = in[15];
  assign out[37] = in[16];
  assign out[36] = in[17];
  assign out[35] = in[18];
  assign out[34] = in[19];
  assign out[33] = in[20];
  assign out[32] = in[21];
  assign out[31] = in[22];
  assign out[30] = in[23];
  assign out[29] = in[24];
  assign out[28] = in[25];
  assign out[27] = in[26];
  assign out[26] = in[27];
  assign out[25] = in[28];
  assign out[24] = in[29];
  assign out[23] = in[30];
  assign out[22] = in[31];
  assign out[21] = in[32];
  assign out[20] = in[33];
  assign out[19] = in[34];
  assign out[18] = in[35];
  assign out[17] = in[36];
  assign out[16] = in[37];
  assign out[15] = in[38];
  assign out[14] = in[39];
  assign out[13] = in[40];
  assign out[12] = in[41];
  assign out[11] = in[42];
  assign out[10] = in[43];
  assign out[9] = in[44];
  assign out[8] = in[45];
  assign out[7] = in[46];
  assign out[6] = in[47];
  assign out[5] = in[48];
  assign out[4] = in[49];
  assign out[3] = in[50];
  assign out[2] = in[51];
  assign out[1] = in[52];
  assign out[0] = in[53];

endmodule



module lowMaskLoHi_inWidth12_topBound972_bottomBound1026
(
  in,
  out
);

  input [11:0] in;
  output [53:0] out;
  wire [53:0] out,reverseOut;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,
  sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,
  sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,
  sv2v_dc_20,sv2v_dc_21,sv2v_dc_22,sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,
  sv2v_dc_27,sv2v_dc_28,sv2v_dc_29,sv2v_dc_30,sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,
  sv2v_dc_34,sv2v_dc_35,sv2v_dc_36,sv2v_dc_37,sv2v_dc_38,sv2v_dc_39,sv2v_dc_40,sv2v_dc_41,
  sv2v_dc_42,sv2v_dc_43,sv2v_dc_44,sv2v_dc_45,sv2v_dc_46,sv2v_dc_47,sv2v_dc_48,
  sv2v_dc_49,sv2v_dc_50,sv2v_dc_51,sv2v_dc_52,sv2v_dc_53,sv2v_dc_54,sv2v_dc_55,
  sv2v_dc_56,sv2v_dc_57,sv2v_dc_58,sv2v_dc_59,sv2v_dc_60,sv2v_dc_61,sv2v_dc_62,
  sv2v_dc_63,sv2v_dc_64,sv2v_dc_65,sv2v_dc_66,sv2v_dc_67,sv2v_dc_68,sv2v_dc_69,sv2v_dc_70,
  sv2v_dc_71,sv2v_dc_72,sv2v_dc_73,sv2v_dc_74,sv2v_dc_75,sv2v_dc_76,sv2v_dc_77,
  sv2v_dc_78,sv2v_dc_79,sv2v_dc_80,sv2v_dc_81,sv2v_dc_82,sv2v_dc_83,sv2v_dc_84,
  sv2v_dc_85,sv2v_dc_86,sv2v_dc_87,sv2v_dc_88,sv2v_dc_89,sv2v_dc_90,sv2v_dc_91,
  sv2v_dc_92,sv2v_dc_93,sv2v_dc_94,sv2v_dc_95,sv2v_dc_96,sv2v_dc_97,sv2v_dc_98,sv2v_dc_99,
  sv2v_dc_100,sv2v_dc_101,sv2v_dc_102,sv2v_dc_103,sv2v_dc_104,sv2v_dc_105,
  sv2v_dc_106,sv2v_dc_107,sv2v_dc_108,sv2v_dc_109,sv2v_dc_110,sv2v_dc_111,sv2v_dc_112,
  sv2v_dc_113,sv2v_dc_114,sv2v_dc_115,sv2v_dc_116,sv2v_dc_117,sv2v_dc_118,sv2v_dc_119,
  sv2v_dc_120,sv2v_dc_121,sv2v_dc_122,sv2v_dc_123,sv2v_dc_124,sv2v_dc_125,
  sv2v_dc_126,sv2v_dc_127,sv2v_dc_128,sv2v_dc_129,sv2v_dc_130,sv2v_dc_131,sv2v_dc_132,
  sv2v_dc_133,sv2v_dc_134,sv2v_dc_135,sv2v_dc_136,sv2v_dc_137,sv2v_dc_138,sv2v_dc_139,
  sv2v_dc_140,sv2v_dc_141,sv2v_dc_142,sv2v_dc_143,sv2v_dc_144,sv2v_dc_145,
  sv2v_dc_146,sv2v_dc_147,sv2v_dc_148,sv2v_dc_149,sv2v_dc_150,sv2v_dc_151,sv2v_dc_152,
  sv2v_dc_153,sv2v_dc_154,sv2v_dc_155,sv2v_dc_156,sv2v_dc_157,sv2v_dc_158,sv2v_dc_159,
  sv2v_dc_160,sv2v_dc_161,sv2v_dc_162,sv2v_dc_163,sv2v_dc_164,sv2v_dc_165,
  sv2v_dc_166,sv2v_dc_167,sv2v_dc_168,sv2v_dc_169,sv2v_dc_170,sv2v_dc_171,sv2v_dc_172,
  sv2v_dc_173,sv2v_dc_174,sv2v_dc_175,sv2v_dc_176,sv2v_dc_177,sv2v_dc_178,sv2v_dc_179,
  sv2v_dc_180,sv2v_dc_181,sv2v_dc_182,sv2v_dc_183,sv2v_dc_184,sv2v_dc_185,
  sv2v_dc_186,sv2v_dc_187,sv2v_dc_188,sv2v_dc_189,sv2v_dc_190,sv2v_dc_191,sv2v_dc_192,
  sv2v_dc_193,sv2v_dc_194,sv2v_dc_195,sv2v_dc_196,sv2v_dc_197,sv2v_dc_198,sv2v_dc_199,
  sv2v_dc_200,sv2v_dc_201,sv2v_dc_202,sv2v_dc_203,sv2v_dc_204,sv2v_dc_205,
  sv2v_dc_206,sv2v_dc_207,sv2v_dc_208,sv2v_dc_209,sv2v_dc_210,sv2v_dc_211,sv2v_dc_212,
  sv2v_dc_213,sv2v_dc_214,sv2v_dc_215,sv2v_dc_216,sv2v_dc_217,sv2v_dc_218,sv2v_dc_219,
  sv2v_dc_220,sv2v_dc_221,sv2v_dc_222,sv2v_dc_223,sv2v_dc_224,sv2v_dc_225,
  sv2v_dc_226,sv2v_dc_227,sv2v_dc_228,sv2v_dc_229,sv2v_dc_230,sv2v_dc_231,sv2v_dc_232,
  sv2v_dc_233,sv2v_dc_234,sv2v_dc_235,sv2v_dc_236,sv2v_dc_237,sv2v_dc_238,sv2v_dc_239,
  sv2v_dc_240,sv2v_dc_241,sv2v_dc_242,sv2v_dc_243,sv2v_dc_244,sv2v_dc_245,
  sv2v_dc_246,sv2v_dc_247,sv2v_dc_248,sv2v_dc_249,sv2v_dc_250,sv2v_dc_251,sv2v_dc_252,
  sv2v_dc_253,sv2v_dc_254,sv2v_dc_255,sv2v_dc_256,sv2v_dc_257,sv2v_dc_258,sv2v_dc_259,
  sv2v_dc_260,sv2v_dc_261,sv2v_dc_262,sv2v_dc_263,sv2v_dc_264,sv2v_dc_265,
  sv2v_dc_266,sv2v_dc_267,sv2v_dc_268,sv2v_dc_269,sv2v_dc_270,sv2v_dc_271,sv2v_dc_272,
  sv2v_dc_273,sv2v_dc_274,sv2v_dc_275,sv2v_dc_276,sv2v_dc_277,sv2v_dc_278,sv2v_dc_279,
  sv2v_dc_280,sv2v_dc_281,sv2v_dc_282,sv2v_dc_283,sv2v_dc_284,sv2v_dc_285,
  sv2v_dc_286,sv2v_dc_287,sv2v_dc_288,sv2v_dc_289,sv2v_dc_290,sv2v_dc_291,sv2v_dc_292,
  sv2v_dc_293,sv2v_dc_294,sv2v_dc_295,sv2v_dc_296,sv2v_dc_297,sv2v_dc_298,sv2v_dc_299,
  sv2v_dc_300,sv2v_dc_301,sv2v_dc_302,sv2v_dc_303,sv2v_dc_304,sv2v_dc_305,
  sv2v_dc_306,sv2v_dc_307,sv2v_dc_308,sv2v_dc_309,sv2v_dc_310,sv2v_dc_311,sv2v_dc_312,
  sv2v_dc_313,sv2v_dc_314,sv2v_dc_315,sv2v_dc_316,sv2v_dc_317,sv2v_dc_318,sv2v_dc_319,
  sv2v_dc_320,sv2v_dc_321,sv2v_dc_322,sv2v_dc_323,sv2v_dc_324,sv2v_dc_325,
  sv2v_dc_326,sv2v_dc_327,sv2v_dc_328,sv2v_dc_329,sv2v_dc_330,sv2v_dc_331,sv2v_dc_332,
  sv2v_dc_333,sv2v_dc_334,sv2v_dc_335,sv2v_dc_336,sv2v_dc_337,sv2v_dc_338,sv2v_dc_339,
  sv2v_dc_340,sv2v_dc_341,sv2v_dc_342,sv2v_dc_343,sv2v_dc_344,sv2v_dc_345,
  sv2v_dc_346,sv2v_dc_347,sv2v_dc_348,sv2v_dc_349,sv2v_dc_350,sv2v_dc_351,sv2v_dc_352,
  sv2v_dc_353,sv2v_dc_354,sv2v_dc_355,sv2v_dc_356,sv2v_dc_357,sv2v_dc_358,sv2v_dc_359,
  sv2v_dc_360,sv2v_dc_361,sv2v_dc_362,sv2v_dc_363,sv2v_dc_364,sv2v_dc_365,
  sv2v_dc_366,sv2v_dc_367,sv2v_dc_368,sv2v_dc_369,sv2v_dc_370,sv2v_dc_371,sv2v_dc_372,
  sv2v_dc_373,sv2v_dc_374,sv2v_dc_375,sv2v_dc_376,sv2v_dc_377,sv2v_dc_378,sv2v_dc_379,
  sv2v_dc_380,sv2v_dc_381,sv2v_dc_382,sv2v_dc_383,sv2v_dc_384,sv2v_dc_385,
  sv2v_dc_386,sv2v_dc_387,sv2v_dc_388,sv2v_dc_389,sv2v_dc_390,sv2v_dc_391,sv2v_dc_392,
  sv2v_dc_393,sv2v_dc_394,sv2v_dc_395,sv2v_dc_396,sv2v_dc_397,sv2v_dc_398,sv2v_dc_399,
  sv2v_dc_400,sv2v_dc_401,sv2v_dc_402,sv2v_dc_403,sv2v_dc_404,sv2v_dc_405,
  sv2v_dc_406,sv2v_dc_407,sv2v_dc_408,sv2v_dc_409,sv2v_dc_410,sv2v_dc_411,sv2v_dc_412,
  sv2v_dc_413,sv2v_dc_414,sv2v_dc_415,sv2v_dc_416,sv2v_dc_417,sv2v_dc_418,sv2v_dc_419,
  sv2v_dc_420,sv2v_dc_421,sv2v_dc_422,sv2v_dc_423,sv2v_dc_424,sv2v_dc_425,
  sv2v_dc_426,sv2v_dc_427,sv2v_dc_428,sv2v_dc_429,sv2v_dc_430,sv2v_dc_431,sv2v_dc_432,
  sv2v_dc_433,sv2v_dc_434,sv2v_dc_435,sv2v_dc_436,sv2v_dc_437,sv2v_dc_438,sv2v_dc_439,
  sv2v_dc_440,sv2v_dc_441,sv2v_dc_442,sv2v_dc_443,sv2v_dc_444,sv2v_dc_445,
  sv2v_dc_446,sv2v_dc_447,sv2v_dc_448,sv2v_dc_449,sv2v_dc_450,sv2v_dc_451,sv2v_dc_452,
  sv2v_dc_453,sv2v_dc_454,sv2v_dc_455,sv2v_dc_456,sv2v_dc_457,sv2v_dc_458,sv2v_dc_459,
  sv2v_dc_460,sv2v_dc_461,sv2v_dc_462,sv2v_dc_463,sv2v_dc_464,sv2v_dc_465,
  sv2v_dc_466,sv2v_dc_467,sv2v_dc_468,sv2v_dc_469,sv2v_dc_470,sv2v_dc_471,sv2v_dc_472,
  sv2v_dc_473,sv2v_dc_474,sv2v_dc_475,sv2v_dc_476,sv2v_dc_477,sv2v_dc_478,sv2v_dc_479,
  sv2v_dc_480,sv2v_dc_481,sv2v_dc_482,sv2v_dc_483,sv2v_dc_484,sv2v_dc_485,
  sv2v_dc_486,sv2v_dc_487,sv2v_dc_488,sv2v_dc_489,sv2v_dc_490,sv2v_dc_491,sv2v_dc_492,
  sv2v_dc_493,sv2v_dc_494,sv2v_dc_495,sv2v_dc_496,sv2v_dc_497,sv2v_dc_498,sv2v_dc_499,
  sv2v_dc_500,sv2v_dc_501,sv2v_dc_502,sv2v_dc_503,sv2v_dc_504,sv2v_dc_505,
  sv2v_dc_506,sv2v_dc_507,sv2v_dc_508,sv2v_dc_509,sv2v_dc_510,sv2v_dc_511,sv2v_dc_512,
  sv2v_dc_513,sv2v_dc_514,sv2v_dc_515,sv2v_dc_516,sv2v_dc_517,sv2v_dc_518,sv2v_dc_519,
  sv2v_dc_520,sv2v_dc_521,sv2v_dc_522,sv2v_dc_523,sv2v_dc_524,sv2v_dc_525,
  sv2v_dc_526,sv2v_dc_527,sv2v_dc_528,sv2v_dc_529,sv2v_dc_530,sv2v_dc_531,sv2v_dc_532,
  sv2v_dc_533,sv2v_dc_534,sv2v_dc_535,sv2v_dc_536,sv2v_dc_537,sv2v_dc_538,sv2v_dc_539,
  sv2v_dc_540,sv2v_dc_541,sv2v_dc_542,sv2v_dc_543,sv2v_dc_544,sv2v_dc_545,
  sv2v_dc_546,sv2v_dc_547,sv2v_dc_548,sv2v_dc_549,sv2v_dc_550,sv2v_dc_551,sv2v_dc_552,
  sv2v_dc_553,sv2v_dc_554,sv2v_dc_555,sv2v_dc_556,sv2v_dc_557,sv2v_dc_558,sv2v_dc_559,
  sv2v_dc_560,sv2v_dc_561,sv2v_dc_562,sv2v_dc_563,sv2v_dc_564,sv2v_dc_565,
  sv2v_dc_566,sv2v_dc_567,sv2v_dc_568,sv2v_dc_569,sv2v_dc_570,sv2v_dc_571,sv2v_dc_572,
  sv2v_dc_573,sv2v_dc_574,sv2v_dc_575,sv2v_dc_576,sv2v_dc_577,sv2v_dc_578,sv2v_dc_579,
  sv2v_dc_580,sv2v_dc_581,sv2v_dc_582,sv2v_dc_583,sv2v_dc_584,sv2v_dc_585,
  sv2v_dc_586,sv2v_dc_587,sv2v_dc_588,sv2v_dc_589,sv2v_dc_590,sv2v_dc_591,sv2v_dc_592,
  sv2v_dc_593,sv2v_dc_594,sv2v_dc_595,sv2v_dc_596,sv2v_dc_597,sv2v_dc_598,sv2v_dc_599,
  sv2v_dc_600,sv2v_dc_601,sv2v_dc_602,sv2v_dc_603,sv2v_dc_604,sv2v_dc_605,
  sv2v_dc_606,sv2v_dc_607,sv2v_dc_608,sv2v_dc_609,sv2v_dc_610,sv2v_dc_611,sv2v_dc_612,
  sv2v_dc_613,sv2v_dc_614,sv2v_dc_615,sv2v_dc_616,sv2v_dc_617,sv2v_dc_618,sv2v_dc_619,
  sv2v_dc_620,sv2v_dc_621,sv2v_dc_622,sv2v_dc_623,sv2v_dc_624,sv2v_dc_625,
  sv2v_dc_626,sv2v_dc_627,sv2v_dc_628,sv2v_dc_629,sv2v_dc_630,sv2v_dc_631,sv2v_dc_632,
  sv2v_dc_633,sv2v_dc_634,sv2v_dc_635,sv2v_dc_636,sv2v_dc_637,sv2v_dc_638,sv2v_dc_639,
  sv2v_dc_640,sv2v_dc_641,sv2v_dc_642,sv2v_dc_643,sv2v_dc_644,sv2v_dc_645,
  sv2v_dc_646,sv2v_dc_647,sv2v_dc_648,sv2v_dc_649,sv2v_dc_650,sv2v_dc_651,sv2v_dc_652,
  sv2v_dc_653,sv2v_dc_654,sv2v_dc_655,sv2v_dc_656,sv2v_dc_657,sv2v_dc_658,sv2v_dc_659,
  sv2v_dc_660,sv2v_dc_661,sv2v_dc_662,sv2v_dc_663,sv2v_dc_664,sv2v_dc_665,
  sv2v_dc_666,sv2v_dc_667,sv2v_dc_668,sv2v_dc_669,sv2v_dc_670,sv2v_dc_671,sv2v_dc_672,
  sv2v_dc_673,sv2v_dc_674,sv2v_dc_675,sv2v_dc_676,sv2v_dc_677,sv2v_dc_678,sv2v_dc_679,
  sv2v_dc_680,sv2v_dc_681,sv2v_dc_682,sv2v_dc_683,sv2v_dc_684,sv2v_dc_685,
  sv2v_dc_686,sv2v_dc_687,sv2v_dc_688,sv2v_dc_689,sv2v_dc_690,sv2v_dc_691,sv2v_dc_692,
  sv2v_dc_693,sv2v_dc_694,sv2v_dc_695,sv2v_dc_696,sv2v_dc_697,sv2v_dc_698,sv2v_dc_699,
  sv2v_dc_700,sv2v_dc_701,sv2v_dc_702,sv2v_dc_703,sv2v_dc_704,sv2v_dc_705,
  sv2v_dc_706,sv2v_dc_707,sv2v_dc_708,sv2v_dc_709,sv2v_dc_710,sv2v_dc_711,sv2v_dc_712,
  sv2v_dc_713,sv2v_dc_714,sv2v_dc_715,sv2v_dc_716,sv2v_dc_717,sv2v_dc_718,sv2v_dc_719,
  sv2v_dc_720,sv2v_dc_721,sv2v_dc_722,sv2v_dc_723,sv2v_dc_724,sv2v_dc_725,
  sv2v_dc_726,sv2v_dc_727,sv2v_dc_728,sv2v_dc_729,sv2v_dc_730,sv2v_dc_731,sv2v_dc_732,
  sv2v_dc_733,sv2v_dc_734,sv2v_dc_735,sv2v_dc_736,sv2v_dc_737,sv2v_dc_738,sv2v_dc_739,
  sv2v_dc_740,sv2v_dc_741,sv2v_dc_742,sv2v_dc_743,sv2v_dc_744,sv2v_dc_745,
  sv2v_dc_746,sv2v_dc_747,sv2v_dc_748,sv2v_dc_749,sv2v_dc_750,sv2v_dc_751,sv2v_dc_752,
  sv2v_dc_753,sv2v_dc_754,sv2v_dc_755,sv2v_dc_756,sv2v_dc_757,sv2v_dc_758,sv2v_dc_759,
  sv2v_dc_760,sv2v_dc_761,sv2v_dc_762,sv2v_dc_763,sv2v_dc_764,sv2v_dc_765,
  sv2v_dc_766,sv2v_dc_767,sv2v_dc_768,sv2v_dc_769,sv2v_dc_770,sv2v_dc_771,sv2v_dc_772,
  sv2v_dc_773,sv2v_dc_774,sv2v_dc_775,sv2v_dc_776,sv2v_dc_777,sv2v_dc_778,sv2v_dc_779,
  sv2v_dc_780,sv2v_dc_781,sv2v_dc_782,sv2v_dc_783,sv2v_dc_784,sv2v_dc_785,
  sv2v_dc_786,sv2v_dc_787,sv2v_dc_788,sv2v_dc_789,sv2v_dc_790,sv2v_dc_791,sv2v_dc_792,
  sv2v_dc_793,sv2v_dc_794,sv2v_dc_795,sv2v_dc_796,sv2v_dc_797,sv2v_dc_798,sv2v_dc_799,
  sv2v_dc_800,sv2v_dc_801,sv2v_dc_802,sv2v_dc_803,sv2v_dc_804,sv2v_dc_805,
  sv2v_dc_806,sv2v_dc_807,sv2v_dc_808,sv2v_dc_809,sv2v_dc_810,sv2v_dc_811,sv2v_dc_812,
  sv2v_dc_813,sv2v_dc_814,sv2v_dc_815,sv2v_dc_816,sv2v_dc_817,sv2v_dc_818,sv2v_dc_819,
  sv2v_dc_820,sv2v_dc_821,sv2v_dc_822,sv2v_dc_823,sv2v_dc_824,sv2v_dc_825,
  sv2v_dc_826,sv2v_dc_827,sv2v_dc_828,sv2v_dc_829,sv2v_dc_830,sv2v_dc_831,sv2v_dc_832,
  sv2v_dc_833,sv2v_dc_834,sv2v_dc_835,sv2v_dc_836,sv2v_dc_837,sv2v_dc_838,sv2v_dc_839,
  sv2v_dc_840,sv2v_dc_841,sv2v_dc_842,sv2v_dc_843,sv2v_dc_844,sv2v_dc_845,
  sv2v_dc_846,sv2v_dc_847,sv2v_dc_848,sv2v_dc_849,sv2v_dc_850,sv2v_dc_851,sv2v_dc_852,
  sv2v_dc_853,sv2v_dc_854,sv2v_dc_855,sv2v_dc_856,sv2v_dc_857,sv2v_dc_858,sv2v_dc_859,
  sv2v_dc_860,sv2v_dc_861,sv2v_dc_862,sv2v_dc_863,sv2v_dc_864,sv2v_dc_865,
  sv2v_dc_866,sv2v_dc_867,sv2v_dc_868,sv2v_dc_869,sv2v_dc_870,sv2v_dc_871,sv2v_dc_872,
  sv2v_dc_873,sv2v_dc_874,sv2v_dc_875,sv2v_dc_876,sv2v_dc_877,sv2v_dc_878,sv2v_dc_879,
  sv2v_dc_880,sv2v_dc_881,sv2v_dc_882,sv2v_dc_883,sv2v_dc_884,sv2v_dc_885,
  sv2v_dc_886,sv2v_dc_887,sv2v_dc_888,sv2v_dc_889,sv2v_dc_890,sv2v_dc_891,sv2v_dc_892,
  sv2v_dc_893,sv2v_dc_894,sv2v_dc_895,sv2v_dc_896,sv2v_dc_897,sv2v_dc_898,sv2v_dc_899,
  sv2v_dc_900,sv2v_dc_901,sv2v_dc_902,sv2v_dc_903,sv2v_dc_904,sv2v_dc_905,
  sv2v_dc_906,sv2v_dc_907,sv2v_dc_908,sv2v_dc_909,sv2v_dc_910,sv2v_dc_911,sv2v_dc_912,
  sv2v_dc_913,sv2v_dc_914,sv2v_dc_915,sv2v_dc_916,sv2v_dc_917,sv2v_dc_918,sv2v_dc_919,
  sv2v_dc_920,sv2v_dc_921,sv2v_dc_922,sv2v_dc_923,sv2v_dc_924,sv2v_dc_925,
  sv2v_dc_926,sv2v_dc_927,sv2v_dc_928,sv2v_dc_929,sv2v_dc_930,sv2v_dc_931,sv2v_dc_932,
  sv2v_dc_933,sv2v_dc_934,sv2v_dc_935,sv2v_dc_936,sv2v_dc_937,sv2v_dc_938,sv2v_dc_939,
  sv2v_dc_940,sv2v_dc_941,sv2v_dc_942,sv2v_dc_943,sv2v_dc_944,sv2v_dc_945,
  sv2v_dc_946,sv2v_dc_947,sv2v_dc_948,sv2v_dc_949,sv2v_dc_950,sv2v_dc_951,sv2v_dc_952,
  sv2v_dc_953,sv2v_dc_954,sv2v_dc_955,sv2v_dc_956,sv2v_dc_957,sv2v_dc_958,sv2v_dc_959,
  sv2v_dc_960,sv2v_dc_961,sv2v_dc_962,sv2v_dc_963,sv2v_dc_964,sv2v_dc_965,
  sv2v_dc_966,sv2v_dc_967,sv2v_dc_968,sv2v_dc_969,sv2v_dc_970,sv2v_dc_971,sv2v_dc_972,
  sv2v_dc_973,sv2v_dc_974,sv2v_dc_975,sv2v_dc_976,sv2v_dc_977,sv2v_dc_978,sv2v_dc_979,
  sv2v_dc_980,sv2v_dc_981,sv2v_dc_982,sv2v_dc_983,sv2v_dc_984,sv2v_dc_985,
  sv2v_dc_986,sv2v_dc_987,sv2v_dc_988,sv2v_dc_989,sv2v_dc_990,sv2v_dc_991,sv2v_dc_992,
  sv2v_dc_993,sv2v_dc_994,sv2v_dc_995,sv2v_dc_996,sv2v_dc_997,sv2v_dc_998,sv2v_dc_999,
  sv2v_dc_1000,sv2v_dc_1001,sv2v_dc_1002,sv2v_dc_1003,sv2v_dc_1004,sv2v_dc_1005,
  sv2v_dc_1006,sv2v_dc_1007,sv2v_dc_1008,sv2v_dc_1009,sv2v_dc_1010,sv2v_dc_1011,
  sv2v_dc_1012,sv2v_dc_1013,sv2v_dc_1014,sv2v_dc_1015,sv2v_dc_1016,sv2v_dc_1017,
  sv2v_dc_1018,sv2v_dc_1019,sv2v_dc_1020,sv2v_dc_1021,sv2v_dc_1022,sv2v_dc_1023,
  sv2v_dc_1024,sv2v_dc_1025,sv2v_dc_1026,sv2v_dc_1027,sv2v_dc_1028,sv2v_dc_1029,
  sv2v_dc_1030,sv2v_dc_1031,sv2v_dc_1032,sv2v_dc_1033,sv2v_dc_1034,sv2v_dc_1035,sv2v_dc_1036,
  sv2v_dc_1037,sv2v_dc_1038,sv2v_dc_1039,sv2v_dc_1040,sv2v_dc_1041,sv2v_dc_1042,
  sv2v_dc_1043,sv2v_dc_1044,sv2v_dc_1045,sv2v_dc_1046,sv2v_dc_1047,sv2v_dc_1048,
  sv2v_dc_1049,sv2v_dc_1050,sv2v_dc_1051,sv2v_dc_1052,sv2v_dc_1053,sv2v_dc_1054,
  sv2v_dc_1055,sv2v_dc_1056,sv2v_dc_1057,sv2v_dc_1058,sv2v_dc_1059,sv2v_dc_1060,
  sv2v_dc_1061,sv2v_dc_1062,sv2v_dc_1063,sv2v_dc_1064,sv2v_dc_1065,sv2v_dc_1066,
  sv2v_dc_1067,sv2v_dc_1068,sv2v_dc_1069,sv2v_dc_1070,sv2v_dc_1071,sv2v_dc_1072,sv2v_dc_1073,
  sv2v_dc_1074,sv2v_dc_1075,sv2v_dc_1076,sv2v_dc_1077,sv2v_dc_1078,sv2v_dc_1079,
  sv2v_dc_1080,sv2v_dc_1081,sv2v_dc_1082,sv2v_dc_1083,sv2v_dc_1084,sv2v_dc_1085,
  sv2v_dc_1086,sv2v_dc_1087,sv2v_dc_1088,sv2v_dc_1089,sv2v_dc_1090,sv2v_dc_1091,
  sv2v_dc_1092,sv2v_dc_1093,sv2v_dc_1094,sv2v_dc_1095,sv2v_dc_1096,sv2v_dc_1097,
  sv2v_dc_1098,sv2v_dc_1099,sv2v_dc_1100,sv2v_dc_1101,sv2v_dc_1102,sv2v_dc_1103,
  sv2v_dc_1104,sv2v_dc_1105,sv2v_dc_1106,sv2v_dc_1107,sv2v_dc_1108,sv2v_dc_1109,
  sv2v_dc_1110,sv2v_dc_1111,sv2v_dc_1112,sv2v_dc_1113,sv2v_dc_1114,sv2v_dc_1115,sv2v_dc_1116,
  sv2v_dc_1117,sv2v_dc_1118,sv2v_dc_1119,sv2v_dc_1120,sv2v_dc_1121,sv2v_dc_1122,
  sv2v_dc_1123,sv2v_dc_1124,sv2v_dc_1125,sv2v_dc_1126,sv2v_dc_1127,sv2v_dc_1128,
  sv2v_dc_1129,sv2v_dc_1130,sv2v_dc_1131,sv2v_dc_1132,sv2v_dc_1133,sv2v_dc_1134,
  sv2v_dc_1135,sv2v_dc_1136,sv2v_dc_1137,sv2v_dc_1138,sv2v_dc_1139,sv2v_dc_1140,
  sv2v_dc_1141,sv2v_dc_1142,sv2v_dc_1143,sv2v_dc_1144,sv2v_dc_1145,sv2v_dc_1146,
  sv2v_dc_1147,sv2v_dc_1148,sv2v_dc_1149,sv2v_dc_1150,sv2v_dc_1151,sv2v_dc_1152,sv2v_dc_1153,
  sv2v_dc_1154,sv2v_dc_1155,sv2v_dc_1156,sv2v_dc_1157,sv2v_dc_1158,sv2v_dc_1159,
  sv2v_dc_1160,sv2v_dc_1161,sv2v_dc_1162,sv2v_dc_1163,sv2v_dc_1164,sv2v_dc_1165,
  sv2v_dc_1166,sv2v_dc_1167,sv2v_dc_1168,sv2v_dc_1169,sv2v_dc_1170,sv2v_dc_1171,
  sv2v_dc_1172,sv2v_dc_1173,sv2v_dc_1174,sv2v_dc_1175,sv2v_dc_1176,sv2v_dc_1177,
  sv2v_dc_1178,sv2v_dc_1179,sv2v_dc_1180,sv2v_dc_1181,sv2v_dc_1182,sv2v_dc_1183,
  sv2v_dc_1184,sv2v_dc_1185,sv2v_dc_1186,sv2v_dc_1187,sv2v_dc_1188,sv2v_dc_1189,
  sv2v_dc_1190,sv2v_dc_1191,sv2v_dc_1192,sv2v_dc_1193,sv2v_dc_1194,sv2v_dc_1195,sv2v_dc_1196,
  sv2v_dc_1197,sv2v_dc_1198,sv2v_dc_1199,sv2v_dc_1200,sv2v_dc_1201,sv2v_dc_1202,
  sv2v_dc_1203,sv2v_dc_1204,sv2v_dc_1205,sv2v_dc_1206,sv2v_dc_1207,sv2v_dc_1208,
  sv2v_dc_1209,sv2v_dc_1210,sv2v_dc_1211,sv2v_dc_1212,sv2v_dc_1213,sv2v_dc_1214,
  sv2v_dc_1215,sv2v_dc_1216,sv2v_dc_1217,sv2v_dc_1218,sv2v_dc_1219,sv2v_dc_1220,
  sv2v_dc_1221,sv2v_dc_1222,sv2v_dc_1223,sv2v_dc_1224,sv2v_dc_1225,sv2v_dc_1226,
  sv2v_dc_1227,sv2v_dc_1228,sv2v_dc_1229,sv2v_dc_1230,sv2v_dc_1231,sv2v_dc_1232,sv2v_dc_1233,
  sv2v_dc_1234,sv2v_dc_1235,sv2v_dc_1236,sv2v_dc_1237,sv2v_dc_1238,sv2v_dc_1239,
  sv2v_dc_1240,sv2v_dc_1241,sv2v_dc_1242,sv2v_dc_1243,sv2v_dc_1244,sv2v_dc_1245,
  sv2v_dc_1246,sv2v_dc_1247,sv2v_dc_1248,sv2v_dc_1249,sv2v_dc_1250,sv2v_dc_1251,
  sv2v_dc_1252,sv2v_dc_1253,sv2v_dc_1254,sv2v_dc_1255,sv2v_dc_1256,sv2v_dc_1257,
  sv2v_dc_1258,sv2v_dc_1259,sv2v_dc_1260,sv2v_dc_1261,sv2v_dc_1262,sv2v_dc_1263,
  sv2v_dc_1264,sv2v_dc_1265,sv2v_dc_1266,sv2v_dc_1267,sv2v_dc_1268,sv2v_dc_1269,
  sv2v_dc_1270,sv2v_dc_1271,sv2v_dc_1272,sv2v_dc_1273,sv2v_dc_1274,sv2v_dc_1275,sv2v_dc_1276,
  sv2v_dc_1277,sv2v_dc_1278,sv2v_dc_1279,sv2v_dc_1280,sv2v_dc_1281,sv2v_dc_1282,
  sv2v_dc_1283,sv2v_dc_1284,sv2v_dc_1285,sv2v_dc_1286,sv2v_dc_1287,sv2v_dc_1288,
  sv2v_dc_1289,sv2v_dc_1290,sv2v_dc_1291,sv2v_dc_1292,sv2v_dc_1293,sv2v_dc_1294,
  sv2v_dc_1295,sv2v_dc_1296,sv2v_dc_1297,sv2v_dc_1298,sv2v_dc_1299,sv2v_dc_1300,
  sv2v_dc_1301,sv2v_dc_1302,sv2v_dc_1303,sv2v_dc_1304,sv2v_dc_1305,sv2v_dc_1306,
  sv2v_dc_1307,sv2v_dc_1308,sv2v_dc_1309,sv2v_dc_1310,sv2v_dc_1311,sv2v_dc_1312,sv2v_dc_1313,
  sv2v_dc_1314,sv2v_dc_1315,sv2v_dc_1316,sv2v_dc_1317,sv2v_dc_1318,sv2v_dc_1319,
  sv2v_dc_1320,sv2v_dc_1321,sv2v_dc_1322,sv2v_dc_1323,sv2v_dc_1324,sv2v_dc_1325,
  sv2v_dc_1326,sv2v_dc_1327,sv2v_dc_1328,sv2v_dc_1329,sv2v_dc_1330,sv2v_dc_1331,
  sv2v_dc_1332,sv2v_dc_1333,sv2v_dc_1334,sv2v_dc_1335,sv2v_dc_1336,sv2v_dc_1337,
  sv2v_dc_1338,sv2v_dc_1339,sv2v_dc_1340,sv2v_dc_1341,sv2v_dc_1342,sv2v_dc_1343,
  sv2v_dc_1344,sv2v_dc_1345,sv2v_dc_1346,sv2v_dc_1347,sv2v_dc_1348,sv2v_dc_1349,
  sv2v_dc_1350,sv2v_dc_1351,sv2v_dc_1352,sv2v_dc_1353,sv2v_dc_1354,sv2v_dc_1355,sv2v_dc_1356,
  sv2v_dc_1357,sv2v_dc_1358,sv2v_dc_1359,sv2v_dc_1360,sv2v_dc_1361,sv2v_dc_1362,
  sv2v_dc_1363,sv2v_dc_1364,sv2v_dc_1365,sv2v_dc_1366,sv2v_dc_1367,sv2v_dc_1368,
  sv2v_dc_1369,sv2v_dc_1370,sv2v_dc_1371,sv2v_dc_1372,sv2v_dc_1373,sv2v_dc_1374,
  sv2v_dc_1375,sv2v_dc_1376,sv2v_dc_1377,sv2v_dc_1378,sv2v_dc_1379,sv2v_dc_1380,
  sv2v_dc_1381,sv2v_dc_1382,sv2v_dc_1383,sv2v_dc_1384,sv2v_dc_1385,sv2v_dc_1386,
  sv2v_dc_1387,sv2v_dc_1388,sv2v_dc_1389,sv2v_dc_1390,sv2v_dc_1391,sv2v_dc_1392,sv2v_dc_1393,
  sv2v_dc_1394,sv2v_dc_1395,sv2v_dc_1396,sv2v_dc_1397,sv2v_dc_1398,sv2v_dc_1399,
  sv2v_dc_1400,sv2v_dc_1401,sv2v_dc_1402,sv2v_dc_1403,sv2v_dc_1404,sv2v_dc_1405,
  sv2v_dc_1406,sv2v_dc_1407,sv2v_dc_1408,sv2v_dc_1409,sv2v_dc_1410,sv2v_dc_1411,
  sv2v_dc_1412,sv2v_dc_1413,sv2v_dc_1414,sv2v_dc_1415,sv2v_dc_1416,sv2v_dc_1417,
  sv2v_dc_1418,sv2v_dc_1419,sv2v_dc_1420,sv2v_dc_1421,sv2v_dc_1422,sv2v_dc_1423,
  sv2v_dc_1424,sv2v_dc_1425,sv2v_dc_1426,sv2v_dc_1427,sv2v_dc_1428,sv2v_dc_1429,
  sv2v_dc_1430,sv2v_dc_1431,sv2v_dc_1432,sv2v_dc_1433,sv2v_dc_1434,sv2v_dc_1435,sv2v_dc_1436,
  sv2v_dc_1437,sv2v_dc_1438,sv2v_dc_1439,sv2v_dc_1440,sv2v_dc_1441,sv2v_dc_1442,
  sv2v_dc_1443,sv2v_dc_1444,sv2v_dc_1445,sv2v_dc_1446,sv2v_dc_1447,sv2v_dc_1448,
  sv2v_dc_1449,sv2v_dc_1450,sv2v_dc_1451,sv2v_dc_1452,sv2v_dc_1453,sv2v_dc_1454,
  sv2v_dc_1455,sv2v_dc_1456,sv2v_dc_1457,sv2v_dc_1458,sv2v_dc_1459,sv2v_dc_1460,
  sv2v_dc_1461,sv2v_dc_1462,sv2v_dc_1463,sv2v_dc_1464,sv2v_dc_1465,sv2v_dc_1466,
  sv2v_dc_1467,sv2v_dc_1468,sv2v_dc_1469,sv2v_dc_1470,sv2v_dc_1471,sv2v_dc_1472,sv2v_dc_1473,
  sv2v_dc_1474,sv2v_dc_1475,sv2v_dc_1476,sv2v_dc_1477,sv2v_dc_1478,sv2v_dc_1479,
  sv2v_dc_1480,sv2v_dc_1481,sv2v_dc_1482,sv2v_dc_1483,sv2v_dc_1484,sv2v_dc_1485,
  sv2v_dc_1486,sv2v_dc_1487,sv2v_dc_1488,sv2v_dc_1489,sv2v_dc_1490,sv2v_dc_1491,
  sv2v_dc_1492,sv2v_dc_1493,sv2v_dc_1494,sv2v_dc_1495,sv2v_dc_1496,sv2v_dc_1497,
  sv2v_dc_1498,sv2v_dc_1499,sv2v_dc_1500,sv2v_dc_1501,sv2v_dc_1502,sv2v_dc_1503,
  sv2v_dc_1504,sv2v_dc_1505,sv2v_dc_1506,sv2v_dc_1507,sv2v_dc_1508,sv2v_dc_1509,
  sv2v_dc_1510,sv2v_dc_1511,sv2v_dc_1512,sv2v_dc_1513,sv2v_dc_1514,sv2v_dc_1515,sv2v_dc_1516,
  sv2v_dc_1517,sv2v_dc_1518,sv2v_dc_1519,sv2v_dc_1520,sv2v_dc_1521,sv2v_dc_1522,
  sv2v_dc_1523,sv2v_dc_1524,sv2v_dc_1525,sv2v_dc_1526,sv2v_dc_1527,sv2v_dc_1528,
  sv2v_dc_1529,sv2v_dc_1530,sv2v_dc_1531,sv2v_dc_1532,sv2v_dc_1533,sv2v_dc_1534,
  sv2v_dc_1535,sv2v_dc_1536,sv2v_dc_1537,sv2v_dc_1538,sv2v_dc_1539,sv2v_dc_1540,
  sv2v_dc_1541,sv2v_dc_1542,sv2v_dc_1543,sv2v_dc_1544,sv2v_dc_1545,sv2v_dc_1546,
  sv2v_dc_1547,sv2v_dc_1548,sv2v_dc_1549,sv2v_dc_1550,sv2v_dc_1551,sv2v_dc_1552,sv2v_dc_1553,
  sv2v_dc_1554,sv2v_dc_1555,sv2v_dc_1556,sv2v_dc_1557,sv2v_dc_1558,sv2v_dc_1559,
  sv2v_dc_1560,sv2v_dc_1561,sv2v_dc_1562,sv2v_dc_1563,sv2v_dc_1564,sv2v_dc_1565,
  sv2v_dc_1566,sv2v_dc_1567,sv2v_dc_1568,sv2v_dc_1569,sv2v_dc_1570,sv2v_dc_1571,
  sv2v_dc_1572,sv2v_dc_1573,sv2v_dc_1574,sv2v_dc_1575,sv2v_dc_1576,sv2v_dc_1577,
  sv2v_dc_1578,sv2v_dc_1579,sv2v_dc_1580,sv2v_dc_1581,sv2v_dc_1582,sv2v_dc_1583,
  sv2v_dc_1584,sv2v_dc_1585,sv2v_dc_1586,sv2v_dc_1587,sv2v_dc_1588,sv2v_dc_1589,
  sv2v_dc_1590,sv2v_dc_1591,sv2v_dc_1592,sv2v_dc_1593,sv2v_dc_1594,sv2v_dc_1595,sv2v_dc_1596,
  sv2v_dc_1597,sv2v_dc_1598,sv2v_dc_1599,sv2v_dc_1600,sv2v_dc_1601,sv2v_dc_1602,
  sv2v_dc_1603,sv2v_dc_1604,sv2v_dc_1605,sv2v_dc_1606,sv2v_dc_1607,sv2v_dc_1608,
  sv2v_dc_1609,sv2v_dc_1610,sv2v_dc_1611,sv2v_dc_1612,sv2v_dc_1613,sv2v_dc_1614,
  sv2v_dc_1615,sv2v_dc_1616,sv2v_dc_1617,sv2v_dc_1618,sv2v_dc_1619,sv2v_dc_1620,
  sv2v_dc_1621,sv2v_dc_1622,sv2v_dc_1623,sv2v_dc_1624,sv2v_dc_1625,sv2v_dc_1626,
  sv2v_dc_1627,sv2v_dc_1628,sv2v_dc_1629,sv2v_dc_1630,sv2v_dc_1631,sv2v_dc_1632,sv2v_dc_1633,
  sv2v_dc_1634,sv2v_dc_1635,sv2v_dc_1636,sv2v_dc_1637,sv2v_dc_1638,sv2v_dc_1639,
  sv2v_dc_1640,sv2v_dc_1641,sv2v_dc_1642,sv2v_dc_1643,sv2v_dc_1644,sv2v_dc_1645,
  sv2v_dc_1646,sv2v_dc_1647,sv2v_dc_1648,sv2v_dc_1649,sv2v_dc_1650,sv2v_dc_1651,
  sv2v_dc_1652,sv2v_dc_1653,sv2v_dc_1654,sv2v_dc_1655,sv2v_dc_1656,sv2v_dc_1657,
  sv2v_dc_1658,sv2v_dc_1659,sv2v_dc_1660,sv2v_dc_1661,sv2v_dc_1662,sv2v_dc_1663,
  sv2v_dc_1664,sv2v_dc_1665,sv2v_dc_1666,sv2v_dc_1667,sv2v_dc_1668,sv2v_dc_1669,
  sv2v_dc_1670,sv2v_dc_1671,sv2v_dc_1672,sv2v_dc_1673,sv2v_dc_1674,sv2v_dc_1675,sv2v_dc_1676,
  sv2v_dc_1677,sv2v_dc_1678,sv2v_dc_1679,sv2v_dc_1680,sv2v_dc_1681,sv2v_dc_1682,
  sv2v_dc_1683,sv2v_dc_1684,sv2v_dc_1685,sv2v_dc_1686,sv2v_dc_1687,sv2v_dc_1688,
  sv2v_dc_1689,sv2v_dc_1690,sv2v_dc_1691,sv2v_dc_1692,sv2v_dc_1693,sv2v_dc_1694,
  sv2v_dc_1695,sv2v_dc_1696,sv2v_dc_1697,sv2v_dc_1698,sv2v_dc_1699,sv2v_dc_1700,
  sv2v_dc_1701,sv2v_dc_1702,sv2v_dc_1703,sv2v_dc_1704,sv2v_dc_1705,sv2v_dc_1706,
  sv2v_dc_1707,sv2v_dc_1708,sv2v_dc_1709,sv2v_dc_1710,sv2v_dc_1711,sv2v_dc_1712,sv2v_dc_1713,
  sv2v_dc_1714,sv2v_dc_1715,sv2v_dc_1716,sv2v_dc_1717,sv2v_dc_1718,sv2v_dc_1719,
  sv2v_dc_1720,sv2v_dc_1721,sv2v_dc_1722,sv2v_dc_1723,sv2v_dc_1724,sv2v_dc_1725,
  sv2v_dc_1726,sv2v_dc_1727,sv2v_dc_1728,sv2v_dc_1729,sv2v_dc_1730,sv2v_dc_1731,
  sv2v_dc_1732,sv2v_dc_1733,sv2v_dc_1734,sv2v_dc_1735,sv2v_dc_1736,sv2v_dc_1737,
  sv2v_dc_1738,sv2v_dc_1739,sv2v_dc_1740,sv2v_dc_1741,sv2v_dc_1742,sv2v_dc_1743,
  sv2v_dc_1744,sv2v_dc_1745,sv2v_dc_1746,sv2v_dc_1747,sv2v_dc_1748,sv2v_dc_1749,
  sv2v_dc_1750,sv2v_dc_1751,sv2v_dc_1752,sv2v_dc_1753,sv2v_dc_1754,sv2v_dc_1755,sv2v_dc_1756,
  sv2v_dc_1757,sv2v_dc_1758,sv2v_dc_1759,sv2v_dc_1760,sv2v_dc_1761,sv2v_dc_1762,
  sv2v_dc_1763,sv2v_dc_1764,sv2v_dc_1765,sv2v_dc_1766,sv2v_dc_1767,sv2v_dc_1768,
  sv2v_dc_1769,sv2v_dc_1770,sv2v_dc_1771,sv2v_dc_1772,sv2v_dc_1773,sv2v_dc_1774,
  sv2v_dc_1775,sv2v_dc_1776,sv2v_dc_1777,sv2v_dc_1778,sv2v_dc_1779,sv2v_dc_1780,
  sv2v_dc_1781,sv2v_dc_1782,sv2v_dc_1783,sv2v_dc_1784,sv2v_dc_1785,sv2v_dc_1786,
  sv2v_dc_1787,sv2v_dc_1788,sv2v_dc_1789,sv2v_dc_1790,sv2v_dc_1791,sv2v_dc_1792,sv2v_dc_1793,
  sv2v_dc_1794,sv2v_dc_1795,sv2v_dc_1796,sv2v_dc_1797,sv2v_dc_1798,sv2v_dc_1799,
  sv2v_dc_1800,sv2v_dc_1801,sv2v_dc_1802,sv2v_dc_1803,sv2v_dc_1804,sv2v_dc_1805,
  sv2v_dc_1806,sv2v_dc_1807,sv2v_dc_1808,sv2v_dc_1809,sv2v_dc_1810,sv2v_dc_1811,
  sv2v_dc_1812,sv2v_dc_1813,sv2v_dc_1814,sv2v_dc_1815,sv2v_dc_1816,sv2v_dc_1817,
  sv2v_dc_1818,sv2v_dc_1819,sv2v_dc_1820,sv2v_dc_1821,sv2v_dc_1822,sv2v_dc_1823,
  sv2v_dc_1824,sv2v_dc_1825,sv2v_dc_1826,sv2v_dc_1827,sv2v_dc_1828,sv2v_dc_1829,
  sv2v_dc_1830,sv2v_dc_1831,sv2v_dc_1832,sv2v_dc_1833,sv2v_dc_1834,sv2v_dc_1835,sv2v_dc_1836,
  sv2v_dc_1837,sv2v_dc_1838,sv2v_dc_1839,sv2v_dc_1840,sv2v_dc_1841,sv2v_dc_1842,
  sv2v_dc_1843,sv2v_dc_1844,sv2v_dc_1845,sv2v_dc_1846,sv2v_dc_1847,sv2v_dc_1848,
  sv2v_dc_1849,sv2v_dc_1850,sv2v_dc_1851,sv2v_dc_1852,sv2v_dc_1853,sv2v_dc_1854,
  sv2v_dc_1855,sv2v_dc_1856,sv2v_dc_1857,sv2v_dc_1858,sv2v_dc_1859,sv2v_dc_1860,
  sv2v_dc_1861,sv2v_dc_1862,sv2v_dc_1863,sv2v_dc_1864,sv2v_dc_1865,sv2v_dc_1866,
  sv2v_dc_1867,sv2v_dc_1868,sv2v_dc_1869,sv2v_dc_1870,sv2v_dc_1871,sv2v_dc_1872,sv2v_dc_1873,
  sv2v_dc_1874,sv2v_dc_1875,sv2v_dc_1876,sv2v_dc_1877,sv2v_dc_1878,sv2v_dc_1879,
  sv2v_dc_1880,sv2v_dc_1881,sv2v_dc_1882,sv2v_dc_1883,sv2v_dc_1884,sv2v_dc_1885,
  sv2v_dc_1886,sv2v_dc_1887,sv2v_dc_1888,sv2v_dc_1889,sv2v_dc_1890,sv2v_dc_1891,
  sv2v_dc_1892,sv2v_dc_1893,sv2v_dc_1894,sv2v_dc_1895,sv2v_dc_1896,sv2v_dc_1897,
  sv2v_dc_1898,sv2v_dc_1899,sv2v_dc_1900,sv2v_dc_1901,sv2v_dc_1902,sv2v_dc_1903,
  sv2v_dc_1904,sv2v_dc_1905,sv2v_dc_1906,sv2v_dc_1907,sv2v_dc_1908,sv2v_dc_1909,
  sv2v_dc_1910,sv2v_dc_1911,sv2v_dc_1912,sv2v_dc_1913,sv2v_dc_1914,sv2v_dc_1915,sv2v_dc_1916,
  sv2v_dc_1917,sv2v_dc_1918,sv2v_dc_1919,sv2v_dc_1920,sv2v_dc_1921,sv2v_dc_1922,
  sv2v_dc_1923,sv2v_dc_1924,sv2v_dc_1925,sv2v_dc_1926,sv2v_dc_1927,sv2v_dc_1928,
  sv2v_dc_1929,sv2v_dc_1930,sv2v_dc_1931,sv2v_dc_1932,sv2v_dc_1933,sv2v_dc_1934,
  sv2v_dc_1935,sv2v_dc_1936,sv2v_dc_1937,sv2v_dc_1938,sv2v_dc_1939,sv2v_dc_1940,
  sv2v_dc_1941,sv2v_dc_1942,sv2v_dc_1943,sv2v_dc_1944,sv2v_dc_1945,sv2v_dc_1946,
  sv2v_dc_1947,sv2v_dc_1948,sv2v_dc_1949,sv2v_dc_1950,sv2v_dc_1951,sv2v_dc_1952,sv2v_dc_1953,
  sv2v_dc_1954,sv2v_dc_1955,sv2v_dc_1956,sv2v_dc_1957,sv2v_dc_1958,sv2v_dc_1959,
  sv2v_dc_1960,sv2v_dc_1961,sv2v_dc_1962,sv2v_dc_1963,sv2v_dc_1964,sv2v_dc_1965,
  sv2v_dc_1966,sv2v_dc_1967,sv2v_dc_1968,sv2v_dc_1969,sv2v_dc_1970,sv2v_dc_1971,
  sv2v_dc_1972,sv2v_dc_1973,sv2v_dc_1974,sv2v_dc_1975,sv2v_dc_1976,sv2v_dc_1977,
  sv2v_dc_1978,sv2v_dc_1979,sv2v_dc_1980,sv2v_dc_1981,sv2v_dc_1982,sv2v_dc_1983,
  sv2v_dc_1984,sv2v_dc_1985,sv2v_dc_1986,sv2v_dc_1987,sv2v_dc_1988,sv2v_dc_1989,
  sv2v_dc_1990,sv2v_dc_1991,sv2v_dc_1992,sv2v_dc_1993,sv2v_dc_1994,sv2v_dc_1995,sv2v_dc_1996,
  sv2v_dc_1997,sv2v_dc_1998,sv2v_dc_1999,sv2v_dc_2000,sv2v_dc_2001,sv2v_dc_2002,
  sv2v_dc_2003,sv2v_dc_2004,sv2v_dc_2005,sv2v_dc_2006,sv2v_dc_2007,sv2v_dc_2008,
  sv2v_dc_2009,sv2v_dc_2010,sv2v_dc_2011,sv2v_dc_2012,sv2v_dc_2013,sv2v_dc_2014,
  sv2v_dc_2015,sv2v_dc_2016,sv2v_dc_2017,sv2v_dc_2018,sv2v_dc_2019,sv2v_dc_2020,
  sv2v_dc_2021,sv2v_dc_2022,sv2v_dc_2023,sv2v_dc_2024,sv2v_dc_2025,sv2v_dc_2026,
  sv2v_dc_2027,sv2v_dc_2028,sv2v_dc_2029,sv2v_dc_2030,sv2v_dc_2031,sv2v_dc_2032,sv2v_dc_2033,
  sv2v_dc_2034,sv2v_dc_2035,sv2v_dc_2036,sv2v_dc_2037,sv2v_dc_2038,sv2v_dc_2039,
  sv2v_dc_2040,sv2v_dc_2041,sv2v_dc_2042,sv2v_dc_2043,sv2v_dc_2044,sv2v_dc_2045,
  sv2v_dc_2046,sv2v_dc_2047,sv2v_dc_2048,sv2v_dc_2049,sv2v_dc_2050,sv2v_dc_2051,
  sv2v_dc_2052,sv2v_dc_2053,sv2v_dc_2054,sv2v_dc_2055,sv2v_dc_2056,sv2v_dc_2057,
  sv2v_dc_2058,sv2v_dc_2059,sv2v_dc_2060,sv2v_dc_2061,sv2v_dc_2062,sv2v_dc_2063,
  sv2v_dc_2064,sv2v_dc_2065,sv2v_dc_2066,sv2v_dc_2067,sv2v_dc_2068,sv2v_dc_2069,
  sv2v_dc_2070,sv2v_dc_2071,sv2v_dc_2072,sv2v_dc_2073,sv2v_dc_2074,sv2v_dc_2075,sv2v_dc_2076,
  sv2v_dc_2077,sv2v_dc_2078,sv2v_dc_2079,sv2v_dc_2080,sv2v_dc_2081,sv2v_dc_2082,
  sv2v_dc_2083,sv2v_dc_2084,sv2v_dc_2085,sv2v_dc_2086,sv2v_dc_2087,sv2v_dc_2088,
  sv2v_dc_2089,sv2v_dc_2090,sv2v_dc_2091,sv2v_dc_2092,sv2v_dc_2093,sv2v_dc_2094,
  sv2v_dc_2095,sv2v_dc_2096,sv2v_dc_2097,sv2v_dc_2098,sv2v_dc_2099,sv2v_dc_2100,
  sv2v_dc_2101,sv2v_dc_2102,sv2v_dc_2103,sv2v_dc_2104,sv2v_dc_2105,sv2v_dc_2106,
  sv2v_dc_2107,sv2v_dc_2108,sv2v_dc_2109,sv2v_dc_2110,sv2v_dc_2111,sv2v_dc_2112,sv2v_dc_2113,
  sv2v_dc_2114,sv2v_dc_2115,sv2v_dc_2116,sv2v_dc_2117,sv2v_dc_2118,sv2v_dc_2119,
  sv2v_dc_2120,sv2v_dc_2121,sv2v_dc_2122,sv2v_dc_2123,sv2v_dc_2124,sv2v_dc_2125,
  sv2v_dc_2126,sv2v_dc_2127,sv2v_dc_2128,sv2v_dc_2129,sv2v_dc_2130,sv2v_dc_2131,
  sv2v_dc_2132,sv2v_dc_2133,sv2v_dc_2134,sv2v_dc_2135,sv2v_dc_2136,sv2v_dc_2137,
  sv2v_dc_2138,sv2v_dc_2139,sv2v_dc_2140,sv2v_dc_2141,sv2v_dc_2142,sv2v_dc_2143,
  sv2v_dc_2144,sv2v_dc_2145,sv2v_dc_2146,sv2v_dc_2147,sv2v_dc_2148,sv2v_dc_2149,
  sv2v_dc_2150,sv2v_dc_2151,sv2v_dc_2152,sv2v_dc_2153,sv2v_dc_2154,sv2v_dc_2155,sv2v_dc_2156,
  sv2v_dc_2157,sv2v_dc_2158,sv2v_dc_2159,sv2v_dc_2160,sv2v_dc_2161,sv2v_dc_2162,
  sv2v_dc_2163,sv2v_dc_2164,sv2v_dc_2165,sv2v_dc_2166,sv2v_dc_2167,sv2v_dc_2168,
  sv2v_dc_2169,sv2v_dc_2170,sv2v_dc_2171,sv2v_dc_2172,sv2v_dc_2173,sv2v_dc_2174,
  sv2v_dc_2175,sv2v_dc_2176,sv2v_dc_2177,sv2v_dc_2178,sv2v_dc_2179,sv2v_dc_2180,
  sv2v_dc_2181,sv2v_dc_2182,sv2v_dc_2183,sv2v_dc_2184,sv2v_dc_2185,sv2v_dc_2186,
  sv2v_dc_2187,sv2v_dc_2188,sv2v_dc_2189,sv2v_dc_2190,sv2v_dc_2191,sv2v_dc_2192,sv2v_dc_2193,
  sv2v_dc_2194,sv2v_dc_2195,sv2v_dc_2196,sv2v_dc_2197,sv2v_dc_2198,sv2v_dc_2199,
  sv2v_dc_2200,sv2v_dc_2201,sv2v_dc_2202,sv2v_dc_2203,sv2v_dc_2204,sv2v_dc_2205,
  sv2v_dc_2206,sv2v_dc_2207,sv2v_dc_2208,sv2v_dc_2209,sv2v_dc_2210,sv2v_dc_2211,
  sv2v_dc_2212,sv2v_dc_2213,sv2v_dc_2214,sv2v_dc_2215,sv2v_dc_2216,sv2v_dc_2217,
  sv2v_dc_2218,sv2v_dc_2219,sv2v_dc_2220,sv2v_dc_2221,sv2v_dc_2222,sv2v_dc_2223,
  sv2v_dc_2224,sv2v_dc_2225,sv2v_dc_2226,sv2v_dc_2227,sv2v_dc_2228,sv2v_dc_2229,
  sv2v_dc_2230,sv2v_dc_2231,sv2v_dc_2232,sv2v_dc_2233,sv2v_dc_2234,sv2v_dc_2235,sv2v_dc_2236,
  sv2v_dc_2237,sv2v_dc_2238,sv2v_dc_2239,sv2v_dc_2240,sv2v_dc_2241,sv2v_dc_2242,
  sv2v_dc_2243,sv2v_dc_2244,sv2v_dc_2245,sv2v_dc_2246,sv2v_dc_2247,sv2v_dc_2248,
  sv2v_dc_2249,sv2v_dc_2250,sv2v_dc_2251,sv2v_dc_2252,sv2v_dc_2253,sv2v_dc_2254,
  sv2v_dc_2255,sv2v_dc_2256,sv2v_dc_2257,sv2v_dc_2258,sv2v_dc_2259,sv2v_dc_2260,
  sv2v_dc_2261,sv2v_dc_2262,sv2v_dc_2263,sv2v_dc_2264,sv2v_dc_2265,sv2v_dc_2266,
  sv2v_dc_2267,sv2v_dc_2268,sv2v_dc_2269,sv2v_dc_2270,sv2v_dc_2271,sv2v_dc_2272,sv2v_dc_2273,
  sv2v_dc_2274,sv2v_dc_2275,sv2v_dc_2276,sv2v_dc_2277,sv2v_dc_2278,sv2v_dc_2279,
  sv2v_dc_2280,sv2v_dc_2281,sv2v_dc_2282,sv2v_dc_2283,sv2v_dc_2284,sv2v_dc_2285,
  sv2v_dc_2286,sv2v_dc_2287,sv2v_dc_2288,sv2v_dc_2289,sv2v_dc_2290,sv2v_dc_2291,
  sv2v_dc_2292,sv2v_dc_2293,sv2v_dc_2294,sv2v_dc_2295,sv2v_dc_2296,sv2v_dc_2297,
  sv2v_dc_2298,sv2v_dc_2299,sv2v_dc_2300,sv2v_dc_2301,sv2v_dc_2302,sv2v_dc_2303,
  sv2v_dc_2304,sv2v_dc_2305,sv2v_dc_2306,sv2v_dc_2307,sv2v_dc_2308,sv2v_dc_2309,
  sv2v_dc_2310,sv2v_dc_2311,sv2v_dc_2312,sv2v_dc_2313,sv2v_dc_2314,sv2v_dc_2315,sv2v_dc_2316,
  sv2v_dc_2317,sv2v_dc_2318,sv2v_dc_2319,sv2v_dc_2320,sv2v_dc_2321,sv2v_dc_2322,
  sv2v_dc_2323,sv2v_dc_2324,sv2v_dc_2325,sv2v_dc_2326,sv2v_dc_2327,sv2v_dc_2328,
  sv2v_dc_2329,sv2v_dc_2330,sv2v_dc_2331,sv2v_dc_2332,sv2v_dc_2333,sv2v_dc_2334,
  sv2v_dc_2335,sv2v_dc_2336,sv2v_dc_2337,sv2v_dc_2338,sv2v_dc_2339,sv2v_dc_2340,
  sv2v_dc_2341,sv2v_dc_2342,sv2v_dc_2343,sv2v_dc_2344,sv2v_dc_2345,sv2v_dc_2346,
  sv2v_dc_2347,sv2v_dc_2348,sv2v_dc_2349,sv2v_dc_2350,sv2v_dc_2351,sv2v_dc_2352,sv2v_dc_2353,
  sv2v_dc_2354,sv2v_dc_2355,sv2v_dc_2356,sv2v_dc_2357,sv2v_dc_2358,sv2v_dc_2359,
  sv2v_dc_2360,sv2v_dc_2361,sv2v_dc_2362,sv2v_dc_2363,sv2v_dc_2364,sv2v_dc_2365,
  sv2v_dc_2366,sv2v_dc_2367,sv2v_dc_2368,sv2v_dc_2369,sv2v_dc_2370,sv2v_dc_2371,
  sv2v_dc_2372,sv2v_dc_2373,sv2v_dc_2374,sv2v_dc_2375,sv2v_dc_2376,sv2v_dc_2377,
  sv2v_dc_2378,sv2v_dc_2379,sv2v_dc_2380,sv2v_dc_2381,sv2v_dc_2382,sv2v_dc_2383,
  sv2v_dc_2384,sv2v_dc_2385,sv2v_dc_2386,sv2v_dc_2387,sv2v_dc_2388,sv2v_dc_2389,
  sv2v_dc_2390,sv2v_dc_2391,sv2v_dc_2392,sv2v_dc_2393,sv2v_dc_2394,sv2v_dc_2395,sv2v_dc_2396,
  sv2v_dc_2397,sv2v_dc_2398,sv2v_dc_2399,sv2v_dc_2400,sv2v_dc_2401,sv2v_dc_2402,
  sv2v_dc_2403,sv2v_dc_2404,sv2v_dc_2405,sv2v_dc_2406,sv2v_dc_2407,sv2v_dc_2408,
  sv2v_dc_2409,sv2v_dc_2410,sv2v_dc_2411,sv2v_dc_2412,sv2v_dc_2413,sv2v_dc_2414,
  sv2v_dc_2415,sv2v_dc_2416,sv2v_dc_2417,sv2v_dc_2418,sv2v_dc_2419,sv2v_dc_2420,
  sv2v_dc_2421,sv2v_dc_2422,sv2v_dc_2423,sv2v_dc_2424,sv2v_dc_2425,sv2v_dc_2426,
  sv2v_dc_2427,sv2v_dc_2428,sv2v_dc_2429,sv2v_dc_2430,sv2v_dc_2431,sv2v_dc_2432,sv2v_dc_2433,
  sv2v_dc_2434,sv2v_dc_2435,sv2v_dc_2436,sv2v_dc_2437,sv2v_dc_2438,sv2v_dc_2439,
  sv2v_dc_2440,sv2v_dc_2441,sv2v_dc_2442,sv2v_dc_2443,sv2v_dc_2444,sv2v_dc_2445,
  sv2v_dc_2446,sv2v_dc_2447,sv2v_dc_2448,sv2v_dc_2449,sv2v_dc_2450,sv2v_dc_2451,
  sv2v_dc_2452,sv2v_dc_2453,sv2v_dc_2454,sv2v_dc_2455,sv2v_dc_2456,sv2v_dc_2457,
  sv2v_dc_2458,sv2v_dc_2459,sv2v_dc_2460,sv2v_dc_2461,sv2v_dc_2462,sv2v_dc_2463,
  sv2v_dc_2464,sv2v_dc_2465,sv2v_dc_2466,sv2v_dc_2467,sv2v_dc_2468,sv2v_dc_2469,
  sv2v_dc_2470,sv2v_dc_2471,sv2v_dc_2472,sv2v_dc_2473,sv2v_dc_2474,sv2v_dc_2475,sv2v_dc_2476,
  sv2v_dc_2477,sv2v_dc_2478,sv2v_dc_2479,sv2v_dc_2480,sv2v_dc_2481,sv2v_dc_2482,
  sv2v_dc_2483,sv2v_dc_2484,sv2v_dc_2485,sv2v_dc_2486,sv2v_dc_2487,sv2v_dc_2488,
  sv2v_dc_2489,sv2v_dc_2490,sv2v_dc_2491,sv2v_dc_2492,sv2v_dc_2493,sv2v_dc_2494,
  sv2v_dc_2495,sv2v_dc_2496,sv2v_dc_2497,sv2v_dc_2498,sv2v_dc_2499,sv2v_dc_2500,
  sv2v_dc_2501,sv2v_dc_2502,sv2v_dc_2503,sv2v_dc_2504,sv2v_dc_2505,sv2v_dc_2506,
  sv2v_dc_2507,sv2v_dc_2508,sv2v_dc_2509,sv2v_dc_2510,sv2v_dc_2511,sv2v_dc_2512,sv2v_dc_2513,
  sv2v_dc_2514,sv2v_dc_2515,sv2v_dc_2516,sv2v_dc_2517,sv2v_dc_2518,sv2v_dc_2519,
  sv2v_dc_2520,sv2v_dc_2521,sv2v_dc_2522,sv2v_dc_2523,sv2v_dc_2524,sv2v_dc_2525,
  sv2v_dc_2526,sv2v_dc_2527,sv2v_dc_2528,sv2v_dc_2529,sv2v_dc_2530,sv2v_dc_2531,
  sv2v_dc_2532,sv2v_dc_2533,sv2v_dc_2534,sv2v_dc_2535,sv2v_dc_2536,sv2v_dc_2537,
  sv2v_dc_2538,sv2v_dc_2539,sv2v_dc_2540,sv2v_dc_2541,sv2v_dc_2542,sv2v_dc_2543,
  sv2v_dc_2544,sv2v_dc_2545,sv2v_dc_2546,sv2v_dc_2547,sv2v_dc_2548,sv2v_dc_2549,
  sv2v_dc_2550,sv2v_dc_2551,sv2v_dc_2552,sv2v_dc_2553,sv2v_dc_2554,sv2v_dc_2555,sv2v_dc_2556,
  sv2v_dc_2557,sv2v_dc_2558,sv2v_dc_2559,sv2v_dc_2560,sv2v_dc_2561,sv2v_dc_2562,
  sv2v_dc_2563,sv2v_dc_2564,sv2v_dc_2565,sv2v_dc_2566,sv2v_dc_2567,sv2v_dc_2568,
  sv2v_dc_2569,sv2v_dc_2570,sv2v_dc_2571,sv2v_dc_2572,sv2v_dc_2573,sv2v_dc_2574,
  sv2v_dc_2575,sv2v_dc_2576,sv2v_dc_2577,sv2v_dc_2578,sv2v_dc_2579,sv2v_dc_2580,
  sv2v_dc_2581,sv2v_dc_2582,sv2v_dc_2583,sv2v_dc_2584,sv2v_dc_2585,sv2v_dc_2586,
  sv2v_dc_2587,sv2v_dc_2588,sv2v_dc_2589,sv2v_dc_2590,sv2v_dc_2591,sv2v_dc_2592,sv2v_dc_2593,
  sv2v_dc_2594,sv2v_dc_2595,sv2v_dc_2596,sv2v_dc_2597,sv2v_dc_2598,sv2v_dc_2599,
  sv2v_dc_2600,sv2v_dc_2601,sv2v_dc_2602,sv2v_dc_2603,sv2v_dc_2604,sv2v_dc_2605,
  sv2v_dc_2606,sv2v_dc_2607,sv2v_dc_2608,sv2v_dc_2609,sv2v_dc_2610,sv2v_dc_2611,
  sv2v_dc_2612,sv2v_dc_2613,sv2v_dc_2614,sv2v_dc_2615,sv2v_dc_2616,sv2v_dc_2617,
  sv2v_dc_2618,sv2v_dc_2619,sv2v_dc_2620,sv2v_dc_2621,sv2v_dc_2622,sv2v_dc_2623,
  sv2v_dc_2624,sv2v_dc_2625,sv2v_dc_2626,sv2v_dc_2627,sv2v_dc_2628,sv2v_dc_2629,
  sv2v_dc_2630,sv2v_dc_2631,sv2v_dc_2632,sv2v_dc_2633,sv2v_dc_2634,sv2v_dc_2635,sv2v_dc_2636,
  sv2v_dc_2637,sv2v_dc_2638,sv2v_dc_2639,sv2v_dc_2640,sv2v_dc_2641,sv2v_dc_2642,
  sv2v_dc_2643,sv2v_dc_2644,sv2v_dc_2645,sv2v_dc_2646,sv2v_dc_2647,sv2v_dc_2648,
  sv2v_dc_2649,sv2v_dc_2650,sv2v_dc_2651,sv2v_dc_2652,sv2v_dc_2653,sv2v_dc_2654,
  sv2v_dc_2655,sv2v_dc_2656,sv2v_dc_2657,sv2v_dc_2658,sv2v_dc_2659,sv2v_dc_2660,
  sv2v_dc_2661,sv2v_dc_2662,sv2v_dc_2663,sv2v_dc_2664,sv2v_dc_2665,sv2v_dc_2666,
  sv2v_dc_2667,sv2v_dc_2668,sv2v_dc_2669,sv2v_dc_2670,sv2v_dc_2671,sv2v_dc_2672,sv2v_dc_2673,
  sv2v_dc_2674,sv2v_dc_2675,sv2v_dc_2676,sv2v_dc_2677,sv2v_dc_2678,sv2v_dc_2679,
  sv2v_dc_2680,sv2v_dc_2681,sv2v_dc_2682,sv2v_dc_2683,sv2v_dc_2684,sv2v_dc_2685,
  sv2v_dc_2686,sv2v_dc_2687,sv2v_dc_2688,sv2v_dc_2689,sv2v_dc_2690,sv2v_dc_2691,
  sv2v_dc_2692,sv2v_dc_2693,sv2v_dc_2694,sv2v_dc_2695,sv2v_dc_2696,sv2v_dc_2697,
  sv2v_dc_2698,sv2v_dc_2699,sv2v_dc_2700,sv2v_dc_2701,sv2v_dc_2702,sv2v_dc_2703,
  sv2v_dc_2704,sv2v_dc_2705,sv2v_dc_2706,sv2v_dc_2707,sv2v_dc_2708,sv2v_dc_2709,
  sv2v_dc_2710,sv2v_dc_2711,sv2v_dc_2712,sv2v_dc_2713,sv2v_dc_2714,sv2v_dc_2715,sv2v_dc_2716,
  sv2v_dc_2717,sv2v_dc_2718,sv2v_dc_2719,sv2v_dc_2720,sv2v_dc_2721,sv2v_dc_2722,
  sv2v_dc_2723,sv2v_dc_2724,sv2v_dc_2725,sv2v_dc_2726,sv2v_dc_2727,sv2v_dc_2728,
  sv2v_dc_2729,sv2v_dc_2730,sv2v_dc_2731,sv2v_dc_2732,sv2v_dc_2733,sv2v_dc_2734,
  sv2v_dc_2735,sv2v_dc_2736,sv2v_dc_2737,sv2v_dc_2738,sv2v_dc_2739,sv2v_dc_2740,
  sv2v_dc_2741,sv2v_dc_2742,sv2v_dc_2743,sv2v_dc_2744,sv2v_dc_2745,sv2v_dc_2746,
  sv2v_dc_2747,sv2v_dc_2748,sv2v_dc_2749,sv2v_dc_2750,sv2v_dc_2751,sv2v_dc_2752,sv2v_dc_2753,
  sv2v_dc_2754,sv2v_dc_2755,sv2v_dc_2756,sv2v_dc_2757,sv2v_dc_2758,sv2v_dc_2759,
  sv2v_dc_2760,sv2v_dc_2761,sv2v_dc_2762,sv2v_dc_2763,sv2v_dc_2764,sv2v_dc_2765,
  sv2v_dc_2766,sv2v_dc_2767,sv2v_dc_2768,sv2v_dc_2769,sv2v_dc_2770,sv2v_dc_2771,
  sv2v_dc_2772,sv2v_dc_2773,sv2v_dc_2774,sv2v_dc_2775,sv2v_dc_2776,sv2v_dc_2777,
  sv2v_dc_2778,sv2v_dc_2779,sv2v_dc_2780,sv2v_dc_2781,sv2v_dc_2782,sv2v_dc_2783,
  sv2v_dc_2784,sv2v_dc_2785,sv2v_dc_2786,sv2v_dc_2787,sv2v_dc_2788,sv2v_dc_2789,
  sv2v_dc_2790,sv2v_dc_2791,sv2v_dc_2792,sv2v_dc_2793,sv2v_dc_2794,sv2v_dc_2795,sv2v_dc_2796,
  sv2v_dc_2797,sv2v_dc_2798,sv2v_dc_2799,sv2v_dc_2800,sv2v_dc_2801,sv2v_dc_2802,
  sv2v_dc_2803,sv2v_dc_2804,sv2v_dc_2805,sv2v_dc_2806,sv2v_dc_2807,sv2v_dc_2808,
  sv2v_dc_2809,sv2v_dc_2810,sv2v_dc_2811,sv2v_dc_2812,sv2v_dc_2813,sv2v_dc_2814,
  sv2v_dc_2815,sv2v_dc_2816,sv2v_dc_2817,sv2v_dc_2818,sv2v_dc_2819,sv2v_dc_2820,
  sv2v_dc_2821,sv2v_dc_2822,sv2v_dc_2823,sv2v_dc_2824,sv2v_dc_2825,sv2v_dc_2826,
  sv2v_dc_2827,sv2v_dc_2828,sv2v_dc_2829,sv2v_dc_2830,sv2v_dc_2831,sv2v_dc_2832,sv2v_dc_2833,
  sv2v_dc_2834,sv2v_dc_2835,sv2v_dc_2836,sv2v_dc_2837,sv2v_dc_2838,sv2v_dc_2839,
  sv2v_dc_2840,sv2v_dc_2841,sv2v_dc_2842,sv2v_dc_2843,sv2v_dc_2844,sv2v_dc_2845,
  sv2v_dc_2846,sv2v_dc_2847,sv2v_dc_2848,sv2v_dc_2849,sv2v_dc_2850,sv2v_dc_2851,
  sv2v_dc_2852,sv2v_dc_2853,sv2v_dc_2854,sv2v_dc_2855,sv2v_dc_2856,sv2v_dc_2857,
  sv2v_dc_2858,sv2v_dc_2859,sv2v_dc_2860,sv2v_dc_2861,sv2v_dc_2862,sv2v_dc_2863,
  sv2v_dc_2864,sv2v_dc_2865,sv2v_dc_2866,sv2v_dc_2867,sv2v_dc_2868,sv2v_dc_2869,
  sv2v_dc_2870,sv2v_dc_2871,sv2v_dc_2872,sv2v_dc_2873,sv2v_dc_2874,sv2v_dc_2875,sv2v_dc_2876,
  sv2v_dc_2877,sv2v_dc_2878,sv2v_dc_2879,sv2v_dc_2880,sv2v_dc_2881,sv2v_dc_2882,
  sv2v_dc_2883,sv2v_dc_2884,sv2v_dc_2885,sv2v_dc_2886,sv2v_dc_2887,sv2v_dc_2888,
  sv2v_dc_2889,sv2v_dc_2890,sv2v_dc_2891,sv2v_dc_2892,sv2v_dc_2893,sv2v_dc_2894,
  sv2v_dc_2895,sv2v_dc_2896,sv2v_dc_2897,sv2v_dc_2898,sv2v_dc_2899,sv2v_dc_2900,
  sv2v_dc_2901,sv2v_dc_2902,sv2v_dc_2903,sv2v_dc_2904,sv2v_dc_2905,sv2v_dc_2906,
  sv2v_dc_2907,sv2v_dc_2908,sv2v_dc_2909,sv2v_dc_2910,sv2v_dc_2911,sv2v_dc_2912,sv2v_dc_2913,
  sv2v_dc_2914,sv2v_dc_2915,sv2v_dc_2916,sv2v_dc_2917,sv2v_dc_2918,sv2v_dc_2919,
  sv2v_dc_2920,sv2v_dc_2921,sv2v_dc_2922,sv2v_dc_2923,sv2v_dc_2924,sv2v_dc_2925,
  sv2v_dc_2926,sv2v_dc_2927,sv2v_dc_2928,sv2v_dc_2929,sv2v_dc_2930,sv2v_dc_2931,
  sv2v_dc_2932,sv2v_dc_2933,sv2v_dc_2934,sv2v_dc_2935,sv2v_dc_2936,sv2v_dc_2937,
  sv2v_dc_2938,sv2v_dc_2939,sv2v_dc_2940,sv2v_dc_2941,sv2v_dc_2942,sv2v_dc_2943,
  sv2v_dc_2944,sv2v_dc_2945,sv2v_dc_2946,sv2v_dc_2947,sv2v_dc_2948,sv2v_dc_2949,
  sv2v_dc_2950,sv2v_dc_2951,sv2v_dc_2952,sv2v_dc_2953,sv2v_dc_2954,sv2v_dc_2955,sv2v_dc_2956,
  sv2v_dc_2957,sv2v_dc_2958,sv2v_dc_2959,sv2v_dc_2960,sv2v_dc_2961,sv2v_dc_2962,
  sv2v_dc_2963,sv2v_dc_2964,sv2v_dc_2965,sv2v_dc_2966,sv2v_dc_2967,sv2v_dc_2968,
  sv2v_dc_2969,sv2v_dc_2970,sv2v_dc_2971,sv2v_dc_2972,sv2v_dc_2973,sv2v_dc_2974,
  sv2v_dc_2975,sv2v_dc_2976,sv2v_dc_2977,sv2v_dc_2978,sv2v_dc_2979,sv2v_dc_2980,
  sv2v_dc_2981,sv2v_dc_2982,sv2v_dc_2983,sv2v_dc_2984,sv2v_dc_2985,sv2v_dc_2986,
  sv2v_dc_2987,sv2v_dc_2988,sv2v_dc_2989,sv2v_dc_2990,sv2v_dc_2991,sv2v_dc_2992,sv2v_dc_2993,
  sv2v_dc_2994,sv2v_dc_2995,sv2v_dc_2996,sv2v_dc_2997,sv2v_dc_2998,sv2v_dc_2999,
  sv2v_dc_3000,sv2v_dc_3001,sv2v_dc_3002,sv2v_dc_3003,sv2v_dc_3004,sv2v_dc_3005,
  sv2v_dc_3006,sv2v_dc_3007,sv2v_dc_3008,sv2v_dc_3009,sv2v_dc_3010,sv2v_dc_3011,
  sv2v_dc_3012,sv2v_dc_3013,sv2v_dc_3014,sv2v_dc_3015,sv2v_dc_3016,sv2v_dc_3017,
  sv2v_dc_3018,sv2v_dc_3019,sv2v_dc_3020,sv2v_dc_3021,sv2v_dc_3022,sv2v_dc_3023,
  sv2v_dc_3024,sv2v_dc_3025,sv2v_dc_3026,sv2v_dc_3027,sv2v_dc_3028,sv2v_dc_3029,
  sv2v_dc_3030,sv2v_dc_3031,sv2v_dc_3032,sv2v_dc_3033,sv2v_dc_3034,sv2v_dc_3035,sv2v_dc_3036,
  sv2v_dc_3037,sv2v_dc_3038,sv2v_dc_3039,sv2v_dc_3040,sv2v_dc_3041,sv2v_dc_3042,
  sv2v_dc_3043,sv2v_dc_3044,sv2v_dc_3045,sv2v_dc_3046,sv2v_dc_3047,sv2v_dc_3048,
  sv2v_dc_3049,sv2v_dc_3050,sv2v_dc_3051,sv2v_dc_3052,sv2v_dc_3053,sv2v_dc_3054,
  sv2v_dc_3055,sv2v_dc_3056,sv2v_dc_3057,sv2v_dc_3058,sv2v_dc_3059,sv2v_dc_3060,
  sv2v_dc_3061,sv2v_dc_3062,sv2v_dc_3063,sv2v_dc_3064,sv2v_dc_3065,sv2v_dc_3066,
  sv2v_dc_3067,sv2v_dc_3068,sv2v_dc_3069,sv2v_dc_3070;

  reverse_width54
  reverse
  (
    .in(reverseOut),
    .out(out)
  );

  assign { sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36, sv2v_dc_37, sv2v_dc_38, sv2v_dc_39, sv2v_dc_40, sv2v_dc_41, sv2v_dc_42, sv2v_dc_43, sv2v_dc_44, sv2v_dc_45, sv2v_dc_46, sv2v_dc_47, sv2v_dc_48, sv2v_dc_49, sv2v_dc_50, sv2v_dc_51, sv2v_dc_52, sv2v_dc_53, sv2v_dc_54, sv2v_dc_55, sv2v_dc_56, sv2v_dc_57, sv2v_dc_58, sv2v_dc_59, sv2v_dc_60, sv2v_dc_61, sv2v_dc_62, sv2v_dc_63, sv2v_dc_64, sv2v_dc_65, sv2v_dc_66, sv2v_dc_67, sv2v_dc_68, sv2v_dc_69, sv2v_dc_70, sv2v_dc_71, sv2v_dc_72, sv2v_dc_73, sv2v_dc_74, sv2v_dc_75, sv2v_dc_76, sv2v_dc_77, sv2v_dc_78, sv2v_dc_79, sv2v_dc_80, sv2v_dc_81, sv2v_dc_82, sv2v_dc_83, sv2v_dc_84, sv2v_dc_85, sv2v_dc_86, sv2v_dc_87, sv2v_dc_88, sv2v_dc_89, sv2v_dc_90, sv2v_dc_91, sv2v_dc_92, sv2v_dc_93, sv2v_dc_94, sv2v_dc_95, sv2v_dc_96, sv2v_dc_97, sv2v_dc_98, sv2v_dc_99, sv2v_dc_100, sv2v_dc_101, sv2v_dc_102, sv2v_dc_103, sv2v_dc_104, sv2v_dc_105, sv2v_dc_106, sv2v_dc_107, sv2v_dc_108, sv2v_dc_109, sv2v_dc_110, sv2v_dc_111, sv2v_dc_112, sv2v_dc_113, sv2v_dc_114, sv2v_dc_115, sv2v_dc_116, sv2v_dc_117, sv2v_dc_118, sv2v_dc_119, sv2v_dc_120, sv2v_dc_121, sv2v_dc_122, sv2v_dc_123, sv2v_dc_124, sv2v_dc_125, sv2v_dc_126, sv2v_dc_127, sv2v_dc_128, sv2v_dc_129, sv2v_dc_130, sv2v_dc_131, sv2v_dc_132, sv2v_dc_133, sv2v_dc_134, sv2v_dc_135, sv2v_dc_136, sv2v_dc_137, sv2v_dc_138, sv2v_dc_139, sv2v_dc_140, sv2v_dc_141, sv2v_dc_142, sv2v_dc_143, sv2v_dc_144, sv2v_dc_145, sv2v_dc_146, sv2v_dc_147, sv2v_dc_148, sv2v_dc_149, sv2v_dc_150, sv2v_dc_151, sv2v_dc_152, sv2v_dc_153, sv2v_dc_154, sv2v_dc_155, sv2v_dc_156, sv2v_dc_157, sv2v_dc_158, sv2v_dc_159, sv2v_dc_160, sv2v_dc_161, sv2v_dc_162, sv2v_dc_163, sv2v_dc_164, sv2v_dc_165, sv2v_dc_166, sv2v_dc_167, sv2v_dc_168, sv2v_dc_169, sv2v_dc_170, sv2v_dc_171, sv2v_dc_172, sv2v_dc_173, sv2v_dc_174, sv2v_dc_175, sv2v_dc_176, sv2v_dc_177, sv2v_dc_178, sv2v_dc_179, sv2v_dc_180, sv2v_dc_181, sv2v_dc_182, sv2v_dc_183, sv2v_dc_184, sv2v_dc_185, sv2v_dc_186, sv2v_dc_187, sv2v_dc_188, sv2v_dc_189, sv2v_dc_190, sv2v_dc_191, sv2v_dc_192, sv2v_dc_193, sv2v_dc_194, sv2v_dc_195, sv2v_dc_196, sv2v_dc_197, sv2v_dc_198, sv2v_dc_199, sv2v_dc_200, sv2v_dc_201, sv2v_dc_202, sv2v_dc_203, sv2v_dc_204, sv2v_dc_205, sv2v_dc_206, sv2v_dc_207, sv2v_dc_208, sv2v_dc_209, sv2v_dc_210, sv2v_dc_211, sv2v_dc_212, sv2v_dc_213, sv2v_dc_214, sv2v_dc_215, sv2v_dc_216, sv2v_dc_217, sv2v_dc_218, sv2v_dc_219, sv2v_dc_220, sv2v_dc_221, sv2v_dc_222, sv2v_dc_223, sv2v_dc_224, sv2v_dc_225, sv2v_dc_226, sv2v_dc_227, sv2v_dc_228, sv2v_dc_229, sv2v_dc_230, sv2v_dc_231, sv2v_dc_232, sv2v_dc_233, sv2v_dc_234, sv2v_dc_235, sv2v_dc_236, sv2v_dc_237, sv2v_dc_238, sv2v_dc_239, sv2v_dc_240, sv2v_dc_241, sv2v_dc_242, sv2v_dc_243, sv2v_dc_244, sv2v_dc_245, sv2v_dc_246, sv2v_dc_247, sv2v_dc_248, sv2v_dc_249, sv2v_dc_250, sv2v_dc_251, sv2v_dc_252, sv2v_dc_253, sv2v_dc_254, sv2v_dc_255, sv2v_dc_256, sv2v_dc_257, sv2v_dc_258, sv2v_dc_259, sv2v_dc_260, sv2v_dc_261, sv2v_dc_262, sv2v_dc_263, sv2v_dc_264, sv2v_dc_265, sv2v_dc_266, sv2v_dc_267, sv2v_dc_268, sv2v_dc_269, sv2v_dc_270, sv2v_dc_271, sv2v_dc_272, sv2v_dc_273, sv2v_dc_274, sv2v_dc_275, sv2v_dc_276, sv2v_dc_277, sv2v_dc_278, sv2v_dc_279, sv2v_dc_280, sv2v_dc_281, sv2v_dc_282, sv2v_dc_283, sv2v_dc_284, sv2v_dc_285, sv2v_dc_286, sv2v_dc_287, sv2v_dc_288, sv2v_dc_289, sv2v_dc_290, sv2v_dc_291, sv2v_dc_292, sv2v_dc_293, sv2v_dc_294, sv2v_dc_295, sv2v_dc_296, sv2v_dc_297, sv2v_dc_298, sv2v_dc_299, sv2v_dc_300, sv2v_dc_301, sv2v_dc_302, sv2v_dc_303, sv2v_dc_304, sv2v_dc_305, sv2v_dc_306, sv2v_dc_307, sv2v_dc_308, sv2v_dc_309, sv2v_dc_310, sv2v_dc_311, sv2v_dc_312, sv2v_dc_313, sv2v_dc_314, sv2v_dc_315, sv2v_dc_316, sv2v_dc_317, sv2v_dc_318, sv2v_dc_319, sv2v_dc_320, sv2v_dc_321, sv2v_dc_322, sv2v_dc_323, sv2v_dc_324, sv2v_dc_325, sv2v_dc_326, sv2v_dc_327, sv2v_dc_328, sv2v_dc_329, sv2v_dc_330, sv2v_dc_331, sv2v_dc_332, sv2v_dc_333, sv2v_dc_334, sv2v_dc_335, sv2v_dc_336, sv2v_dc_337, sv2v_dc_338, sv2v_dc_339, sv2v_dc_340, sv2v_dc_341, sv2v_dc_342, sv2v_dc_343, sv2v_dc_344, sv2v_dc_345, sv2v_dc_346, sv2v_dc_347, sv2v_dc_348, sv2v_dc_349, sv2v_dc_350, sv2v_dc_351, sv2v_dc_352, sv2v_dc_353, sv2v_dc_354, sv2v_dc_355, sv2v_dc_356, sv2v_dc_357, sv2v_dc_358, sv2v_dc_359, sv2v_dc_360, sv2v_dc_361, sv2v_dc_362, sv2v_dc_363, sv2v_dc_364, sv2v_dc_365, sv2v_dc_366, sv2v_dc_367, sv2v_dc_368, sv2v_dc_369, sv2v_dc_370, sv2v_dc_371, sv2v_dc_372, sv2v_dc_373, sv2v_dc_374, sv2v_dc_375, sv2v_dc_376, sv2v_dc_377, sv2v_dc_378, sv2v_dc_379, sv2v_dc_380, sv2v_dc_381, sv2v_dc_382, sv2v_dc_383, sv2v_dc_384, sv2v_dc_385, sv2v_dc_386, sv2v_dc_387, sv2v_dc_388, sv2v_dc_389, sv2v_dc_390, sv2v_dc_391, sv2v_dc_392, sv2v_dc_393, sv2v_dc_394, sv2v_dc_395, sv2v_dc_396, sv2v_dc_397, sv2v_dc_398, sv2v_dc_399, sv2v_dc_400, sv2v_dc_401, sv2v_dc_402, sv2v_dc_403, sv2v_dc_404, sv2v_dc_405, sv2v_dc_406, sv2v_dc_407, sv2v_dc_408, sv2v_dc_409, sv2v_dc_410, sv2v_dc_411, sv2v_dc_412, sv2v_dc_413, sv2v_dc_414, sv2v_dc_415, sv2v_dc_416, sv2v_dc_417, sv2v_dc_418, sv2v_dc_419, sv2v_dc_420, sv2v_dc_421, sv2v_dc_422, sv2v_dc_423, sv2v_dc_424, sv2v_dc_425, sv2v_dc_426, sv2v_dc_427, sv2v_dc_428, sv2v_dc_429, sv2v_dc_430, sv2v_dc_431, sv2v_dc_432, sv2v_dc_433, sv2v_dc_434, sv2v_dc_435, sv2v_dc_436, sv2v_dc_437, sv2v_dc_438, sv2v_dc_439, sv2v_dc_440, sv2v_dc_441, sv2v_dc_442, sv2v_dc_443, sv2v_dc_444, sv2v_dc_445, sv2v_dc_446, sv2v_dc_447, sv2v_dc_448, sv2v_dc_449, sv2v_dc_450, sv2v_dc_451, sv2v_dc_452, sv2v_dc_453, sv2v_dc_454, sv2v_dc_455, sv2v_dc_456, sv2v_dc_457, sv2v_dc_458, sv2v_dc_459, sv2v_dc_460, sv2v_dc_461, sv2v_dc_462, sv2v_dc_463, sv2v_dc_464, sv2v_dc_465, sv2v_dc_466, sv2v_dc_467, sv2v_dc_468, sv2v_dc_469, sv2v_dc_470, sv2v_dc_471, sv2v_dc_472, sv2v_dc_473, sv2v_dc_474, sv2v_dc_475, sv2v_dc_476, sv2v_dc_477, sv2v_dc_478, sv2v_dc_479, sv2v_dc_480, sv2v_dc_481, sv2v_dc_482, sv2v_dc_483, sv2v_dc_484, sv2v_dc_485, sv2v_dc_486, sv2v_dc_487, sv2v_dc_488, sv2v_dc_489, sv2v_dc_490, sv2v_dc_491, sv2v_dc_492, sv2v_dc_493, sv2v_dc_494, sv2v_dc_495, sv2v_dc_496, sv2v_dc_497, sv2v_dc_498, sv2v_dc_499, sv2v_dc_500, sv2v_dc_501, sv2v_dc_502, sv2v_dc_503, sv2v_dc_504, sv2v_dc_505, sv2v_dc_506, sv2v_dc_507, sv2v_dc_508, sv2v_dc_509, sv2v_dc_510, sv2v_dc_511, sv2v_dc_512, sv2v_dc_513, sv2v_dc_514, sv2v_dc_515, sv2v_dc_516, sv2v_dc_517, sv2v_dc_518, sv2v_dc_519, sv2v_dc_520, sv2v_dc_521, sv2v_dc_522, sv2v_dc_523, sv2v_dc_524, sv2v_dc_525, sv2v_dc_526, sv2v_dc_527, sv2v_dc_528, sv2v_dc_529, sv2v_dc_530, sv2v_dc_531, sv2v_dc_532, sv2v_dc_533, sv2v_dc_534, sv2v_dc_535, sv2v_dc_536, sv2v_dc_537, sv2v_dc_538, sv2v_dc_539, sv2v_dc_540, sv2v_dc_541, sv2v_dc_542, sv2v_dc_543, sv2v_dc_544, sv2v_dc_545, sv2v_dc_546, sv2v_dc_547, sv2v_dc_548, sv2v_dc_549, sv2v_dc_550, sv2v_dc_551, sv2v_dc_552, sv2v_dc_553, sv2v_dc_554, sv2v_dc_555, sv2v_dc_556, sv2v_dc_557, sv2v_dc_558, sv2v_dc_559, sv2v_dc_560, sv2v_dc_561, sv2v_dc_562, sv2v_dc_563, sv2v_dc_564, sv2v_dc_565, sv2v_dc_566, sv2v_dc_567, sv2v_dc_568, sv2v_dc_569, sv2v_dc_570, sv2v_dc_571, sv2v_dc_572, sv2v_dc_573, sv2v_dc_574, sv2v_dc_575, sv2v_dc_576, sv2v_dc_577, sv2v_dc_578, sv2v_dc_579, sv2v_dc_580, sv2v_dc_581, sv2v_dc_582, sv2v_dc_583, sv2v_dc_584, sv2v_dc_585, sv2v_dc_586, sv2v_dc_587, sv2v_dc_588, sv2v_dc_589, sv2v_dc_590, sv2v_dc_591, sv2v_dc_592, sv2v_dc_593, sv2v_dc_594, sv2v_dc_595, sv2v_dc_596, sv2v_dc_597, sv2v_dc_598, sv2v_dc_599, sv2v_dc_600, sv2v_dc_601, sv2v_dc_602, sv2v_dc_603, sv2v_dc_604, sv2v_dc_605, sv2v_dc_606, sv2v_dc_607, sv2v_dc_608, sv2v_dc_609, sv2v_dc_610, sv2v_dc_611, sv2v_dc_612, sv2v_dc_613, sv2v_dc_614, sv2v_dc_615, sv2v_dc_616, sv2v_dc_617, sv2v_dc_618, sv2v_dc_619, sv2v_dc_620, sv2v_dc_621, sv2v_dc_622, sv2v_dc_623, sv2v_dc_624, sv2v_dc_625, sv2v_dc_626, sv2v_dc_627, sv2v_dc_628, sv2v_dc_629, sv2v_dc_630, sv2v_dc_631, sv2v_dc_632, sv2v_dc_633, sv2v_dc_634, sv2v_dc_635, sv2v_dc_636, sv2v_dc_637, sv2v_dc_638, sv2v_dc_639, sv2v_dc_640, sv2v_dc_641, sv2v_dc_642, sv2v_dc_643, sv2v_dc_644, sv2v_dc_645, sv2v_dc_646, sv2v_dc_647, sv2v_dc_648, sv2v_dc_649, sv2v_dc_650, sv2v_dc_651, sv2v_dc_652, sv2v_dc_653, sv2v_dc_654, sv2v_dc_655, sv2v_dc_656, sv2v_dc_657, sv2v_dc_658, sv2v_dc_659, sv2v_dc_660, sv2v_dc_661, sv2v_dc_662, sv2v_dc_663, sv2v_dc_664, sv2v_dc_665, sv2v_dc_666, sv2v_dc_667, sv2v_dc_668, sv2v_dc_669, sv2v_dc_670, sv2v_dc_671, sv2v_dc_672, sv2v_dc_673, sv2v_dc_674, sv2v_dc_675, sv2v_dc_676, sv2v_dc_677, sv2v_dc_678, sv2v_dc_679, sv2v_dc_680, sv2v_dc_681, sv2v_dc_682, sv2v_dc_683, sv2v_dc_684, sv2v_dc_685, sv2v_dc_686, sv2v_dc_687, sv2v_dc_688, sv2v_dc_689, sv2v_dc_690, sv2v_dc_691, sv2v_dc_692, sv2v_dc_693, sv2v_dc_694, sv2v_dc_695, sv2v_dc_696, sv2v_dc_697, sv2v_dc_698, sv2v_dc_699, sv2v_dc_700, sv2v_dc_701, sv2v_dc_702, sv2v_dc_703, sv2v_dc_704, sv2v_dc_705, sv2v_dc_706, sv2v_dc_707, sv2v_dc_708, sv2v_dc_709, sv2v_dc_710, sv2v_dc_711, sv2v_dc_712, sv2v_dc_713, sv2v_dc_714, sv2v_dc_715, sv2v_dc_716, sv2v_dc_717, sv2v_dc_718, sv2v_dc_719, sv2v_dc_720, sv2v_dc_721, sv2v_dc_722, sv2v_dc_723, sv2v_dc_724, sv2v_dc_725, sv2v_dc_726, sv2v_dc_727, sv2v_dc_728, sv2v_dc_729, sv2v_dc_730, sv2v_dc_731, sv2v_dc_732, sv2v_dc_733, sv2v_dc_734, sv2v_dc_735, sv2v_dc_736, sv2v_dc_737, sv2v_dc_738, sv2v_dc_739, sv2v_dc_740, sv2v_dc_741, sv2v_dc_742, sv2v_dc_743, sv2v_dc_744, sv2v_dc_745, sv2v_dc_746, sv2v_dc_747, sv2v_dc_748, sv2v_dc_749, sv2v_dc_750, sv2v_dc_751, sv2v_dc_752, sv2v_dc_753, sv2v_dc_754, sv2v_dc_755, sv2v_dc_756, sv2v_dc_757, sv2v_dc_758, sv2v_dc_759, sv2v_dc_760, sv2v_dc_761, sv2v_dc_762, sv2v_dc_763, sv2v_dc_764, sv2v_dc_765, sv2v_dc_766, sv2v_dc_767, sv2v_dc_768, sv2v_dc_769, sv2v_dc_770, sv2v_dc_771, sv2v_dc_772, sv2v_dc_773, sv2v_dc_774, sv2v_dc_775, sv2v_dc_776, sv2v_dc_777, sv2v_dc_778, sv2v_dc_779, sv2v_dc_780, sv2v_dc_781, sv2v_dc_782, sv2v_dc_783, sv2v_dc_784, sv2v_dc_785, sv2v_dc_786, sv2v_dc_787, sv2v_dc_788, sv2v_dc_789, sv2v_dc_790, sv2v_dc_791, sv2v_dc_792, sv2v_dc_793, sv2v_dc_794, sv2v_dc_795, sv2v_dc_796, sv2v_dc_797, sv2v_dc_798, sv2v_dc_799, sv2v_dc_800, sv2v_dc_801, sv2v_dc_802, sv2v_dc_803, sv2v_dc_804, sv2v_dc_805, sv2v_dc_806, sv2v_dc_807, sv2v_dc_808, sv2v_dc_809, sv2v_dc_810, sv2v_dc_811, sv2v_dc_812, sv2v_dc_813, sv2v_dc_814, sv2v_dc_815, sv2v_dc_816, sv2v_dc_817, sv2v_dc_818, sv2v_dc_819, sv2v_dc_820, sv2v_dc_821, sv2v_dc_822, sv2v_dc_823, sv2v_dc_824, sv2v_dc_825, sv2v_dc_826, sv2v_dc_827, sv2v_dc_828, sv2v_dc_829, sv2v_dc_830, sv2v_dc_831, sv2v_dc_832, sv2v_dc_833, sv2v_dc_834, sv2v_dc_835, sv2v_dc_836, sv2v_dc_837, sv2v_dc_838, sv2v_dc_839, sv2v_dc_840, sv2v_dc_841, sv2v_dc_842, sv2v_dc_843, sv2v_dc_844, sv2v_dc_845, sv2v_dc_846, sv2v_dc_847, sv2v_dc_848, sv2v_dc_849, sv2v_dc_850, sv2v_dc_851, sv2v_dc_852, sv2v_dc_853, sv2v_dc_854, sv2v_dc_855, sv2v_dc_856, sv2v_dc_857, sv2v_dc_858, sv2v_dc_859, sv2v_dc_860, sv2v_dc_861, sv2v_dc_862, sv2v_dc_863, sv2v_dc_864, sv2v_dc_865, sv2v_dc_866, sv2v_dc_867, sv2v_dc_868, sv2v_dc_869, sv2v_dc_870, sv2v_dc_871, sv2v_dc_872, sv2v_dc_873, sv2v_dc_874, sv2v_dc_875, sv2v_dc_876, sv2v_dc_877, sv2v_dc_878, sv2v_dc_879, sv2v_dc_880, sv2v_dc_881, sv2v_dc_882, sv2v_dc_883, sv2v_dc_884, sv2v_dc_885, sv2v_dc_886, sv2v_dc_887, sv2v_dc_888, sv2v_dc_889, sv2v_dc_890, sv2v_dc_891, sv2v_dc_892, sv2v_dc_893, sv2v_dc_894, sv2v_dc_895, sv2v_dc_896, sv2v_dc_897, sv2v_dc_898, sv2v_dc_899, sv2v_dc_900, sv2v_dc_901, sv2v_dc_902, sv2v_dc_903, sv2v_dc_904, sv2v_dc_905, sv2v_dc_906, sv2v_dc_907, sv2v_dc_908, sv2v_dc_909, sv2v_dc_910, sv2v_dc_911, sv2v_dc_912, sv2v_dc_913, sv2v_dc_914, sv2v_dc_915, sv2v_dc_916, sv2v_dc_917, sv2v_dc_918, sv2v_dc_919, sv2v_dc_920, sv2v_dc_921, sv2v_dc_922, sv2v_dc_923, sv2v_dc_924, sv2v_dc_925, sv2v_dc_926, sv2v_dc_927, sv2v_dc_928, sv2v_dc_929, sv2v_dc_930, sv2v_dc_931, sv2v_dc_932, sv2v_dc_933, sv2v_dc_934, sv2v_dc_935, sv2v_dc_936, sv2v_dc_937, sv2v_dc_938, sv2v_dc_939, sv2v_dc_940, sv2v_dc_941, sv2v_dc_942, sv2v_dc_943, sv2v_dc_944, sv2v_dc_945, sv2v_dc_946, sv2v_dc_947, sv2v_dc_948, sv2v_dc_949, sv2v_dc_950, sv2v_dc_951, sv2v_dc_952, sv2v_dc_953, sv2v_dc_954, sv2v_dc_955, sv2v_dc_956, sv2v_dc_957, sv2v_dc_958, sv2v_dc_959, sv2v_dc_960, sv2v_dc_961, sv2v_dc_962, sv2v_dc_963, sv2v_dc_964, sv2v_dc_965, sv2v_dc_966, sv2v_dc_967, sv2v_dc_968, sv2v_dc_969, sv2v_dc_970, sv2v_dc_971, sv2v_dc_972, sv2v_dc_973, sv2v_dc_974, sv2v_dc_975, sv2v_dc_976, sv2v_dc_977, sv2v_dc_978, sv2v_dc_979, sv2v_dc_980, sv2v_dc_981, sv2v_dc_982, sv2v_dc_983, sv2v_dc_984, sv2v_dc_985, sv2v_dc_986, sv2v_dc_987, sv2v_dc_988, sv2v_dc_989, sv2v_dc_990, sv2v_dc_991, sv2v_dc_992, sv2v_dc_993, sv2v_dc_994, sv2v_dc_995, sv2v_dc_996, sv2v_dc_997, sv2v_dc_998, sv2v_dc_999, sv2v_dc_1000, sv2v_dc_1001, sv2v_dc_1002, sv2v_dc_1003, sv2v_dc_1004, sv2v_dc_1005, sv2v_dc_1006, sv2v_dc_1007, sv2v_dc_1008, sv2v_dc_1009, sv2v_dc_1010, sv2v_dc_1011, sv2v_dc_1012, sv2v_dc_1013, sv2v_dc_1014, sv2v_dc_1015, sv2v_dc_1016, sv2v_dc_1017, sv2v_dc_1018, sv2v_dc_1019, sv2v_dc_1020, sv2v_dc_1021, sv2v_dc_1022, sv2v_dc_1023, sv2v_dc_1024, sv2v_dc_1025, sv2v_dc_1026, sv2v_dc_1027, sv2v_dc_1028, sv2v_dc_1029, sv2v_dc_1030, sv2v_dc_1031, sv2v_dc_1032, sv2v_dc_1033, sv2v_dc_1034, sv2v_dc_1035, sv2v_dc_1036, sv2v_dc_1037, sv2v_dc_1038, sv2v_dc_1039, sv2v_dc_1040, sv2v_dc_1041, sv2v_dc_1042, sv2v_dc_1043, sv2v_dc_1044, sv2v_dc_1045, sv2v_dc_1046, sv2v_dc_1047, sv2v_dc_1048, sv2v_dc_1049, sv2v_dc_1050, sv2v_dc_1051, sv2v_dc_1052, sv2v_dc_1053, sv2v_dc_1054, sv2v_dc_1055, sv2v_dc_1056, sv2v_dc_1057, sv2v_dc_1058, sv2v_dc_1059, sv2v_dc_1060, sv2v_dc_1061, sv2v_dc_1062, sv2v_dc_1063, sv2v_dc_1064, sv2v_dc_1065, sv2v_dc_1066, sv2v_dc_1067, sv2v_dc_1068, sv2v_dc_1069, sv2v_dc_1070, sv2v_dc_1071, sv2v_dc_1072, sv2v_dc_1073, sv2v_dc_1074, sv2v_dc_1075, sv2v_dc_1076, sv2v_dc_1077, sv2v_dc_1078, sv2v_dc_1079, sv2v_dc_1080, sv2v_dc_1081, sv2v_dc_1082, sv2v_dc_1083, sv2v_dc_1084, sv2v_dc_1085, sv2v_dc_1086, sv2v_dc_1087, sv2v_dc_1088, sv2v_dc_1089, sv2v_dc_1090, sv2v_dc_1091, sv2v_dc_1092, sv2v_dc_1093, sv2v_dc_1094, sv2v_dc_1095, sv2v_dc_1096, sv2v_dc_1097, sv2v_dc_1098, sv2v_dc_1099, sv2v_dc_1100, sv2v_dc_1101, sv2v_dc_1102, sv2v_dc_1103, sv2v_dc_1104, sv2v_dc_1105, sv2v_dc_1106, sv2v_dc_1107, sv2v_dc_1108, sv2v_dc_1109, sv2v_dc_1110, sv2v_dc_1111, sv2v_dc_1112, sv2v_dc_1113, sv2v_dc_1114, sv2v_dc_1115, sv2v_dc_1116, sv2v_dc_1117, sv2v_dc_1118, sv2v_dc_1119, sv2v_dc_1120, sv2v_dc_1121, sv2v_dc_1122, sv2v_dc_1123, sv2v_dc_1124, sv2v_dc_1125, sv2v_dc_1126, sv2v_dc_1127, sv2v_dc_1128, sv2v_dc_1129, sv2v_dc_1130, sv2v_dc_1131, sv2v_dc_1132, sv2v_dc_1133, sv2v_dc_1134, sv2v_dc_1135, sv2v_dc_1136, sv2v_dc_1137, sv2v_dc_1138, sv2v_dc_1139, sv2v_dc_1140, sv2v_dc_1141, sv2v_dc_1142, sv2v_dc_1143, sv2v_dc_1144, sv2v_dc_1145, sv2v_dc_1146, sv2v_dc_1147, sv2v_dc_1148, sv2v_dc_1149, sv2v_dc_1150, sv2v_dc_1151, sv2v_dc_1152, sv2v_dc_1153, sv2v_dc_1154, sv2v_dc_1155, sv2v_dc_1156, sv2v_dc_1157, sv2v_dc_1158, sv2v_dc_1159, sv2v_dc_1160, sv2v_dc_1161, sv2v_dc_1162, sv2v_dc_1163, sv2v_dc_1164, sv2v_dc_1165, sv2v_dc_1166, sv2v_dc_1167, sv2v_dc_1168, sv2v_dc_1169, sv2v_dc_1170, sv2v_dc_1171, sv2v_dc_1172, sv2v_dc_1173, sv2v_dc_1174, sv2v_dc_1175, sv2v_dc_1176, sv2v_dc_1177, sv2v_dc_1178, sv2v_dc_1179, sv2v_dc_1180, sv2v_dc_1181, sv2v_dc_1182, sv2v_dc_1183, sv2v_dc_1184, sv2v_dc_1185, sv2v_dc_1186, sv2v_dc_1187, sv2v_dc_1188, sv2v_dc_1189, sv2v_dc_1190, sv2v_dc_1191, sv2v_dc_1192, sv2v_dc_1193, sv2v_dc_1194, sv2v_dc_1195, sv2v_dc_1196, sv2v_dc_1197, sv2v_dc_1198, sv2v_dc_1199, sv2v_dc_1200, sv2v_dc_1201, sv2v_dc_1202, sv2v_dc_1203, sv2v_dc_1204, sv2v_dc_1205, sv2v_dc_1206, sv2v_dc_1207, sv2v_dc_1208, sv2v_dc_1209, sv2v_dc_1210, sv2v_dc_1211, sv2v_dc_1212, sv2v_dc_1213, sv2v_dc_1214, sv2v_dc_1215, sv2v_dc_1216, sv2v_dc_1217, sv2v_dc_1218, sv2v_dc_1219, sv2v_dc_1220, sv2v_dc_1221, sv2v_dc_1222, sv2v_dc_1223, sv2v_dc_1224, sv2v_dc_1225, sv2v_dc_1226, sv2v_dc_1227, sv2v_dc_1228, sv2v_dc_1229, sv2v_dc_1230, sv2v_dc_1231, sv2v_dc_1232, sv2v_dc_1233, sv2v_dc_1234, sv2v_dc_1235, sv2v_dc_1236, sv2v_dc_1237, sv2v_dc_1238, sv2v_dc_1239, sv2v_dc_1240, sv2v_dc_1241, sv2v_dc_1242, sv2v_dc_1243, sv2v_dc_1244, sv2v_dc_1245, sv2v_dc_1246, sv2v_dc_1247, sv2v_dc_1248, sv2v_dc_1249, sv2v_dc_1250, sv2v_dc_1251, sv2v_dc_1252, sv2v_dc_1253, sv2v_dc_1254, sv2v_dc_1255, sv2v_dc_1256, sv2v_dc_1257, sv2v_dc_1258, sv2v_dc_1259, sv2v_dc_1260, sv2v_dc_1261, sv2v_dc_1262, sv2v_dc_1263, sv2v_dc_1264, sv2v_dc_1265, sv2v_dc_1266, sv2v_dc_1267, sv2v_dc_1268, sv2v_dc_1269, sv2v_dc_1270, sv2v_dc_1271, sv2v_dc_1272, sv2v_dc_1273, sv2v_dc_1274, sv2v_dc_1275, sv2v_dc_1276, sv2v_dc_1277, sv2v_dc_1278, sv2v_dc_1279, sv2v_dc_1280, sv2v_dc_1281, sv2v_dc_1282, sv2v_dc_1283, sv2v_dc_1284, sv2v_dc_1285, sv2v_dc_1286, sv2v_dc_1287, sv2v_dc_1288, sv2v_dc_1289, sv2v_dc_1290, sv2v_dc_1291, sv2v_dc_1292, sv2v_dc_1293, sv2v_dc_1294, sv2v_dc_1295, sv2v_dc_1296, sv2v_dc_1297, sv2v_dc_1298, sv2v_dc_1299, sv2v_dc_1300, sv2v_dc_1301, sv2v_dc_1302, sv2v_dc_1303, sv2v_dc_1304, sv2v_dc_1305, sv2v_dc_1306, sv2v_dc_1307, sv2v_dc_1308, sv2v_dc_1309, sv2v_dc_1310, sv2v_dc_1311, sv2v_dc_1312, sv2v_dc_1313, sv2v_dc_1314, sv2v_dc_1315, sv2v_dc_1316, sv2v_dc_1317, sv2v_dc_1318, sv2v_dc_1319, sv2v_dc_1320, sv2v_dc_1321, sv2v_dc_1322, sv2v_dc_1323, sv2v_dc_1324, sv2v_dc_1325, sv2v_dc_1326, sv2v_dc_1327, sv2v_dc_1328, sv2v_dc_1329, sv2v_dc_1330, sv2v_dc_1331, sv2v_dc_1332, sv2v_dc_1333, sv2v_dc_1334, sv2v_dc_1335, sv2v_dc_1336, sv2v_dc_1337, sv2v_dc_1338, sv2v_dc_1339, sv2v_dc_1340, sv2v_dc_1341, sv2v_dc_1342, sv2v_dc_1343, sv2v_dc_1344, sv2v_dc_1345, sv2v_dc_1346, sv2v_dc_1347, sv2v_dc_1348, sv2v_dc_1349, sv2v_dc_1350, sv2v_dc_1351, sv2v_dc_1352, sv2v_dc_1353, sv2v_dc_1354, sv2v_dc_1355, sv2v_dc_1356, sv2v_dc_1357, sv2v_dc_1358, sv2v_dc_1359, sv2v_dc_1360, sv2v_dc_1361, sv2v_dc_1362, sv2v_dc_1363, sv2v_dc_1364, sv2v_dc_1365, sv2v_dc_1366, sv2v_dc_1367, sv2v_dc_1368, sv2v_dc_1369, sv2v_dc_1370, sv2v_dc_1371, sv2v_dc_1372, sv2v_dc_1373, sv2v_dc_1374, sv2v_dc_1375, sv2v_dc_1376, sv2v_dc_1377, sv2v_dc_1378, sv2v_dc_1379, sv2v_dc_1380, sv2v_dc_1381, sv2v_dc_1382, sv2v_dc_1383, sv2v_dc_1384, sv2v_dc_1385, sv2v_dc_1386, sv2v_dc_1387, sv2v_dc_1388, sv2v_dc_1389, sv2v_dc_1390, sv2v_dc_1391, sv2v_dc_1392, sv2v_dc_1393, sv2v_dc_1394, sv2v_dc_1395, sv2v_dc_1396, sv2v_dc_1397, sv2v_dc_1398, sv2v_dc_1399, sv2v_dc_1400, sv2v_dc_1401, sv2v_dc_1402, sv2v_dc_1403, sv2v_dc_1404, sv2v_dc_1405, sv2v_dc_1406, sv2v_dc_1407, sv2v_dc_1408, sv2v_dc_1409, sv2v_dc_1410, sv2v_dc_1411, sv2v_dc_1412, sv2v_dc_1413, sv2v_dc_1414, sv2v_dc_1415, sv2v_dc_1416, sv2v_dc_1417, sv2v_dc_1418, sv2v_dc_1419, sv2v_dc_1420, sv2v_dc_1421, sv2v_dc_1422, sv2v_dc_1423, sv2v_dc_1424, sv2v_dc_1425, sv2v_dc_1426, sv2v_dc_1427, sv2v_dc_1428, sv2v_dc_1429, sv2v_dc_1430, sv2v_dc_1431, sv2v_dc_1432, sv2v_dc_1433, sv2v_dc_1434, sv2v_dc_1435, sv2v_dc_1436, sv2v_dc_1437, sv2v_dc_1438, sv2v_dc_1439, sv2v_dc_1440, sv2v_dc_1441, sv2v_dc_1442, sv2v_dc_1443, sv2v_dc_1444, sv2v_dc_1445, sv2v_dc_1446, sv2v_dc_1447, sv2v_dc_1448, sv2v_dc_1449, sv2v_dc_1450, sv2v_dc_1451, sv2v_dc_1452, sv2v_dc_1453, sv2v_dc_1454, sv2v_dc_1455, sv2v_dc_1456, sv2v_dc_1457, sv2v_dc_1458, sv2v_dc_1459, sv2v_dc_1460, sv2v_dc_1461, sv2v_dc_1462, sv2v_dc_1463, sv2v_dc_1464, sv2v_dc_1465, sv2v_dc_1466, sv2v_dc_1467, sv2v_dc_1468, sv2v_dc_1469, sv2v_dc_1470, sv2v_dc_1471, sv2v_dc_1472, sv2v_dc_1473, sv2v_dc_1474, sv2v_dc_1475, sv2v_dc_1476, sv2v_dc_1477, sv2v_dc_1478, sv2v_dc_1479, sv2v_dc_1480, sv2v_dc_1481, sv2v_dc_1482, sv2v_dc_1483, sv2v_dc_1484, sv2v_dc_1485, sv2v_dc_1486, sv2v_dc_1487, sv2v_dc_1488, sv2v_dc_1489, sv2v_dc_1490, sv2v_dc_1491, sv2v_dc_1492, sv2v_dc_1493, sv2v_dc_1494, sv2v_dc_1495, sv2v_dc_1496, sv2v_dc_1497, sv2v_dc_1498, sv2v_dc_1499, sv2v_dc_1500, sv2v_dc_1501, sv2v_dc_1502, sv2v_dc_1503, sv2v_dc_1504, sv2v_dc_1505, sv2v_dc_1506, sv2v_dc_1507, sv2v_dc_1508, sv2v_dc_1509, sv2v_dc_1510, sv2v_dc_1511, sv2v_dc_1512, sv2v_dc_1513, sv2v_dc_1514, sv2v_dc_1515, sv2v_dc_1516, sv2v_dc_1517, sv2v_dc_1518, sv2v_dc_1519, sv2v_dc_1520, sv2v_dc_1521, sv2v_dc_1522, sv2v_dc_1523, sv2v_dc_1524, sv2v_dc_1525, sv2v_dc_1526, sv2v_dc_1527, sv2v_dc_1528, sv2v_dc_1529, sv2v_dc_1530, sv2v_dc_1531, sv2v_dc_1532, sv2v_dc_1533, sv2v_dc_1534, sv2v_dc_1535, sv2v_dc_1536, sv2v_dc_1537, sv2v_dc_1538, sv2v_dc_1539, sv2v_dc_1540, sv2v_dc_1541, sv2v_dc_1542, sv2v_dc_1543, sv2v_dc_1544, sv2v_dc_1545, sv2v_dc_1546, sv2v_dc_1547, sv2v_dc_1548, sv2v_dc_1549, sv2v_dc_1550, sv2v_dc_1551, sv2v_dc_1552, sv2v_dc_1553, sv2v_dc_1554, sv2v_dc_1555, sv2v_dc_1556, sv2v_dc_1557, sv2v_dc_1558, sv2v_dc_1559, sv2v_dc_1560, sv2v_dc_1561, sv2v_dc_1562, sv2v_dc_1563, sv2v_dc_1564, sv2v_dc_1565, sv2v_dc_1566, sv2v_dc_1567, sv2v_dc_1568, sv2v_dc_1569, sv2v_dc_1570, sv2v_dc_1571, sv2v_dc_1572, sv2v_dc_1573, sv2v_dc_1574, sv2v_dc_1575, sv2v_dc_1576, sv2v_dc_1577, sv2v_dc_1578, sv2v_dc_1579, sv2v_dc_1580, sv2v_dc_1581, sv2v_dc_1582, sv2v_dc_1583, sv2v_dc_1584, sv2v_dc_1585, sv2v_dc_1586, sv2v_dc_1587, sv2v_dc_1588, sv2v_dc_1589, sv2v_dc_1590, sv2v_dc_1591, sv2v_dc_1592, sv2v_dc_1593, sv2v_dc_1594, sv2v_dc_1595, sv2v_dc_1596, sv2v_dc_1597, sv2v_dc_1598, sv2v_dc_1599, sv2v_dc_1600, sv2v_dc_1601, sv2v_dc_1602, sv2v_dc_1603, sv2v_dc_1604, sv2v_dc_1605, sv2v_dc_1606, sv2v_dc_1607, sv2v_dc_1608, sv2v_dc_1609, sv2v_dc_1610, sv2v_dc_1611, sv2v_dc_1612, sv2v_dc_1613, sv2v_dc_1614, sv2v_dc_1615, sv2v_dc_1616, sv2v_dc_1617, sv2v_dc_1618, sv2v_dc_1619, sv2v_dc_1620, sv2v_dc_1621, sv2v_dc_1622, sv2v_dc_1623, sv2v_dc_1624, sv2v_dc_1625, sv2v_dc_1626, sv2v_dc_1627, sv2v_dc_1628, sv2v_dc_1629, sv2v_dc_1630, sv2v_dc_1631, sv2v_dc_1632, sv2v_dc_1633, sv2v_dc_1634, sv2v_dc_1635, sv2v_dc_1636, sv2v_dc_1637, sv2v_dc_1638, sv2v_dc_1639, sv2v_dc_1640, sv2v_dc_1641, sv2v_dc_1642, sv2v_dc_1643, sv2v_dc_1644, sv2v_dc_1645, sv2v_dc_1646, sv2v_dc_1647, sv2v_dc_1648, sv2v_dc_1649, sv2v_dc_1650, sv2v_dc_1651, sv2v_dc_1652, sv2v_dc_1653, sv2v_dc_1654, sv2v_dc_1655, sv2v_dc_1656, sv2v_dc_1657, sv2v_dc_1658, sv2v_dc_1659, sv2v_dc_1660, sv2v_dc_1661, sv2v_dc_1662, sv2v_dc_1663, sv2v_dc_1664, sv2v_dc_1665, sv2v_dc_1666, sv2v_dc_1667, sv2v_dc_1668, sv2v_dc_1669, sv2v_dc_1670, sv2v_dc_1671, sv2v_dc_1672, sv2v_dc_1673, sv2v_dc_1674, sv2v_dc_1675, sv2v_dc_1676, sv2v_dc_1677, sv2v_dc_1678, sv2v_dc_1679, sv2v_dc_1680, sv2v_dc_1681, sv2v_dc_1682, sv2v_dc_1683, sv2v_dc_1684, sv2v_dc_1685, sv2v_dc_1686, sv2v_dc_1687, sv2v_dc_1688, sv2v_dc_1689, sv2v_dc_1690, sv2v_dc_1691, sv2v_dc_1692, sv2v_dc_1693, sv2v_dc_1694, sv2v_dc_1695, sv2v_dc_1696, sv2v_dc_1697, sv2v_dc_1698, sv2v_dc_1699, sv2v_dc_1700, sv2v_dc_1701, sv2v_dc_1702, sv2v_dc_1703, sv2v_dc_1704, sv2v_dc_1705, sv2v_dc_1706, sv2v_dc_1707, sv2v_dc_1708, sv2v_dc_1709, sv2v_dc_1710, sv2v_dc_1711, sv2v_dc_1712, sv2v_dc_1713, sv2v_dc_1714, sv2v_dc_1715, sv2v_dc_1716, sv2v_dc_1717, sv2v_dc_1718, sv2v_dc_1719, sv2v_dc_1720, sv2v_dc_1721, sv2v_dc_1722, sv2v_dc_1723, sv2v_dc_1724, sv2v_dc_1725, sv2v_dc_1726, sv2v_dc_1727, sv2v_dc_1728, sv2v_dc_1729, sv2v_dc_1730, sv2v_dc_1731, sv2v_dc_1732, sv2v_dc_1733, sv2v_dc_1734, sv2v_dc_1735, sv2v_dc_1736, sv2v_dc_1737, sv2v_dc_1738, sv2v_dc_1739, sv2v_dc_1740, sv2v_dc_1741, sv2v_dc_1742, sv2v_dc_1743, sv2v_dc_1744, sv2v_dc_1745, sv2v_dc_1746, sv2v_dc_1747, sv2v_dc_1748, sv2v_dc_1749, sv2v_dc_1750, sv2v_dc_1751, sv2v_dc_1752, sv2v_dc_1753, sv2v_dc_1754, sv2v_dc_1755, sv2v_dc_1756, sv2v_dc_1757, sv2v_dc_1758, sv2v_dc_1759, sv2v_dc_1760, sv2v_dc_1761, sv2v_dc_1762, sv2v_dc_1763, sv2v_dc_1764, sv2v_dc_1765, sv2v_dc_1766, sv2v_dc_1767, sv2v_dc_1768, sv2v_dc_1769, sv2v_dc_1770, sv2v_dc_1771, sv2v_dc_1772, sv2v_dc_1773, sv2v_dc_1774, sv2v_dc_1775, sv2v_dc_1776, sv2v_dc_1777, sv2v_dc_1778, sv2v_dc_1779, sv2v_dc_1780, sv2v_dc_1781, sv2v_dc_1782, sv2v_dc_1783, sv2v_dc_1784, sv2v_dc_1785, sv2v_dc_1786, sv2v_dc_1787, sv2v_dc_1788, sv2v_dc_1789, sv2v_dc_1790, sv2v_dc_1791, sv2v_dc_1792, sv2v_dc_1793, sv2v_dc_1794, sv2v_dc_1795, sv2v_dc_1796, sv2v_dc_1797, sv2v_dc_1798, sv2v_dc_1799, sv2v_dc_1800, sv2v_dc_1801, sv2v_dc_1802, sv2v_dc_1803, sv2v_dc_1804, sv2v_dc_1805, sv2v_dc_1806, sv2v_dc_1807, sv2v_dc_1808, sv2v_dc_1809, sv2v_dc_1810, sv2v_dc_1811, sv2v_dc_1812, sv2v_dc_1813, sv2v_dc_1814, sv2v_dc_1815, sv2v_dc_1816, sv2v_dc_1817, sv2v_dc_1818, sv2v_dc_1819, sv2v_dc_1820, sv2v_dc_1821, sv2v_dc_1822, sv2v_dc_1823, sv2v_dc_1824, sv2v_dc_1825, sv2v_dc_1826, sv2v_dc_1827, sv2v_dc_1828, sv2v_dc_1829, sv2v_dc_1830, sv2v_dc_1831, sv2v_dc_1832, sv2v_dc_1833, sv2v_dc_1834, sv2v_dc_1835, sv2v_dc_1836, sv2v_dc_1837, sv2v_dc_1838, sv2v_dc_1839, sv2v_dc_1840, sv2v_dc_1841, sv2v_dc_1842, sv2v_dc_1843, sv2v_dc_1844, sv2v_dc_1845, sv2v_dc_1846, sv2v_dc_1847, sv2v_dc_1848, sv2v_dc_1849, sv2v_dc_1850, sv2v_dc_1851, sv2v_dc_1852, sv2v_dc_1853, sv2v_dc_1854, sv2v_dc_1855, sv2v_dc_1856, sv2v_dc_1857, sv2v_dc_1858, sv2v_dc_1859, sv2v_dc_1860, sv2v_dc_1861, sv2v_dc_1862, sv2v_dc_1863, sv2v_dc_1864, sv2v_dc_1865, sv2v_dc_1866, sv2v_dc_1867, sv2v_dc_1868, sv2v_dc_1869, sv2v_dc_1870, sv2v_dc_1871, sv2v_dc_1872, sv2v_dc_1873, sv2v_dc_1874, sv2v_dc_1875, sv2v_dc_1876, sv2v_dc_1877, sv2v_dc_1878, sv2v_dc_1879, sv2v_dc_1880, sv2v_dc_1881, sv2v_dc_1882, sv2v_dc_1883, sv2v_dc_1884, sv2v_dc_1885, sv2v_dc_1886, sv2v_dc_1887, sv2v_dc_1888, sv2v_dc_1889, sv2v_dc_1890, sv2v_dc_1891, sv2v_dc_1892, sv2v_dc_1893, sv2v_dc_1894, sv2v_dc_1895, sv2v_dc_1896, sv2v_dc_1897, sv2v_dc_1898, sv2v_dc_1899, sv2v_dc_1900, sv2v_dc_1901, sv2v_dc_1902, sv2v_dc_1903, sv2v_dc_1904, sv2v_dc_1905, sv2v_dc_1906, sv2v_dc_1907, sv2v_dc_1908, sv2v_dc_1909, sv2v_dc_1910, sv2v_dc_1911, sv2v_dc_1912, sv2v_dc_1913, sv2v_dc_1914, sv2v_dc_1915, sv2v_dc_1916, sv2v_dc_1917, sv2v_dc_1918, sv2v_dc_1919, sv2v_dc_1920, sv2v_dc_1921, sv2v_dc_1922, sv2v_dc_1923, sv2v_dc_1924, sv2v_dc_1925, sv2v_dc_1926, sv2v_dc_1927, sv2v_dc_1928, sv2v_dc_1929, sv2v_dc_1930, sv2v_dc_1931, sv2v_dc_1932, sv2v_dc_1933, sv2v_dc_1934, sv2v_dc_1935, sv2v_dc_1936, sv2v_dc_1937, sv2v_dc_1938, sv2v_dc_1939, sv2v_dc_1940, sv2v_dc_1941, sv2v_dc_1942, sv2v_dc_1943, sv2v_dc_1944, sv2v_dc_1945, sv2v_dc_1946, sv2v_dc_1947, sv2v_dc_1948, sv2v_dc_1949, sv2v_dc_1950, sv2v_dc_1951, sv2v_dc_1952, sv2v_dc_1953, sv2v_dc_1954, sv2v_dc_1955, sv2v_dc_1956, sv2v_dc_1957, sv2v_dc_1958, sv2v_dc_1959, sv2v_dc_1960, sv2v_dc_1961, sv2v_dc_1962, sv2v_dc_1963, sv2v_dc_1964, sv2v_dc_1965, sv2v_dc_1966, sv2v_dc_1967, sv2v_dc_1968, sv2v_dc_1969, sv2v_dc_1970, sv2v_dc_1971, sv2v_dc_1972, sv2v_dc_1973, sv2v_dc_1974, sv2v_dc_1975, sv2v_dc_1976, sv2v_dc_1977, sv2v_dc_1978, sv2v_dc_1979, sv2v_dc_1980, sv2v_dc_1981, sv2v_dc_1982, sv2v_dc_1983, sv2v_dc_1984, sv2v_dc_1985, sv2v_dc_1986, sv2v_dc_1987, sv2v_dc_1988, sv2v_dc_1989, sv2v_dc_1990, sv2v_dc_1991, sv2v_dc_1992, sv2v_dc_1993, sv2v_dc_1994, sv2v_dc_1995, sv2v_dc_1996, sv2v_dc_1997, sv2v_dc_1998, sv2v_dc_1999, sv2v_dc_2000, sv2v_dc_2001, sv2v_dc_2002, sv2v_dc_2003, sv2v_dc_2004, sv2v_dc_2005, sv2v_dc_2006, sv2v_dc_2007, sv2v_dc_2008, sv2v_dc_2009, sv2v_dc_2010, sv2v_dc_2011, sv2v_dc_2012, sv2v_dc_2013, sv2v_dc_2014, sv2v_dc_2015, sv2v_dc_2016, sv2v_dc_2017, sv2v_dc_2018, sv2v_dc_2019, sv2v_dc_2020, sv2v_dc_2021, sv2v_dc_2022, sv2v_dc_2023, sv2v_dc_2024, sv2v_dc_2025, sv2v_dc_2026, sv2v_dc_2027, sv2v_dc_2028, sv2v_dc_2029, sv2v_dc_2030, sv2v_dc_2031, sv2v_dc_2032, sv2v_dc_2033, sv2v_dc_2034, sv2v_dc_2035, sv2v_dc_2036, sv2v_dc_2037, sv2v_dc_2038, sv2v_dc_2039, sv2v_dc_2040, sv2v_dc_2041, sv2v_dc_2042, sv2v_dc_2043, sv2v_dc_2044, sv2v_dc_2045, sv2v_dc_2046, sv2v_dc_2047, sv2v_dc_2048, sv2v_dc_2049, sv2v_dc_2050, sv2v_dc_2051, sv2v_dc_2052, sv2v_dc_2053, sv2v_dc_2054, sv2v_dc_2055, sv2v_dc_2056, sv2v_dc_2057, sv2v_dc_2058, sv2v_dc_2059, sv2v_dc_2060, sv2v_dc_2061, sv2v_dc_2062, sv2v_dc_2063, sv2v_dc_2064, sv2v_dc_2065, sv2v_dc_2066, sv2v_dc_2067, sv2v_dc_2068, sv2v_dc_2069, sv2v_dc_2070, sv2v_dc_2071, sv2v_dc_2072, sv2v_dc_2073, sv2v_dc_2074, sv2v_dc_2075, sv2v_dc_2076, sv2v_dc_2077, sv2v_dc_2078, sv2v_dc_2079, sv2v_dc_2080, sv2v_dc_2081, sv2v_dc_2082, sv2v_dc_2083, sv2v_dc_2084, sv2v_dc_2085, sv2v_dc_2086, sv2v_dc_2087, sv2v_dc_2088, sv2v_dc_2089, sv2v_dc_2090, sv2v_dc_2091, sv2v_dc_2092, sv2v_dc_2093, sv2v_dc_2094, sv2v_dc_2095, sv2v_dc_2096, sv2v_dc_2097, sv2v_dc_2098, sv2v_dc_2099, sv2v_dc_2100, sv2v_dc_2101, sv2v_dc_2102, sv2v_dc_2103, sv2v_dc_2104, sv2v_dc_2105, sv2v_dc_2106, sv2v_dc_2107, sv2v_dc_2108, sv2v_dc_2109, sv2v_dc_2110, sv2v_dc_2111, sv2v_dc_2112, sv2v_dc_2113, sv2v_dc_2114, sv2v_dc_2115, sv2v_dc_2116, sv2v_dc_2117, sv2v_dc_2118, sv2v_dc_2119, sv2v_dc_2120, sv2v_dc_2121, sv2v_dc_2122, sv2v_dc_2123, sv2v_dc_2124, sv2v_dc_2125, sv2v_dc_2126, sv2v_dc_2127, sv2v_dc_2128, sv2v_dc_2129, sv2v_dc_2130, sv2v_dc_2131, sv2v_dc_2132, sv2v_dc_2133, sv2v_dc_2134, sv2v_dc_2135, sv2v_dc_2136, sv2v_dc_2137, sv2v_dc_2138, sv2v_dc_2139, sv2v_dc_2140, sv2v_dc_2141, sv2v_dc_2142, sv2v_dc_2143, sv2v_dc_2144, sv2v_dc_2145, sv2v_dc_2146, sv2v_dc_2147, sv2v_dc_2148, sv2v_dc_2149, sv2v_dc_2150, sv2v_dc_2151, sv2v_dc_2152, sv2v_dc_2153, sv2v_dc_2154, sv2v_dc_2155, sv2v_dc_2156, sv2v_dc_2157, sv2v_dc_2158, sv2v_dc_2159, sv2v_dc_2160, sv2v_dc_2161, sv2v_dc_2162, sv2v_dc_2163, sv2v_dc_2164, sv2v_dc_2165, sv2v_dc_2166, sv2v_dc_2167, sv2v_dc_2168, sv2v_dc_2169, sv2v_dc_2170, sv2v_dc_2171, sv2v_dc_2172, sv2v_dc_2173, sv2v_dc_2174, sv2v_dc_2175, sv2v_dc_2176, sv2v_dc_2177, sv2v_dc_2178, sv2v_dc_2179, sv2v_dc_2180, sv2v_dc_2181, sv2v_dc_2182, sv2v_dc_2183, sv2v_dc_2184, sv2v_dc_2185, sv2v_dc_2186, sv2v_dc_2187, sv2v_dc_2188, sv2v_dc_2189, sv2v_dc_2190, sv2v_dc_2191, sv2v_dc_2192, sv2v_dc_2193, sv2v_dc_2194, sv2v_dc_2195, sv2v_dc_2196, sv2v_dc_2197, sv2v_dc_2198, sv2v_dc_2199, sv2v_dc_2200, sv2v_dc_2201, sv2v_dc_2202, sv2v_dc_2203, sv2v_dc_2204, sv2v_dc_2205, sv2v_dc_2206, sv2v_dc_2207, sv2v_dc_2208, sv2v_dc_2209, sv2v_dc_2210, sv2v_dc_2211, sv2v_dc_2212, sv2v_dc_2213, sv2v_dc_2214, sv2v_dc_2215, sv2v_dc_2216, sv2v_dc_2217, sv2v_dc_2218, sv2v_dc_2219, sv2v_dc_2220, sv2v_dc_2221, sv2v_dc_2222, sv2v_dc_2223, sv2v_dc_2224, sv2v_dc_2225, sv2v_dc_2226, sv2v_dc_2227, sv2v_dc_2228, sv2v_dc_2229, sv2v_dc_2230, sv2v_dc_2231, sv2v_dc_2232, sv2v_dc_2233, sv2v_dc_2234, sv2v_dc_2235, sv2v_dc_2236, sv2v_dc_2237, sv2v_dc_2238, sv2v_dc_2239, sv2v_dc_2240, sv2v_dc_2241, sv2v_dc_2242, sv2v_dc_2243, sv2v_dc_2244, sv2v_dc_2245, sv2v_dc_2246, sv2v_dc_2247, sv2v_dc_2248, sv2v_dc_2249, sv2v_dc_2250, sv2v_dc_2251, sv2v_dc_2252, sv2v_dc_2253, sv2v_dc_2254, sv2v_dc_2255, sv2v_dc_2256, sv2v_dc_2257, sv2v_dc_2258, sv2v_dc_2259, sv2v_dc_2260, sv2v_dc_2261, sv2v_dc_2262, sv2v_dc_2263, sv2v_dc_2264, sv2v_dc_2265, sv2v_dc_2266, sv2v_dc_2267, sv2v_dc_2268, sv2v_dc_2269, sv2v_dc_2270, sv2v_dc_2271, sv2v_dc_2272, sv2v_dc_2273, sv2v_dc_2274, sv2v_dc_2275, sv2v_dc_2276, sv2v_dc_2277, sv2v_dc_2278, sv2v_dc_2279, sv2v_dc_2280, sv2v_dc_2281, sv2v_dc_2282, sv2v_dc_2283, sv2v_dc_2284, sv2v_dc_2285, sv2v_dc_2286, sv2v_dc_2287, sv2v_dc_2288, sv2v_dc_2289, sv2v_dc_2290, sv2v_dc_2291, sv2v_dc_2292, sv2v_dc_2293, sv2v_dc_2294, sv2v_dc_2295, sv2v_dc_2296, sv2v_dc_2297, sv2v_dc_2298, sv2v_dc_2299, sv2v_dc_2300, sv2v_dc_2301, sv2v_dc_2302, sv2v_dc_2303, sv2v_dc_2304, sv2v_dc_2305, sv2v_dc_2306, sv2v_dc_2307, sv2v_dc_2308, sv2v_dc_2309, sv2v_dc_2310, sv2v_dc_2311, sv2v_dc_2312, sv2v_dc_2313, sv2v_dc_2314, sv2v_dc_2315, sv2v_dc_2316, sv2v_dc_2317, sv2v_dc_2318, sv2v_dc_2319, sv2v_dc_2320, sv2v_dc_2321, sv2v_dc_2322, sv2v_dc_2323, sv2v_dc_2324, sv2v_dc_2325, sv2v_dc_2326, sv2v_dc_2327, sv2v_dc_2328, sv2v_dc_2329, sv2v_dc_2330, sv2v_dc_2331, sv2v_dc_2332, sv2v_dc_2333, sv2v_dc_2334, sv2v_dc_2335, sv2v_dc_2336, sv2v_dc_2337, sv2v_dc_2338, sv2v_dc_2339, sv2v_dc_2340, sv2v_dc_2341, sv2v_dc_2342, sv2v_dc_2343, sv2v_dc_2344, sv2v_dc_2345, sv2v_dc_2346, sv2v_dc_2347, sv2v_dc_2348, sv2v_dc_2349, sv2v_dc_2350, sv2v_dc_2351, sv2v_dc_2352, sv2v_dc_2353, sv2v_dc_2354, sv2v_dc_2355, sv2v_dc_2356, sv2v_dc_2357, sv2v_dc_2358, sv2v_dc_2359, sv2v_dc_2360, sv2v_dc_2361, sv2v_dc_2362, sv2v_dc_2363, sv2v_dc_2364, sv2v_dc_2365, sv2v_dc_2366, sv2v_dc_2367, sv2v_dc_2368, sv2v_dc_2369, sv2v_dc_2370, sv2v_dc_2371, sv2v_dc_2372, sv2v_dc_2373, sv2v_dc_2374, sv2v_dc_2375, sv2v_dc_2376, sv2v_dc_2377, sv2v_dc_2378, sv2v_dc_2379, sv2v_dc_2380, sv2v_dc_2381, sv2v_dc_2382, sv2v_dc_2383, sv2v_dc_2384, sv2v_dc_2385, sv2v_dc_2386, sv2v_dc_2387, sv2v_dc_2388, sv2v_dc_2389, sv2v_dc_2390, sv2v_dc_2391, sv2v_dc_2392, sv2v_dc_2393, sv2v_dc_2394, sv2v_dc_2395, sv2v_dc_2396, sv2v_dc_2397, sv2v_dc_2398, sv2v_dc_2399, sv2v_dc_2400, sv2v_dc_2401, sv2v_dc_2402, sv2v_dc_2403, sv2v_dc_2404, sv2v_dc_2405, sv2v_dc_2406, sv2v_dc_2407, sv2v_dc_2408, sv2v_dc_2409, sv2v_dc_2410, sv2v_dc_2411, sv2v_dc_2412, sv2v_dc_2413, sv2v_dc_2414, sv2v_dc_2415, sv2v_dc_2416, sv2v_dc_2417, sv2v_dc_2418, sv2v_dc_2419, sv2v_dc_2420, sv2v_dc_2421, sv2v_dc_2422, sv2v_dc_2423, sv2v_dc_2424, sv2v_dc_2425, sv2v_dc_2426, sv2v_dc_2427, sv2v_dc_2428, sv2v_dc_2429, sv2v_dc_2430, sv2v_dc_2431, sv2v_dc_2432, sv2v_dc_2433, sv2v_dc_2434, sv2v_dc_2435, sv2v_dc_2436, sv2v_dc_2437, sv2v_dc_2438, sv2v_dc_2439, sv2v_dc_2440, sv2v_dc_2441, sv2v_dc_2442, sv2v_dc_2443, sv2v_dc_2444, sv2v_dc_2445, sv2v_dc_2446, sv2v_dc_2447, sv2v_dc_2448, sv2v_dc_2449, sv2v_dc_2450, sv2v_dc_2451, sv2v_dc_2452, sv2v_dc_2453, sv2v_dc_2454, sv2v_dc_2455, sv2v_dc_2456, sv2v_dc_2457, sv2v_dc_2458, sv2v_dc_2459, sv2v_dc_2460, sv2v_dc_2461, sv2v_dc_2462, sv2v_dc_2463, sv2v_dc_2464, sv2v_dc_2465, sv2v_dc_2466, sv2v_dc_2467, sv2v_dc_2468, sv2v_dc_2469, sv2v_dc_2470, sv2v_dc_2471, sv2v_dc_2472, sv2v_dc_2473, sv2v_dc_2474, sv2v_dc_2475, sv2v_dc_2476, sv2v_dc_2477, sv2v_dc_2478, sv2v_dc_2479, sv2v_dc_2480, sv2v_dc_2481, sv2v_dc_2482, sv2v_dc_2483, sv2v_dc_2484, sv2v_dc_2485, sv2v_dc_2486, sv2v_dc_2487, sv2v_dc_2488, sv2v_dc_2489, sv2v_dc_2490, sv2v_dc_2491, sv2v_dc_2492, sv2v_dc_2493, sv2v_dc_2494, sv2v_dc_2495, sv2v_dc_2496, sv2v_dc_2497, sv2v_dc_2498, sv2v_dc_2499, sv2v_dc_2500, sv2v_dc_2501, sv2v_dc_2502, sv2v_dc_2503, sv2v_dc_2504, sv2v_dc_2505, sv2v_dc_2506, sv2v_dc_2507, sv2v_dc_2508, sv2v_dc_2509, sv2v_dc_2510, sv2v_dc_2511, sv2v_dc_2512, sv2v_dc_2513, sv2v_dc_2514, sv2v_dc_2515, sv2v_dc_2516, sv2v_dc_2517, sv2v_dc_2518, sv2v_dc_2519, sv2v_dc_2520, sv2v_dc_2521, sv2v_dc_2522, sv2v_dc_2523, sv2v_dc_2524, sv2v_dc_2525, sv2v_dc_2526, sv2v_dc_2527, sv2v_dc_2528, sv2v_dc_2529, sv2v_dc_2530, sv2v_dc_2531, sv2v_dc_2532, sv2v_dc_2533, sv2v_dc_2534, sv2v_dc_2535, sv2v_dc_2536, sv2v_dc_2537, sv2v_dc_2538, sv2v_dc_2539, sv2v_dc_2540, sv2v_dc_2541, sv2v_dc_2542, sv2v_dc_2543, sv2v_dc_2544, sv2v_dc_2545, sv2v_dc_2546, sv2v_dc_2547, sv2v_dc_2548, sv2v_dc_2549, sv2v_dc_2550, sv2v_dc_2551, sv2v_dc_2552, sv2v_dc_2553, sv2v_dc_2554, sv2v_dc_2555, sv2v_dc_2556, sv2v_dc_2557, sv2v_dc_2558, sv2v_dc_2559, sv2v_dc_2560, sv2v_dc_2561, sv2v_dc_2562, sv2v_dc_2563, sv2v_dc_2564, sv2v_dc_2565, sv2v_dc_2566, sv2v_dc_2567, sv2v_dc_2568, sv2v_dc_2569, sv2v_dc_2570, sv2v_dc_2571, sv2v_dc_2572, sv2v_dc_2573, sv2v_dc_2574, sv2v_dc_2575, sv2v_dc_2576, sv2v_dc_2577, sv2v_dc_2578, sv2v_dc_2579, sv2v_dc_2580, sv2v_dc_2581, sv2v_dc_2582, sv2v_dc_2583, sv2v_dc_2584, sv2v_dc_2585, sv2v_dc_2586, sv2v_dc_2587, sv2v_dc_2588, sv2v_dc_2589, sv2v_dc_2590, sv2v_dc_2591, sv2v_dc_2592, sv2v_dc_2593, sv2v_dc_2594, sv2v_dc_2595, sv2v_dc_2596, sv2v_dc_2597, sv2v_dc_2598, sv2v_dc_2599, sv2v_dc_2600, sv2v_dc_2601, sv2v_dc_2602, sv2v_dc_2603, sv2v_dc_2604, sv2v_dc_2605, sv2v_dc_2606, sv2v_dc_2607, sv2v_dc_2608, sv2v_dc_2609, sv2v_dc_2610, sv2v_dc_2611, sv2v_dc_2612, sv2v_dc_2613, sv2v_dc_2614, sv2v_dc_2615, sv2v_dc_2616, sv2v_dc_2617, sv2v_dc_2618, sv2v_dc_2619, sv2v_dc_2620, sv2v_dc_2621, sv2v_dc_2622, sv2v_dc_2623, sv2v_dc_2624, sv2v_dc_2625, sv2v_dc_2626, sv2v_dc_2627, sv2v_dc_2628, sv2v_dc_2629, sv2v_dc_2630, sv2v_dc_2631, sv2v_dc_2632, sv2v_dc_2633, sv2v_dc_2634, sv2v_dc_2635, sv2v_dc_2636, sv2v_dc_2637, sv2v_dc_2638, sv2v_dc_2639, sv2v_dc_2640, sv2v_dc_2641, sv2v_dc_2642, sv2v_dc_2643, sv2v_dc_2644, sv2v_dc_2645, sv2v_dc_2646, sv2v_dc_2647, sv2v_dc_2648, sv2v_dc_2649, sv2v_dc_2650, sv2v_dc_2651, sv2v_dc_2652, sv2v_dc_2653, sv2v_dc_2654, sv2v_dc_2655, sv2v_dc_2656, sv2v_dc_2657, sv2v_dc_2658, sv2v_dc_2659, sv2v_dc_2660, sv2v_dc_2661, sv2v_dc_2662, sv2v_dc_2663, sv2v_dc_2664, sv2v_dc_2665, sv2v_dc_2666, sv2v_dc_2667, sv2v_dc_2668, sv2v_dc_2669, sv2v_dc_2670, sv2v_dc_2671, sv2v_dc_2672, sv2v_dc_2673, sv2v_dc_2674, sv2v_dc_2675, sv2v_dc_2676, sv2v_dc_2677, sv2v_dc_2678, sv2v_dc_2679, sv2v_dc_2680, sv2v_dc_2681, sv2v_dc_2682, sv2v_dc_2683, sv2v_dc_2684, sv2v_dc_2685, sv2v_dc_2686, sv2v_dc_2687, sv2v_dc_2688, sv2v_dc_2689, sv2v_dc_2690, sv2v_dc_2691, sv2v_dc_2692, sv2v_dc_2693, sv2v_dc_2694, sv2v_dc_2695, sv2v_dc_2696, sv2v_dc_2697, sv2v_dc_2698, sv2v_dc_2699, sv2v_dc_2700, sv2v_dc_2701, sv2v_dc_2702, sv2v_dc_2703, sv2v_dc_2704, sv2v_dc_2705, sv2v_dc_2706, sv2v_dc_2707, sv2v_dc_2708, sv2v_dc_2709, sv2v_dc_2710, sv2v_dc_2711, sv2v_dc_2712, sv2v_dc_2713, sv2v_dc_2714, sv2v_dc_2715, sv2v_dc_2716, sv2v_dc_2717, sv2v_dc_2718, sv2v_dc_2719, sv2v_dc_2720, sv2v_dc_2721, sv2v_dc_2722, sv2v_dc_2723, sv2v_dc_2724, sv2v_dc_2725, sv2v_dc_2726, sv2v_dc_2727, sv2v_dc_2728, sv2v_dc_2729, sv2v_dc_2730, sv2v_dc_2731, sv2v_dc_2732, sv2v_dc_2733, sv2v_dc_2734, sv2v_dc_2735, sv2v_dc_2736, sv2v_dc_2737, sv2v_dc_2738, sv2v_dc_2739, sv2v_dc_2740, sv2v_dc_2741, sv2v_dc_2742, sv2v_dc_2743, sv2v_dc_2744, sv2v_dc_2745, sv2v_dc_2746, sv2v_dc_2747, sv2v_dc_2748, sv2v_dc_2749, sv2v_dc_2750, sv2v_dc_2751, sv2v_dc_2752, sv2v_dc_2753, sv2v_dc_2754, sv2v_dc_2755, sv2v_dc_2756, sv2v_dc_2757, sv2v_dc_2758, sv2v_dc_2759, sv2v_dc_2760, sv2v_dc_2761, sv2v_dc_2762, sv2v_dc_2763, sv2v_dc_2764, sv2v_dc_2765, sv2v_dc_2766, sv2v_dc_2767, sv2v_dc_2768, sv2v_dc_2769, sv2v_dc_2770, sv2v_dc_2771, sv2v_dc_2772, sv2v_dc_2773, sv2v_dc_2774, sv2v_dc_2775, sv2v_dc_2776, sv2v_dc_2777, sv2v_dc_2778, sv2v_dc_2779, sv2v_dc_2780, sv2v_dc_2781, sv2v_dc_2782, sv2v_dc_2783, sv2v_dc_2784, sv2v_dc_2785, sv2v_dc_2786, sv2v_dc_2787, sv2v_dc_2788, sv2v_dc_2789, sv2v_dc_2790, sv2v_dc_2791, sv2v_dc_2792, sv2v_dc_2793, sv2v_dc_2794, sv2v_dc_2795, sv2v_dc_2796, sv2v_dc_2797, sv2v_dc_2798, sv2v_dc_2799, sv2v_dc_2800, sv2v_dc_2801, sv2v_dc_2802, sv2v_dc_2803, sv2v_dc_2804, sv2v_dc_2805, sv2v_dc_2806, sv2v_dc_2807, sv2v_dc_2808, sv2v_dc_2809, sv2v_dc_2810, sv2v_dc_2811, sv2v_dc_2812, sv2v_dc_2813, sv2v_dc_2814, sv2v_dc_2815, sv2v_dc_2816, sv2v_dc_2817, sv2v_dc_2818, sv2v_dc_2819, sv2v_dc_2820, sv2v_dc_2821, sv2v_dc_2822, sv2v_dc_2823, sv2v_dc_2824, sv2v_dc_2825, sv2v_dc_2826, sv2v_dc_2827, sv2v_dc_2828, sv2v_dc_2829, sv2v_dc_2830, sv2v_dc_2831, sv2v_dc_2832, sv2v_dc_2833, sv2v_dc_2834, sv2v_dc_2835, sv2v_dc_2836, sv2v_dc_2837, sv2v_dc_2838, sv2v_dc_2839, sv2v_dc_2840, sv2v_dc_2841, sv2v_dc_2842, sv2v_dc_2843, sv2v_dc_2844, sv2v_dc_2845, sv2v_dc_2846, sv2v_dc_2847, sv2v_dc_2848, sv2v_dc_2849, sv2v_dc_2850, sv2v_dc_2851, sv2v_dc_2852, sv2v_dc_2853, sv2v_dc_2854, sv2v_dc_2855, sv2v_dc_2856, sv2v_dc_2857, sv2v_dc_2858, sv2v_dc_2859, sv2v_dc_2860, sv2v_dc_2861, sv2v_dc_2862, sv2v_dc_2863, sv2v_dc_2864, sv2v_dc_2865, sv2v_dc_2866, sv2v_dc_2867, sv2v_dc_2868, sv2v_dc_2869, sv2v_dc_2870, sv2v_dc_2871, sv2v_dc_2872, sv2v_dc_2873, sv2v_dc_2874, sv2v_dc_2875, sv2v_dc_2876, sv2v_dc_2877, sv2v_dc_2878, sv2v_dc_2879, sv2v_dc_2880, sv2v_dc_2881, sv2v_dc_2882, sv2v_dc_2883, sv2v_dc_2884, sv2v_dc_2885, sv2v_dc_2886, sv2v_dc_2887, sv2v_dc_2888, sv2v_dc_2889, sv2v_dc_2890, sv2v_dc_2891, sv2v_dc_2892, sv2v_dc_2893, sv2v_dc_2894, sv2v_dc_2895, sv2v_dc_2896, sv2v_dc_2897, sv2v_dc_2898, sv2v_dc_2899, sv2v_dc_2900, sv2v_dc_2901, sv2v_dc_2902, sv2v_dc_2903, sv2v_dc_2904, sv2v_dc_2905, sv2v_dc_2906, sv2v_dc_2907, sv2v_dc_2908, sv2v_dc_2909, sv2v_dc_2910, sv2v_dc_2911, sv2v_dc_2912, sv2v_dc_2913, sv2v_dc_2914, sv2v_dc_2915, sv2v_dc_2916, sv2v_dc_2917, sv2v_dc_2918, sv2v_dc_2919, sv2v_dc_2920, sv2v_dc_2921, sv2v_dc_2922, sv2v_dc_2923, sv2v_dc_2924, sv2v_dc_2925, sv2v_dc_2926, sv2v_dc_2927, sv2v_dc_2928, sv2v_dc_2929, sv2v_dc_2930, sv2v_dc_2931, sv2v_dc_2932, sv2v_dc_2933, sv2v_dc_2934, sv2v_dc_2935, sv2v_dc_2936, sv2v_dc_2937, sv2v_dc_2938, sv2v_dc_2939, sv2v_dc_2940, sv2v_dc_2941, sv2v_dc_2942, sv2v_dc_2943, sv2v_dc_2944, sv2v_dc_2945, sv2v_dc_2946, sv2v_dc_2947, sv2v_dc_2948, sv2v_dc_2949, sv2v_dc_2950, sv2v_dc_2951, sv2v_dc_2952, sv2v_dc_2953, sv2v_dc_2954, sv2v_dc_2955, sv2v_dc_2956, sv2v_dc_2957, sv2v_dc_2958, sv2v_dc_2959, sv2v_dc_2960, sv2v_dc_2961, sv2v_dc_2962, sv2v_dc_2963, sv2v_dc_2964, sv2v_dc_2965, sv2v_dc_2966, sv2v_dc_2967, sv2v_dc_2968, sv2v_dc_2969, sv2v_dc_2970, sv2v_dc_2971, sv2v_dc_2972, sv2v_dc_2973, sv2v_dc_2974, sv2v_dc_2975, sv2v_dc_2976, sv2v_dc_2977, sv2v_dc_2978, sv2v_dc_2979, sv2v_dc_2980, sv2v_dc_2981, sv2v_dc_2982, sv2v_dc_2983, sv2v_dc_2984, sv2v_dc_2985, sv2v_dc_2986, sv2v_dc_2987, sv2v_dc_2988, sv2v_dc_2989, sv2v_dc_2990, sv2v_dc_2991, sv2v_dc_2992, sv2v_dc_2993, sv2v_dc_2994, sv2v_dc_2995, sv2v_dc_2996, sv2v_dc_2997, sv2v_dc_2998, sv2v_dc_2999, sv2v_dc_3000, sv2v_dc_3001, sv2v_dc_3002, sv2v_dc_3003, sv2v_dc_3004, sv2v_dc_3005, sv2v_dc_3006, sv2v_dc_3007, sv2v_dc_3008, sv2v_dc_3009, sv2v_dc_3010, sv2v_dc_3011, sv2v_dc_3012, sv2v_dc_3013, sv2v_dc_3014, sv2v_dc_3015, sv2v_dc_3016, sv2v_dc_3017, sv2v_dc_3018, sv2v_dc_3019, sv2v_dc_3020, sv2v_dc_3021, sv2v_dc_3022, sv2v_dc_3023, sv2v_dc_3024, sv2v_dc_3025, sv2v_dc_3026, sv2v_dc_3027, sv2v_dc_3028, sv2v_dc_3029, sv2v_dc_3030, sv2v_dc_3031, sv2v_dc_3032, sv2v_dc_3033, sv2v_dc_3034, sv2v_dc_3035, sv2v_dc_3036, sv2v_dc_3037, sv2v_dc_3038, sv2v_dc_3039, sv2v_dc_3040, sv2v_dc_3041, sv2v_dc_3042, sv2v_dc_3043, sv2v_dc_3044, sv2v_dc_3045, sv2v_dc_3046, sv2v_dc_3047, sv2v_dc_3048, sv2v_dc_3049, sv2v_dc_3050, sv2v_dc_3051, sv2v_dc_3052, sv2v_dc_3053, sv2v_dc_3054, sv2v_dc_3055, sv2v_dc_3056, sv2v_dc_3057, sv2v_dc_3058, sv2v_dc_3059, sv2v_dc_3060, sv2v_dc_3061, sv2v_dc_3062, sv2v_dc_3063, sv2v_dc_3064, sv2v_dc_3065, sv2v_dc_3066, sv2v_dc_3067, sv2v_dc_3068, sv2v_dc_3069, sv2v_dc_3070, reverseOut } = $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) >>> { N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11 };
  assign N0 = ~in[11];
  assign N1 = ~in[10];
  assign N2 = ~in[9];
  assign N3 = ~in[8];
  assign N4 = ~in[7];
  assign N5 = ~in[6];
  assign N6 = ~in[5];
  assign N7 = ~in[4];
  assign N8 = ~in[3];
  assign N9 = ~in[2];
  assign N10 = ~in[1];
  assign N11 = ~in[0];

endmodule



module roundAnyRawFNToRecFN_inExpWidth11_inSigWidth55_outExpWidth11_outSigWidth53
(
  control,
  invalidExc,
  infiniteExc,
  in_isNaN,
  in_isInf,
  in_isZero,
  in_sign,
  in_sExp,
  in_sig,
  roundingMode,
  out,
  exceptionFlags
);

  input [0:0] control;
  input [12:0] in_sExp;
  input [55:0] in_sig;
  input [2:0] roundingMode;
  output [64:0] out;
  output [4:0] exceptionFlags;
  input invalidExc;
  input infiniteExc;
  input in_isNaN;
  input in_isInf;
  input in_isZero;
  input in_sign;
  wire [64:0] out;
  wire [4:0] exceptionFlags;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,exceptionFlags_4_,
  exceptionFlags_3_,roundMagUp,isNaNOut,_0_net__11_,\genblk2.roundPosBit ,\genblk2.anyRoundExtra ,
  \genblk2.anyRound ,\genblk2.roundIncr ,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,
  N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,
  N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,
  N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,
  N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,
  N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,
  N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,
  N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,
  N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,
  N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,
  N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,
  N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,
  N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,
  N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,
  N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,
  N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,
  N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,
  N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,
  N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,
  N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,
  N343,N344,N345,N346,common_overflow,common_totalUnderflow,
  \genblk2.unboundedRange_roundPosBit ,\genblk2.unboundedRange_anyRound ,
  \genblk2.unboundedRange_roundIncr ,\genblk2.roundCarry ,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  common_underflow,common_inexact,notNaN_isSpecialInfOut,commonCase,overflow_roundMagUp,
  pegMinNonzeroMagOut,pegMaxFiniteMagOut,notNaN_isInfOut,N356,N357,N358,N359,N360,N361,
  N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,
  N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,
  N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,
  N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,
  N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,
  N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,
  N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,
  N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,
  N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,
  N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,
  N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,
  N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,
  N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,
  N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,
  N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,
  N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,
  N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,
  N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,
  N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,
  N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,
  N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,
  N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
  N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,
  N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,
  N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,
  N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,
  N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,
  N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,
  N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,
  N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,
  N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,
  N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,
  N874;
  wire [53:0] \genblk2.genblk1.roundMask_main ;
  wire [2:2] \genblk2.roundMask ;
  wire [55:0] \genblk2.roundPosMask ;
  wire [54:0] \genblk2.roundedSig ;
  wire [13:0] \genblk2.sRoundedExp ;
  wire [51:0] common_fractOut;
  assign exceptionFlags_4_ = invalidExc;
  assign exceptionFlags[4] = exceptionFlags_4_;
  assign exceptionFlags_3_ = infiniteExc;
  assign exceptionFlags[3] = exceptionFlags_3_;

  lowMaskLoHi_inWidth12_topBound972_bottomBound1026
  \genblk2.genblk1.lowMask_roundMask 
  (
    .in({ _0_net__11_, in_sExp[10:0] }),
    .out(\genblk2.genblk1.roundMask_main )
  );

  assign common_overflow = $signed(\genblk2.sRoundedExp [13:10]) >= $signed({ 1'b0, 1'b1, 1'b1 });
  assign common_totalUnderflow = $signed(\genblk2.sRoundedExp ) < $signed({ 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0 });
  assign N348 = $signed(in_sExp[12:11]) <= $signed(1'b0);
  assign N413 = ~roundingMode[2];
  assign N414 = ~roundingMode[1];
  assign N415 = N414 | N413;
  assign N416 = roundingMode[0] | N415;
  assign N417 = ~N416;
  assign N418 = roundingMode[1] | N413;
  assign N419 = roundingMode[0] | N418;
  assign N420 = ~N419;
  assign N421 = roundingMode[1] | roundingMode[2];
  assign N422 = roundingMode[0] | N421;
  assign N423 = ~N422;
  assign N424 = N414 | roundingMode[2];
  assign N425 = roundingMode[0] | N424;
  assign N426 = ~N425;
  assign N427 = ~roundingMode[0];
  assign N428 = N427 | N424;
  assign N429 = ~N428;
  assign { N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125 } = { N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124 } + 1'b1;
  assign \genblk2.sRoundedExp  = { in_sExp[12:12], in_sExp } + \genblk2.roundedSig [54:53];
  assign { N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17 } = (N0)? { \genblk2.genblk1.roundMask_main [53:1], \genblk2.roundMask [2:2] } : 
                                                                                                                                                                                                                                                                                            (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N15;
  assign { N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237 } = (N1)? \genblk2.roundPosMask [55:1] : 
                                                                                                                                                                                                                                                                                                                                                        (N236)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = N235;
  assign \genblk2.roundedSig  = (N2)? { N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234 } : 
                                (N3)? { N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345 } : 1'b0;
  assign N2 = \genblk2.roundIncr ;
  assign N3 = N14;
  assign common_fractOut = (N4)? \genblk2.roundedSig [52:1] : 
                           (N5)? \genblk2.roundedSig [51:0] : 1'b0;
  assign N4 = in_sig[55];
  assign N5 = N346;
  assign \genblk2.unboundedRange_roundPosBit  = (N4)? in_sig[2] : 
                                                (N5)? in_sig[1] : 1'b0;
  assign \genblk2.roundCarry  = (N4)? \genblk2.roundedSig [54] : 
                                (N5)? \genblk2.roundedSig [53] : 1'b0;
  assign N347 = (N4)? \genblk2.genblk1.roundMask_main [1] : 
                (N5)? \genblk2.roundMask [2] : 1'b0;
  assign N351 = (N6)? N347 : 
                (N7)? 1'b0 : 1'b0;
  assign N6 = N349;
  assign N7 = N350;
  assign N352 = (N4)? \genblk2.genblk1.roundMask_main [2] : 
                (N5)? \genblk2.genblk1.roundMask_main [1] : 1'b0;
  assign N355 = (N8)? N354 : 
                (N9)? 1'b0 : 1'b0;
  assign N8 = control[0];
  assign N9 = N353;
  assign out[64] = (N10)? 1'b0 : 
                   (N11)? in_sign : 1'b0;
  assign N10 = isNaNOut;
  assign N11 = N837;
  assign N359 = (N12)? common_fractOut[51] : 
                (N358)? 1'b0 : 1'b0;
  assign N12 = N357;
  assign { N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362 } = (N13)? common_fractOut[50:0] : 
                                                                                                                                                                                                                                                                                                                                (N361)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = N360;
  assign roundMagUp = N430 | N432;
  assign N430 = N426 & in_sign;
  assign N432 = N429 & N431;
  assign N431 = ~in_sign;
  assign isNaNOut = exceptionFlags_4_ | N434;
  assign N434 = N433 & in_isNaN;
  assign N433 = ~exceptionFlags_3_;
  assign _0_net__11_ = in_sExp[11] | 1'b0;
  assign \genblk2.roundMask [2] = \genblk2.genblk1.roundMask_main [0] | in_sig[55];
  assign \genblk2.roundPosMask [55] = N435 & \genblk2.genblk1.roundMask_main [53];
  assign N435 = ~1'b0;
  assign \genblk2.roundPosMask [54] = N436 & \genblk2.genblk1.roundMask_main [52];
  assign N436 = ~\genblk2.genblk1.roundMask_main [53];
  assign \genblk2.roundPosMask [53] = N437 & \genblk2.genblk1.roundMask_main [51];
  assign N437 = ~\genblk2.genblk1.roundMask_main [52];
  assign \genblk2.roundPosMask [52] = N438 & \genblk2.genblk1.roundMask_main [50];
  assign N438 = ~\genblk2.genblk1.roundMask_main [51];
  assign \genblk2.roundPosMask [51] = N439 & \genblk2.genblk1.roundMask_main [49];
  assign N439 = ~\genblk2.genblk1.roundMask_main [50];
  assign \genblk2.roundPosMask [50] = N440 & \genblk2.genblk1.roundMask_main [48];
  assign N440 = ~\genblk2.genblk1.roundMask_main [49];
  assign \genblk2.roundPosMask [49] = N441 & \genblk2.genblk1.roundMask_main [47];
  assign N441 = ~\genblk2.genblk1.roundMask_main [48];
  assign \genblk2.roundPosMask [48] = N442 & \genblk2.genblk1.roundMask_main [46];
  assign N442 = ~\genblk2.genblk1.roundMask_main [47];
  assign \genblk2.roundPosMask [47] = N443 & \genblk2.genblk1.roundMask_main [45];
  assign N443 = ~\genblk2.genblk1.roundMask_main [46];
  assign \genblk2.roundPosMask [46] = N444 & \genblk2.genblk1.roundMask_main [44];
  assign N444 = ~\genblk2.genblk1.roundMask_main [45];
  assign \genblk2.roundPosMask [45] = N445 & \genblk2.genblk1.roundMask_main [43];
  assign N445 = ~\genblk2.genblk1.roundMask_main [44];
  assign \genblk2.roundPosMask [44] = N446 & \genblk2.genblk1.roundMask_main [42];
  assign N446 = ~\genblk2.genblk1.roundMask_main [43];
  assign \genblk2.roundPosMask [43] = N447 & \genblk2.genblk1.roundMask_main [41];
  assign N447 = ~\genblk2.genblk1.roundMask_main [42];
  assign \genblk2.roundPosMask [42] = N448 & \genblk2.genblk1.roundMask_main [40];
  assign N448 = ~\genblk2.genblk1.roundMask_main [41];
  assign \genblk2.roundPosMask [41] = N449 & \genblk2.genblk1.roundMask_main [39];
  assign N449 = ~\genblk2.genblk1.roundMask_main [40];
  assign \genblk2.roundPosMask [40] = N450 & \genblk2.genblk1.roundMask_main [38];
  assign N450 = ~\genblk2.genblk1.roundMask_main [39];
  assign \genblk2.roundPosMask [39] = N451 & \genblk2.genblk1.roundMask_main [37];
  assign N451 = ~\genblk2.genblk1.roundMask_main [38];
  assign \genblk2.roundPosMask [38] = N452 & \genblk2.genblk1.roundMask_main [36];
  assign N452 = ~\genblk2.genblk1.roundMask_main [37];
  assign \genblk2.roundPosMask [37] = N453 & \genblk2.genblk1.roundMask_main [35];
  assign N453 = ~\genblk2.genblk1.roundMask_main [36];
  assign \genblk2.roundPosMask [36] = N454 & \genblk2.genblk1.roundMask_main [34];
  assign N454 = ~\genblk2.genblk1.roundMask_main [35];
  assign \genblk2.roundPosMask [35] = N455 & \genblk2.genblk1.roundMask_main [33];
  assign N455 = ~\genblk2.genblk1.roundMask_main [34];
  assign \genblk2.roundPosMask [34] = N456 & \genblk2.genblk1.roundMask_main [32];
  assign N456 = ~\genblk2.genblk1.roundMask_main [33];
  assign \genblk2.roundPosMask [33] = N457 & \genblk2.genblk1.roundMask_main [31];
  assign N457 = ~\genblk2.genblk1.roundMask_main [32];
  assign \genblk2.roundPosMask [32] = N458 & \genblk2.genblk1.roundMask_main [30];
  assign N458 = ~\genblk2.genblk1.roundMask_main [31];
  assign \genblk2.roundPosMask [31] = N459 & \genblk2.genblk1.roundMask_main [29];
  assign N459 = ~\genblk2.genblk1.roundMask_main [30];
  assign \genblk2.roundPosMask [30] = N460 & \genblk2.genblk1.roundMask_main [28];
  assign N460 = ~\genblk2.genblk1.roundMask_main [29];
  assign \genblk2.roundPosMask [29] = N461 & \genblk2.genblk1.roundMask_main [27];
  assign N461 = ~\genblk2.genblk1.roundMask_main [28];
  assign \genblk2.roundPosMask [28] = N462 & \genblk2.genblk1.roundMask_main [26];
  assign N462 = ~\genblk2.genblk1.roundMask_main [27];
  assign \genblk2.roundPosMask [27] = N463 & \genblk2.genblk1.roundMask_main [25];
  assign N463 = ~\genblk2.genblk1.roundMask_main [26];
  assign \genblk2.roundPosMask [26] = N464 & \genblk2.genblk1.roundMask_main [24];
  assign N464 = ~\genblk2.genblk1.roundMask_main [25];
  assign \genblk2.roundPosMask [25] = N465 & \genblk2.genblk1.roundMask_main [23];
  assign N465 = ~\genblk2.genblk1.roundMask_main [24];
  assign \genblk2.roundPosMask [24] = N466 & \genblk2.genblk1.roundMask_main [22];
  assign N466 = ~\genblk2.genblk1.roundMask_main [23];
  assign \genblk2.roundPosMask [23] = N467 & \genblk2.genblk1.roundMask_main [21];
  assign N467 = ~\genblk2.genblk1.roundMask_main [22];
  assign \genblk2.roundPosMask [22] = N468 & \genblk2.genblk1.roundMask_main [20];
  assign N468 = ~\genblk2.genblk1.roundMask_main [21];
  assign \genblk2.roundPosMask [21] = N469 & \genblk2.genblk1.roundMask_main [19];
  assign N469 = ~\genblk2.genblk1.roundMask_main [20];
  assign \genblk2.roundPosMask [20] = N470 & \genblk2.genblk1.roundMask_main [18];
  assign N470 = ~\genblk2.genblk1.roundMask_main [19];
  assign \genblk2.roundPosMask [19] = N471 & \genblk2.genblk1.roundMask_main [17];
  assign N471 = ~\genblk2.genblk1.roundMask_main [18];
  assign \genblk2.roundPosMask [18] = N472 & \genblk2.genblk1.roundMask_main [16];
  assign N472 = ~\genblk2.genblk1.roundMask_main [17];
  assign \genblk2.roundPosMask [17] = N473 & \genblk2.genblk1.roundMask_main [15];
  assign N473 = ~\genblk2.genblk1.roundMask_main [16];
  assign \genblk2.roundPosMask [16] = N474 & \genblk2.genblk1.roundMask_main [14];
  assign N474 = ~\genblk2.genblk1.roundMask_main [15];
  assign \genblk2.roundPosMask [15] = N475 & \genblk2.genblk1.roundMask_main [13];
  assign N475 = ~\genblk2.genblk1.roundMask_main [14];
  assign \genblk2.roundPosMask [14] = N476 & \genblk2.genblk1.roundMask_main [12];
  assign N476 = ~\genblk2.genblk1.roundMask_main [13];
  assign \genblk2.roundPosMask [13] = N477 & \genblk2.genblk1.roundMask_main [11];
  assign N477 = ~\genblk2.genblk1.roundMask_main [12];
  assign \genblk2.roundPosMask [12] = N478 & \genblk2.genblk1.roundMask_main [10];
  assign N478 = ~\genblk2.genblk1.roundMask_main [11];
  assign \genblk2.roundPosMask [11] = N479 & \genblk2.genblk1.roundMask_main [9];
  assign N479 = ~\genblk2.genblk1.roundMask_main [10];
  assign \genblk2.roundPosMask [10] = N480 & \genblk2.genblk1.roundMask_main [8];
  assign N480 = ~\genblk2.genblk1.roundMask_main [9];
  assign \genblk2.roundPosMask [9] = N481 & \genblk2.genblk1.roundMask_main [7];
  assign N481 = ~\genblk2.genblk1.roundMask_main [8];
  assign \genblk2.roundPosMask [8] = N482 & \genblk2.genblk1.roundMask_main [6];
  assign N482 = ~\genblk2.genblk1.roundMask_main [7];
  assign \genblk2.roundPosMask [7] = N483 & \genblk2.genblk1.roundMask_main [5];
  assign N483 = ~\genblk2.genblk1.roundMask_main [6];
  assign \genblk2.roundPosMask [6] = N484 & \genblk2.genblk1.roundMask_main [4];
  assign N484 = ~\genblk2.genblk1.roundMask_main [5];
  assign \genblk2.roundPosMask [5] = N485 & \genblk2.genblk1.roundMask_main [3];
  assign N485 = ~\genblk2.genblk1.roundMask_main [4];
  assign \genblk2.roundPosMask [4] = N486 & \genblk2.genblk1.roundMask_main [2];
  assign N486 = ~\genblk2.genblk1.roundMask_main [3];
  assign \genblk2.roundPosMask [3] = N487 & \genblk2.genblk1.roundMask_main [1];
  assign N487 = ~\genblk2.genblk1.roundMask_main [2];
  assign \genblk2.roundPosMask [2] = N488 & \genblk2.roundMask [2];
  assign N488 = ~\genblk2.genblk1.roundMask_main [1];
  assign \genblk2.roundPosMask [1] = N489 & 1'b1;
  assign N489 = ~\genblk2.roundMask [2];
  assign \genblk2.roundPosMask [0] = N490 & 1'b1;
  assign N490 = ~1'b1;
  assign \genblk2.roundPosBit  = N595 | N601;
  assign N595 = N593 | N594;
  assign N593 = N591 | N592;
  assign N591 = N589 | N590;
  assign N589 = N587 | N588;
  assign N587 = N585 | N586;
  assign N585 = N583 | N584;
  assign N583 = N581 | N582;
  assign N581 = N579 | N580;
  assign N579 = N577 | N578;
  assign N577 = N575 | N576;
  assign N575 = N573 | N574;
  assign N573 = N571 | N572;
  assign N571 = N569 | N570;
  assign N569 = N567 | N568;
  assign N567 = N565 | N566;
  assign N565 = N563 | N564;
  assign N563 = N561 | N562;
  assign N561 = N559 | N560;
  assign N559 = N557 | N558;
  assign N557 = N555 | N556;
  assign N555 = N553 | N554;
  assign N553 = N551 | N552;
  assign N551 = N549 | N550;
  assign N549 = N547 | N548;
  assign N547 = N545 | N546;
  assign N545 = N543 | N544;
  assign N543 = N541 | N542;
  assign N541 = N539 | N540;
  assign N539 = N537 | N538;
  assign N537 = N535 | N536;
  assign N535 = N533 | N534;
  assign N533 = N531 | N532;
  assign N531 = N529 | N530;
  assign N529 = N527 | N528;
  assign N527 = N525 | N526;
  assign N525 = N523 | N524;
  assign N523 = N521 | N522;
  assign N521 = N519 | N520;
  assign N519 = N517 | N518;
  assign N517 = N515 | N516;
  assign N515 = N513 | N514;
  assign N513 = N511 | N512;
  assign N511 = N509 | N510;
  assign N509 = N507 | N508;
  assign N507 = N505 | N506;
  assign N505 = N503 | N504;
  assign N503 = N501 | N502;
  assign N501 = N499 | N500;
  assign N499 = N497 | N498;
  assign N497 = N495 | N496;
  assign N495 = N493 | N494;
  assign N493 = N491 | N492;
  assign N491 = in_sig[55] & \genblk2.roundPosMask [55];
  assign N492 = in_sig[54] & \genblk2.roundPosMask [54];
  assign N494 = in_sig[53] & \genblk2.roundPosMask [53];
  assign N496 = in_sig[52] & \genblk2.roundPosMask [52];
  assign N498 = in_sig[51] & \genblk2.roundPosMask [51];
  assign N500 = in_sig[50] & \genblk2.roundPosMask [50];
  assign N502 = in_sig[49] & \genblk2.roundPosMask [49];
  assign N504 = in_sig[48] & \genblk2.roundPosMask [48];
  assign N506 = in_sig[47] & \genblk2.roundPosMask [47];
  assign N508 = in_sig[46] & \genblk2.roundPosMask [46];
  assign N510 = in_sig[45] & \genblk2.roundPosMask [45];
  assign N512 = in_sig[44] & \genblk2.roundPosMask [44];
  assign N514 = in_sig[43] & \genblk2.roundPosMask [43];
  assign N516 = in_sig[42] & \genblk2.roundPosMask [42];
  assign N518 = in_sig[41] & \genblk2.roundPosMask [41];
  assign N520 = in_sig[40] & \genblk2.roundPosMask [40];
  assign N522 = in_sig[39] & \genblk2.roundPosMask [39];
  assign N524 = in_sig[38] & \genblk2.roundPosMask [38];
  assign N526 = in_sig[37] & \genblk2.roundPosMask [37];
  assign N528 = in_sig[36] & \genblk2.roundPosMask [36];
  assign N530 = in_sig[35] & \genblk2.roundPosMask [35];
  assign N532 = in_sig[34] & \genblk2.roundPosMask [34];
  assign N534 = in_sig[33] & \genblk2.roundPosMask [33];
  assign N536 = in_sig[32] & \genblk2.roundPosMask [32];
  assign N538 = in_sig[31] & \genblk2.roundPosMask [31];
  assign N540 = in_sig[30] & \genblk2.roundPosMask [30];
  assign N542 = in_sig[29] & \genblk2.roundPosMask [29];
  assign N544 = in_sig[28] & \genblk2.roundPosMask [28];
  assign N546 = in_sig[27] & \genblk2.roundPosMask [27];
  assign N548 = in_sig[26] & \genblk2.roundPosMask [26];
  assign N550 = in_sig[25] & \genblk2.roundPosMask [25];
  assign N552 = in_sig[24] & \genblk2.roundPosMask [24];
  assign N554 = in_sig[23] & \genblk2.roundPosMask [23];
  assign N556 = in_sig[22] & \genblk2.roundPosMask [22];
  assign N558 = in_sig[21] & \genblk2.roundPosMask [21];
  assign N560 = in_sig[20] & \genblk2.roundPosMask [20];
  assign N562 = in_sig[19] & \genblk2.roundPosMask [19];
  assign N564 = in_sig[18] & \genblk2.roundPosMask [18];
  assign N566 = in_sig[17] & \genblk2.roundPosMask [17];
  assign N568 = in_sig[16] & \genblk2.roundPosMask [16];
  assign N570 = in_sig[15] & \genblk2.roundPosMask [15];
  assign N572 = in_sig[14] & \genblk2.roundPosMask [14];
  assign N574 = in_sig[13] & \genblk2.roundPosMask [13];
  assign N576 = in_sig[12] & \genblk2.roundPosMask [12];
  assign N578 = in_sig[11] & \genblk2.roundPosMask [11];
  assign N580 = in_sig[10] & \genblk2.roundPosMask [10];
  assign N582 = in_sig[9] & \genblk2.roundPosMask [9];
  assign N584 = in_sig[8] & \genblk2.roundPosMask [8];
  assign N586 = in_sig[7] & \genblk2.roundPosMask [7];
  assign N588 = in_sig[6] & \genblk2.roundPosMask [6];
  assign N590 = in_sig[5] & \genblk2.roundPosMask [5];
  assign N592 = in_sig[4] & \genblk2.roundPosMask [4];
  assign N594 = in_sig[3] & \genblk2.roundPosMask [3];
  assign N601 = N600 & N435;
  assign N600 = N598 | N599;
  assign N598 = N596 | N597;
  assign N596 = in_sig[2] & \genblk2.roundPosMask [2];
  assign N597 = in_sig[1] & \genblk2.roundPosMask [1];
  assign N599 = in_sig[0] & \genblk2.roundPosMask [0];
  assign \genblk2.anyRoundExtra  = N706 | N712;
  assign N706 = N704 | N705;
  assign N704 = N702 | N703;
  assign N702 = N700 | N701;
  assign N700 = N698 | N699;
  assign N698 = N696 | N697;
  assign N696 = N694 | N695;
  assign N694 = N692 | N693;
  assign N692 = N690 | N691;
  assign N690 = N688 | N689;
  assign N688 = N686 | N687;
  assign N686 = N684 | N685;
  assign N684 = N682 | N683;
  assign N682 = N680 | N681;
  assign N680 = N678 | N679;
  assign N678 = N676 | N677;
  assign N676 = N674 | N675;
  assign N674 = N672 | N673;
  assign N672 = N670 | N671;
  assign N670 = N668 | N669;
  assign N668 = N666 | N667;
  assign N666 = N664 | N665;
  assign N664 = N662 | N663;
  assign N662 = N660 | N661;
  assign N660 = N658 | N659;
  assign N658 = N656 | N657;
  assign N656 = N654 | N655;
  assign N654 = N652 | N653;
  assign N652 = N650 | N651;
  assign N650 = N648 | N649;
  assign N648 = N646 | N647;
  assign N646 = N644 | N645;
  assign N644 = N642 | N643;
  assign N642 = N640 | N641;
  assign N640 = N638 | N639;
  assign N638 = N636 | N637;
  assign N636 = N634 | N635;
  assign N634 = N632 | N633;
  assign N632 = N630 | N631;
  assign N630 = N628 | N629;
  assign N628 = N626 | N627;
  assign N626 = N624 | N625;
  assign N624 = N622 | N623;
  assign N622 = N620 | N621;
  assign N620 = N618 | N619;
  assign N618 = N616 | N617;
  assign N616 = N614 | N615;
  assign N614 = N612 | N613;
  assign N612 = N610 | N611;
  assign N610 = N608 | N609;
  assign N608 = N606 | N607;
  assign N606 = N604 | N605;
  assign N604 = N602 | N603;
  assign N602 = in_sig[55] & 1'b0;
  assign N603 = in_sig[54] & \genblk2.genblk1.roundMask_main [53];
  assign N605 = in_sig[53] & \genblk2.genblk1.roundMask_main [52];
  assign N607 = in_sig[52] & \genblk2.genblk1.roundMask_main [51];
  assign N609 = in_sig[51] & \genblk2.genblk1.roundMask_main [50];
  assign N611 = in_sig[50] & \genblk2.genblk1.roundMask_main [49];
  assign N613 = in_sig[49] & \genblk2.genblk1.roundMask_main [48];
  assign N615 = in_sig[48] & \genblk2.genblk1.roundMask_main [47];
  assign N617 = in_sig[47] & \genblk2.genblk1.roundMask_main [46];
  assign N619 = in_sig[46] & \genblk2.genblk1.roundMask_main [45];
  assign N621 = in_sig[45] & \genblk2.genblk1.roundMask_main [44];
  assign N623 = in_sig[44] & \genblk2.genblk1.roundMask_main [43];
  assign N625 = in_sig[43] & \genblk2.genblk1.roundMask_main [42];
  assign N627 = in_sig[42] & \genblk2.genblk1.roundMask_main [41];
  assign N629 = in_sig[41] & \genblk2.genblk1.roundMask_main [40];
  assign N631 = in_sig[40] & \genblk2.genblk1.roundMask_main [39];
  assign N633 = in_sig[39] & \genblk2.genblk1.roundMask_main [38];
  assign N635 = in_sig[38] & \genblk2.genblk1.roundMask_main [37];
  assign N637 = in_sig[37] & \genblk2.genblk1.roundMask_main [36];
  assign N639 = in_sig[36] & \genblk2.genblk1.roundMask_main [35];
  assign N641 = in_sig[35] & \genblk2.genblk1.roundMask_main [34];
  assign N643 = in_sig[34] & \genblk2.genblk1.roundMask_main [33];
  assign N645 = in_sig[33] & \genblk2.genblk1.roundMask_main [32];
  assign N647 = in_sig[32] & \genblk2.genblk1.roundMask_main [31];
  assign N649 = in_sig[31] & \genblk2.genblk1.roundMask_main [30];
  assign N651 = in_sig[30] & \genblk2.genblk1.roundMask_main [29];
  assign N653 = in_sig[29] & \genblk2.genblk1.roundMask_main [28];
  assign N655 = in_sig[28] & \genblk2.genblk1.roundMask_main [27];
  assign N657 = in_sig[27] & \genblk2.genblk1.roundMask_main [26];
  assign N659 = in_sig[26] & \genblk2.genblk1.roundMask_main [25];
  assign N661 = in_sig[25] & \genblk2.genblk1.roundMask_main [24];
  assign N663 = in_sig[24] & \genblk2.genblk1.roundMask_main [23];
  assign N665 = in_sig[23] & \genblk2.genblk1.roundMask_main [22];
  assign N667 = in_sig[22] & \genblk2.genblk1.roundMask_main [21];
  assign N669 = in_sig[21] & \genblk2.genblk1.roundMask_main [20];
  assign N671 = in_sig[20] & \genblk2.genblk1.roundMask_main [19];
  assign N673 = in_sig[19] & \genblk2.genblk1.roundMask_main [18];
  assign N675 = in_sig[18] & \genblk2.genblk1.roundMask_main [17];
  assign N677 = in_sig[17] & \genblk2.genblk1.roundMask_main [16];
  assign N679 = in_sig[16] & \genblk2.genblk1.roundMask_main [15];
  assign N681 = in_sig[15] & \genblk2.genblk1.roundMask_main [14];
  assign N683 = in_sig[14] & \genblk2.genblk1.roundMask_main [13];
  assign N685 = in_sig[13] & \genblk2.genblk1.roundMask_main [12];
  assign N687 = in_sig[12] & \genblk2.genblk1.roundMask_main [11];
  assign N689 = in_sig[11] & \genblk2.genblk1.roundMask_main [10];
  assign N691 = in_sig[10] & \genblk2.genblk1.roundMask_main [9];
  assign N693 = in_sig[9] & \genblk2.genblk1.roundMask_main [8];
  assign N695 = in_sig[8] & \genblk2.genblk1.roundMask_main [7];
  assign N697 = in_sig[7] & \genblk2.genblk1.roundMask_main [6];
  assign N699 = in_sig[6] & \genblk2.genblk1.roundMask_main [5];
  assign N701 = in_sig[5] & \genblk2.genblk1.roundMask_main [4];
  assign N703 = in_sig[4] & \genblk2.genblk1.roundMask_main [3];
  assign N705 = in_sig[3] & \genblk2.genblk1.roundMask_main [2];
  assign N712 = N711 & N435;
  assign N711 = N709 | N710;
  assign N709 = N707 | N708;
  assign N707 = in_sig[2] & \genblk2.genblk1.roundMask_main [1];
  assign N708 = in_sig[1] & \genblk2.roundMask [2];
  assign N710 = in_sig[0] & 1'b1;
  assign \genblk2.anyRound  = \genblk2.roundPosBit  | \genblk2.anyRoundExtra ;
  assign \genblk2.roundIncr  = N714 | N715;
  assign N714 = N713 & \genblk2.roundPosBit ;
  assign N713 = N423 | N420;
  assign N715 = roundMagUp & \genblk2.anyRound ;
  assign N14 = ~\genblk2.roundIncr ;
  assign N15 = N716 & N717;
  assign N716 = N423 & \genblk2.roundPosBit ;
  assign N717 = ~\genblk2.anyRoundExtra ;
  assign N16 = ~N15;
  assign N71 = in_sig[55] | \genblk2.genblk1.roundMask_main [53];
  assign N72 = in_sig[54] | \genblk2.genblk1.roundMask_main [52];
  assign N73 = in_sig[53] | \genblk2.genblk1.roundMask_main [51];
  assign N74 = in_sig[52] | \genblk2.genblk1.roundMask_main [50];
  assign N75 = in_sig[51] | \genblk2.genblk1.roundMask_main [49];
  assign N76 = in_sig[50] | \genblk2.genblk1.roundMask_main [48];
  assign N77 = in_sig[49] | \genblk2.genblk1.roundMask_main [47];
  assign N78 = in_sig[48] | \genblk2.genblk1.roundMask_main [46];
  assign N79 = in_sig[47] | \genblk2.genblk1.roundMask_main [45];
  assign N80 = in_sig[46] | \genblk2.genblk1.roundMask_main [44];
  assign N81 = in_sig[45] | \genblk2.genblk1.roundMask_main [43];
  assign N82 = in_sig[44] | \genblk2.genblk1.roundMask_main [42];
  assign N83 = in_sig[43] | \genblk2.genblk1.roundMask_main [41];
  assign N84 = in_sig[42] | \genblk2.genblk1.roundMask_main [40];
  assign N85 = in_sig[41] | \genblk2.genblk1.roundMask_main [39];
  assign N86 = in_sig[40] | \genblk2.genblk1.roundMask_main [38];
  assign N87 = in_sig[39] | \genblk2.genblk1.roundMask_main [37];
  assign N88 = in_sig[38] | \genblk2.genblk1.roundMask_main [36];
  assign N89 = in_sig[37] | \genblk2.genblk1.roundMask_main [35];
  assign N90 = in_sig[36] | \genblk2.genblk1.roundMask_main [34];
  assign N91 = in_sig[35] | \genblk2.genblk1.roundMask_main [33];
  assign N92 = in_sig[34] | \genblk2.genblk1.roundMask_main [32];
  assign N93 = in_sig[33] | \genblk2.genblk1.roundMask_main [31];
  assign N94 = in_sig[32] | \genblk2.genblk1.roundMask_main [30];
  assign N95 = in_sig[31] | \genblk2.genblk1.roundMask_main [29];
  assign N96 = in_sig[30] | \genblk2.genblk1.roundMask_main [28];
  assign N97 = in_sig[29] | \genblk2.genblk1.roundMask_main [27];
  assign N98 = in_sig[28] | \genblk2.genblk1.roundMask_main [26];
  assign N99 = in_sig[27] | \genblk2.genblk1.roundMask_main [25];
  assign N100 = in_sig[26] | \genblk2.genblk1.roundMask_main [24];
  assign N101 = in_sig[25] | \genblk2.genblk1.roundMask_main [23];
  assign N102 = in_sig[24] | \genblk2.genblk1.roundMask_main [22];
  assign N103 = in_sig[23] | \genblk2.genblk1.roundMask_main [21];
  assign N104 = in_sig[22] | \genblk2.genblk1.roundMask_main [20];
  assign N105 = in_sig[21] | \genblk2.genblk1.roundMask_main [19];
  assign N106 = in_sig[20] | \genblk2.genblk1.roundMask_main [18];
  assign N107 = in_sig[19] | \genblk2.genblk1.roundMask_main [17];
  assign N108 = in_sig[18] | \genblk2.genblk1.roundMask_main [16];
  assign N109 = in_sig[17] | \genblk2.genblk1.roundMask_main [15];
  assign N110 = in_sig[16] | \genblk2.genblk1.roundMask_main [14];
  assign N111 = in_sig[15] | \genblk2.genblk1.roundMask_main [13];
  assign N112 = in_sig[14] | \genblk2.genblk1.roundMask_main [12];
  assign N113 = in_sig[13] | \genblk2.genblk1.roundMask_main [11];
  assign N114 = in_sig[12] | \genblk2.genblk1.roundMask_main [10];
  assign N115 = in_sig[11] | \genblk2.genblk1.roundMask_main [9];
  assign N116 = in_sig[10] | \genblk2.genblk1.roundMask_main [8];
  assign N117 = in_sig[9] | \genblk2.genblk1.roundMask_main [7];
  assign N118 = in_sig[8] | \genblk2.genblk1.roundMask_main [6];
  assign N119 = in_sig[7] | \genblk2.genblk1.roundMask_main [5];
  assign N120 = in_sig[6] | \genblk2.genblk1.roundMask_main [4];
  assign N121 = in_sig[5] | \genblk2.genblk1.roundMask_main [3];
  assign N122 = in_sig[4] | \genblk2.genblk1.roundMask_main [2];
  assign N123 = in_sig[3] | \genblk2.genblk1.roundMask_main [1];
  assign N124 = in_sig[2] | \genblk2.roundMask [2];
  assign N180 = N179 & N718;
  assign N718 = ~N70;
  assign N181 = N178 & N719;
  assign N719 = ~N69;
  assign N182 = N177 & N720;
  assign N720 = ~N68;
  assign N183 = N176 & N721;
  assign N721 = ~N67;
  assign N184 = N175 & N722;
  assign N722 = ~N66;
  assign N185 = N174 & N723;
  assign N723 = ~N65;
  assign N186 = N173 & N724;
  assign N724 = ~N64;
  assign N187 = N172 & N725;
  assign N725 = ~N63;
  assign N188 = N171 & N726;
  assign N726 = ~N62;
  assign N189 = N170 & N727;
  assign N727 = ~N61;
  assign N190 = N169 & N728;
  assign N728 = ~N60;
  assign N191 = N168 & N729;
  assign N729 = ~N59;
  assign N192 = N167 & N730;
  assign N730 = ~N58;
  assign N193 = N166 & N731;
  assign N731 = ~N57;
  assign N194 = N165 & N732;
  assign N732 = ~N56;
  assign N195 = N164 & N733;
  assign N733 = ~N55;
  assign N196 = N163 & N734;
  assign N734 = ~N54;
  assign N197 = N162 & N735;
  assign N735 = ~N53;
  assign N198 = N161 & N736;
  assign N736 = ~N52;
  assign N199 = N160 & N737;
  assign N737 = ~N51;
  assign N200 = N159 & N738;
  assign N738 = ~N50;
  assign N201 = N158 & N739;
  assign N739 = ~N49;
  assign N202 = N157 & N740;
  assign N740 = ~N48;
  assign N203 = N156 & N741;
  assign N741 = ~N47;
  assign N204 = N155 & N742;
  assign N742 = ~N46;
  assign N205 = N154 & N743;
  assign N743 = ~N45;
  assign N206 = N153 & N744;
  assign N744 = ~N44;
  assign N207 = N152 & N745;
  assign N745 = ~N43;
  assign N208 = N151 & N746;
  assign N746 = ~N42;
  assign N209 = N150 & N747;
  assign N747 = ~N41;
  assign N210 = N149 & N748;
  assign N748 = ~N40;
  assign N211 = N148 & N749;
  assign N749 = ~N39;
  assign N212 = N147 & N750;
  assign N750 = ~N38;
  assign N213 = N146 & N751;
  assign N751 = ~N37;
  assign N214 = N145 & N752;
  assign N752 = ~N36;
  assign N215 = N144 & N753;
  assign N753 = ~N35;
  assign N216 = N143 & N754;
  assign N754 = ~N34;
  assign N217 = N142 & N755;
  assign N755 = ~N33;
  assign N218 = N141 & N756;
  assign N756 = ~N32;
  assign N219 = N140 & N757;
  assign N757 = ~N31;
  assign N220 = N139 & N758;
  assign N758 = ~N30;
  assign N221 = N138 & N759;
  assign N759 = ~N29;
  assign N222 = N137 & N760;
  assign N760 = ~N28;
  assign N223 = N136 & N761;
  assign N761 = ~N27;
  assign N224 = N135 & N762;
  assign N762 = ~N26;
  assign N225 = N134 & N763;
  assign N763 = ~N25;
  assign N226 = N133 & N764;
  assign N764 = ~N24;
  assign N227 = N132 & N765;
  assign N765 = ~N23;
  assign N228 = N131 & N766;
  assign N766 = ~N22;
  assign N229 = N130 & N767;
  assign N767 = ~N21;
  assign N230 = N129 & N768;
  assign N768 = ~N20;
  assign N231 = N128 & N769;
  assign N769 = ~N19;
  assign N232 = N127 & N770;
  assign N770 = ~N18;
  assign N233 = N126 & N771;
  assign N771 = ~N17;
  assign N234 = N125 & N772;
  assign N772 = ~N15;
  assign N235 = N417 & \genblk2.anyRound ;
  assign N236 = ~N235;
  assign N292 = N773 | N290;
  assign N773 = in_sig[55] & N436;
  assign N293 = N774 | N289;
  assign N774 = in_sig[54] & N437;
  assign N294 = N775 | N288;
  assign N775 = in_sig[53] & N438;
  assign N295 = N776 | N287;
  assign N776 = in_sig[52] & N439;
  assign N296 = N777 | N286;
  assign N777 = in_sig[51] & N440;
  assign N297 = N778 | N285;
  assign N778 = in_sig[50] & N441;
  assign N298 = N779 | N284;
  assign N779 = in_sig[49] & N442;
  assign N299 = N780 | N283;
  assign N780 = in_sig[48] & N443;
  assign N300 = N781 | N282;
  assign N781 = in_sig[47] & N444;
  assign N301 = N782 | N281;
  assign N782 = in_sig[46] & N445;
  assign N302 = N783 | N280;
  assign N783 = in_sig[45] & N446;
  assign N303 = N784 | N279;
  assign N784 = in_sig[44] & N447;
  assign N304 = N785 | N278;
  assign N785 = in_sig[43] & N448;
  assign N305 = N786 | N277;
  assign N786 = in_sig[42] & N449;
  assign N306 = N787 | N276;
  assign N787 = in_sig[41] & N450;
  assign N307 = N788 | N275;
  assign N788 = in_sig[40] & N451;
  assign N308 = N789 | N274;
  assign N789 = in_sig[39] & N452;
  assign N309 = N790 | N273;
  assign N790 = in_sig[38] & N453;
  assign N310 = N791 | N272;
  assign N791 = in_sig[37] & N454;
  assign N311 = N792 | N271;
  assign N792 = in_sig[36] & N455;
  assign N312 = N793 | N270;
  assign N793 = in_sig[35] & N456;
  assign N313 = N794 | N269;
  assign N794 = in_sig[34] & N457;
  assign N314 = N795 | N268;
  assign N795 = in_sig[33] & N458;
  assign N315 = N796 | N267;
  assign N796 = in_sig[32] & N459;
  assign N316 = N797 | N266;
  assign N797 = in_sig[31] & N460;
  assign N317 = N798 | N265;
  assign N798 = in_sig[30] & N461;
  assign N318 = N799 | N264;
  assign N799 = in_sig[29] & N462;
  assign N319 = N800 | N263;
  assign N800 = in_sig[28] & N463;
  assign N320 = N801 | N262;
  assign N801 = in_sig[27] & N464;
  assign N321 = N802 | N261;
  assign N802 = in_sig[26] & N465;
  assign N322 = N803 | N260;
  assign N803 = in_sig[25] & N466;
  assign N323 = N804 | N259;
  assign N804 = in_sig[24] & N467;
  assign N324 = N805 | N258;
  assign N805 = in_sig[23] & N468;
  assign N325 = N806 | N257;
  assign N806 = in_sig[22] & N469;
  assign N326 = N807 | N256;
  assign N807 = in_sig[21] & N470;
  assign N327 = N808 | N255;
  assign N808 = in_sig[20] & N471;
  assign N328 = N809 | N254;
  assign N809 = in_sig[19] & N472;
  assign N329 = N810 | N253;
  assign N810 = in_sig[18] & N473;
  assign N330 = N811 | N252;
  assign N811 = in_sig[17] & N474;
  assign N331 = N812 | N251;
  assign N812 = in_sig[16] & N475;
  assign N332 = N813 | N250;
  assign N813 = in_sig[15] & N476;
  assign N333 = N814 | N249;
  assign N814 = in_sig[14] & N477;
  assign N334 = N815 | N248;
  assign N815 = in_sig[13] & N478;
  assign N335 = N816 | N247;
  assign N816 = in_sig[12] & N479;
  assign N336 = N817 | N246;
  assign N817 = in_sig[11] & N480;
  assign N337 = N818 | N245;
  assign N818 = in_sig[10] & N481;
  assign N338 = N819 | N244;
  assign N819 = in_sig[9] & N482;
  assign N339 = N820 | N243;
  assign N820 = in_sig[8] & N483;
  assign N340 = N821 | N242;
  assign N821 = in_sig[7] & N484;
  assign N341 = N822 | N241;
  assign N822 = in_sig[6] & N485;
  assign N342 = N823 | N240;
  assign N823 = in_sig[5] & N486;
  assign N343 = N824 | N239;
  assign N824 = in_sig[4] & N487;
  assign N344 = N825 | N238;
  assign N825 = in_sig[3] & N488;
  assign N345 = N826 | N237;
  assign N826 = in_sig[2] & N489;
  assign N346 = ~in_sig[55];
  assign \genblk2.unboundedRange_anyRound  = N827 | N828;
  assign N827 = in_sig[55] & in_sig[2];
  assign N828 = in_sig[1] | in_sig[0];
  assign \genblk2.unboundedRange_roundIncr  = N830 | N831;
  assign N830 = N829 & \genblk2.unboundedRange_roundPosBit ;
  assign N829 = N423 | N420;
  assign N831 = roundMagUp & \genblk2.unboundedRange_anyRound ;
  assign N349 = \genblk2.anyRound  & N348;
  assign N350 = ~N349;
  assign N353 = ~control[0];
  assign N354 = ~N352;
  assign common_underflow = common_totalUnderflow | N836;
  assign N836 = N351 & N835;
  assign N835 = ~N834;
  assign N834 = N833 & \genblk2.unboundedRange_roundIncr ;
  assign N833 = N832 & \genblk2.roundPosBit ;
  assign N832 = N355 & \genblk2.roundCarry ;
  assign common_inexact = common_totalUnderflow | \genblk2.anyRound ;
  assign notNaN_isSpecialInfOut = exceptionFlags_3_ | in_isInf;
  assign commonCase = N839 & N840;
  assign N839 = N837 & N838;
  assign N837 = ~isNaNOut;
  assign N838 = ~notNaN_isSpecialInfOut;
  assign N840 = ~in_isZero;
  assign exceptionFlags[2] = commonCase & common_overflow;
  assign exceptionFlags[1] = commonCase & common_underflow;
  assign exceptionFlags[0] = exceptionFlags[2] | N841;
  assign N841 = commonCase & common_inexact;
  assign overflow_roundMagUp = N842 | roundMagUp;
  assign N842 = N423 | N420;
  assign pegMinNonzeroMagOut = N843 & N844;
  assign N843 = commonCase & common_totalUnderflow;
  assign N844 = roundMagUp | N417;
  assign pegMaxFiniteMagOut = exceptionFlags[2] & N845;
  assign N845 = ~overflow_roundMagUp;
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | N846;
  assign N846 = exceptionFlags[2] & overflow_roundMagUp;
  assign N356 = in_isZero | common_totalUnderflow;
  assign out[63] = N852 | isNaNOut;
  assign N852 = N851 | notNaN_isInfOut;
  assign N851 = N850 | pegMaxFiniteMagOut;
  assign N850 = N848 & N849;
  assign N848 = \genblk2.sRoundedExp [11] & N847;
  assign N847 = ~N356;
  assign N849 = ~pegMinNonzeroMagOut;
  assign out[62] = N857 | isNaNOut;
  assign N857 = N856 | notNaN_isInfOut;
  assign N856 = N854 & N855;
  assign N854 = N853 & N849;
  assign N853 = \genblk2.sRoundedExp [10] & N847;
  assign N855 = ~pegMaxFiniteMagOut;
  assign out[61] = N862 | isNaNOut;
  assign N862 = N861 | pegMaxFiniteMagOut;
  assign N861 = N860 | pegMinNonzeroMagOut;
  assign N860 = N858 & N859;
  assign N858 = \genblk2.sRoundedExp [9] & N847;
  assign N859 = ~notNaN_isInfOut;
  assign out[60] = N863 | pegMaxFiniteMagOut;
  assign N863 = \genblk2.sRoundedExp [8] | pegMinNonzeroMagOut;
  assign out[59] = N864 | pegMaxFiniteMagOut;
  assign N864 = \genblk2.sRoundedExp [7] | pegMinNonzeroMagOut;
  assign out[58] = N865 | pegMaxFiniteMagOut;
  assign N865 = \genblk2.sRoundedExp [6] | pegMinNonzeroMagOut;
  assign out[57] = N866 | pegMaxFiniteMagOut;
  assign N866 = \genblk2.sRoundedExp [5] & N849;
  assign out[56] = N867 | pegMaxFiniteMagOut;
  assign N867 = \genblk2.sRoundedExp [4] & N849;
  assign out[55] = N868 | pegMaxFiniteMagOut;
  assign N868 = \genblk2.sRoundedExp [3] | pegMinNonzeroMagOut;
  assign out[54] = N869 | pegMaxFiniteMagOut;
  assign N869 = \genblk2.sRoundedExp [2] | pegMinNonzeroMagOut;
  assign out[53] = N870 | pegMaxFiniteMagOut;
  assign N870 = \genblk2.sRoundedExp [1] | pegMinNonzeroMagOut;
  assign out[52] = N871 | pegMaxFiniteMagOut;
  assign N871 = \genblk2.sRoundedExp [0] & N849;
  assign N357 = N840 & N872;
  assign N872 = ~common_totalUnderflow;
  assign N358 = ~N357;
  assign N360 = N873 & N872;
  assign N873 = N837 & N840;
  assign N361 = ~N360;
  assign out[51] = N874 | pegMaxFiniteMagOut;
  assign N874 = isNaNOut | N359;
  assign out[50] = N412 | pegMaxFiniteMagOut;
  assign out[49] = N411 | pegMaxFiniteMagOut;
  assign out[48] = N410 | pegMaxFiniteMagOut;
  assign out[47] = N409 | pegMaxFiniteMagOut;
  assign out[46] = N408 | pegMaxFiniteMagOut;
  assign out[45] = N407 | pegMaxFiniteMagOut;
  assign out[44] = N406 | pegMaxFiniteMagOut;
  assign out[43] = N405 | pegMaxFiniteMagOut;
  assign out[42] = N404 | pegMaxFiniteMagOut;
  assign out[41] = N403 | pegMaxFiniteMagOut;
  assign out[40] = N402 | pegMaxFiniteMagOut;
  assign out[39] = N401 | pegMaxFiniteMagOut;
  assign out[38] = N400 | pegMaxFiniteMagOut;
  assign out[37] = N399 | pegMaxFiniteMagOut;
  assign out[36] = N398 | pegMaxFiniteMagOut;
  assign out[35] = N397 | pegMaxFiniteMagOut;
  assign out[34] = N396 | pegMaxFiniteMagOut;
  assign out[33] = N395 | pegMaxFiniteMagOut;
  assign out[32] = N394 | pegMaxFiniteMagOut;
  assign out[31] = N393 | pegMaxFiniteMagOut;
  assign out[30] = N392 | pegMaxFiniteMagOut;
  assign out[29] = N391 | pegMaxFiniteMagOut;
  assign out[28] = N390 | pegMaxFiniteMagOut;
  assign out[27] = N389 | pegMaxFiniteMagOut;
  assign out[26] = N388 | pegMaxFiniteMagOut;
  assign out[25] = N387 | pegMaxFiniteMagOut;
  assign out[24] = N386 | pegMaxFiniteMagOut;
  assign out[23] = N385 | pegMaxFiniteMagOut;
  assign out[22] = N384 | pegMaxFiniteMagOut;
  assign out[21] = N383 | pegMaxFiniteMagOut;
  assign out[20] = N382 | pegMaxFiniteMagOut;
  assign out[19] = N381 | pegMaxFiniteMagOut;
  assign out[18] = N380 | pegMaxFiniteMagOut;
  assign out[17] = N379 | pegMaxFiniteMagOut;
  assign out[16] = N378 | pegMaxFiniteMagOut;
  assign out[15] = N377 | pegMaxFiniteMagOut;
  assign out[14] = N376 | pegMaxFiniteMagOut;
  assign out[13] = N375 | pegMaxFiniteMagOut;
  assign out[12] = N374 | pegMaxFiniteMagOut;
  assign out[11] = N373 | pegMaxFiniteMagOut;
  assign out[10] = N372 | pegMaxFiniteMagOut;
  assign out[9] = N371 | pegMaxFiniteMagOut;
  assign out[8] = N370 | pegMaxFiniteMagOut;
  assign out[7] = N369 | pegMaxFiniteMagOut;
  assign out[6] = N368 | pegMaxFiniteMagOut;
  assign out[5] = N367 | pegMaxFiniteMagOut;
  assign out[4] = N366 | pegMaxFiniteMagOut;
  assign out[3] = N365 | pegMaxFiniteMagOut;
  assign out[2] = N364 | pegMaxFiniteMagOut;
  assign out[1] = N363 | pegMaxFiniteMagOut;
  assign out[0] = N362 | pegMaxFiniteMagOut;

endmodule



module reverse_width25
(
  in,
  out
);

  input [24:0] in;
  output [24:0] out;
  wire [24:0] out;
  assign out[24] = in[0];
  assign out[23] = in[1];
  assign out[22] = in[2];
  assign out[21] = in[3];
  assign out[20] = in[4];
  assign out[19] = in[5];
  assign out[18] = in[6];
  assign out[17] = in[7];
  assign out[16] = in[8];
  assign out[15] = in[9];
  assign out[14] = in[10];
  assign out[13] = in[11];
  assign out[12] = in[12];
  assign out[11] = in[13];
  assign out[10] = in[14];
  assign out[9] = in[15];
  assign out[8] = in[16];
  assign out[7] = in[17];
  assign out[6] = in[18];
  assign out[5] = in[19];
  assign out[4] = in[20];
  assign out[3] = in[21];
  assign out[2] = in[22];
  assign out[1] = in[23];
  assign out[0] = in[24];

endmodule



module lowMaskLoHi_inWidth9_topBound105_bottomBound130
(
  in,
  out
);

  input [8:0] in;
  output [24:0] out;
  wire [24:0] out,reverseOut;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,
  sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,
  sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,
  sv2v_dc_21,sv2v_dc_22,sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,sv2v_dc_27,
  sv2v_dc_28,sv2v_dc_29,sv2v_dc_30,sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,sv2v_dc_34,
  sv2v_dc_35,sv2v_dc_36,sv2v_dc_37,sv2v_dc_38,sv2v_dc_39,sv2v_dc_40,sv2v_dc_41,sv2v_dc_42,
  sv2v_dc_43,sv2v_dc_44,sv2v_dc_45,sv2v_dc_46,sv2v_dc_47,sv2v_dc_48,sv2v_dc_49,
  sv2v_dc_50,sv2v_dc_51,sv2v_dc_52,sv2v_dc_53,sv2v_dc_54,sv2v_dc_55,sv2v_dc_56,
  sv2v_dc_57,sv2v_dc_58,sv2v_dc_59,sv2v_dc_60,sv2v_dc_61,sv2v_dc_62,sv2v_dc_63,
  sv2v_dc_64,sv2v_dc_65,sv2v_dc_66,sv2v_dc_67,sv2v_dc_68,sv2v_dc_69,sv2v_dc_70,sv2v_dc_71,
  sv2v_dc_72,sv2v_dc_73,sv2v_dc_74,sv2v_dc_75,sv2v_dc_76,sv2v_dc_77,sv2v_dc_78,
  sv2v_dc_79,sv2v_dc_80,sv2v_dc_81,sv2v_dc_82,sv2v_dc_83,sv2v_dc_84,sv2v_dc_85,
  sv2v_dc_86,sv2v_dc_87,sv2v_dc_88,sv2v_dc_89,sv2v_dc_90,sv2v_dc_91,sv2v_dc_92,
  sv2v_dc_93,sv2v_dc_94,sv2v_dc_95,sv2v_dc_96,sv2v_dc_97,sv2v_dc_98,sv2v_dc_99,sv2v_dc_100,
  sv2v_dc_101,sv2v_dc_102,sv2v_dc_103,sv2v_dc_104,sv2v_dc_105,sv2v_dc_106,
  sv2v_dc_107,sv2v_dc_108,sv2v_dc_109,sv2v_dc_110,sv2v_dc_111,sv2v_dc_112,sv2v_dc_113,
  sv2v_dc_114,sv2v_dc_115,sv2v_dc_116,sv2v_dc_117,sv2v_dc_118,sv2v_dc_119,sv2v_dc_120,
  sv2v_dc_121,sv2v_dc_122,sv2v_dc_123,sv2v_dc_124,sv2v_dc_125,sv2v_dc_126,
  sv2v_dc_127,sv2v_dc_128,sv2v_dc_129,sv2v_dc_130,sv2v_dc_131,sv2v_dc_132,sv2v_dc_133,
  sv2v_dc_134,sv2v_dc_135,sv2v_dc_136,sv2v_dc_137,sv2v_dc_138,sv2v_dc_139,sv2v_dc_140,
  sv2v_dc_141,sv2v_dc_142,sv2v_dc_143,sv2v_dc_144,sv2v_dc_145,sv2v_dc_146,
  sv2v_dc_147,sv2v_dc_148,sv2v_dc_149,sv2v_dc_150,sv2v_dc_151,sv2v_dc_152,sv2v_dc_153,
  sv2v_dc_154,sv2v_dc_155,sv2v_dc_156,sv2v_dc_157,sv2v_dc_158,sv2v_dc_159,sv2v_dc_160,
  sv2v_dc_161,sv2v_dc_162,sv2v_dc_163,sv2v_dc_164,sv2v_dc_165,sv2v_dc_166,
  sv2v_dc_167,sv2v_dc_168,sv2v_dc_169,sv2v_dc_170,sv2v_dc_171,sv2v_dc_172,sv2v_dc_173,
  sv2v_dc_174,sv2v_dc_175,sv2v_dc_176,sv2v_dc_177,sv2v_dc_178,sv2v_dc_179,sv2v_dc_180,
  sv2v_dc_181,sv2v_dc_182,sv2v_dc_183,sv2v_dc_184,sv2v_dc_185,sv2v_dc_186,
  sv2v_dc_187,sv2v_dc_188,sv2v_dc_189,sv2v_dc_190,sv2v_dc_191,sv2v_dc_192,sv2v_dc_193,
  sv2v_dc_194,sv2v_dc_195,sv2v_dc_196,sv2v_dc_197,sv2v_dc_198,sv2v_dc_199,sv2v_dc_200,
  sv2v_dc_201,sv2v_dc_202,sv2v_dc_203,sv2v_dc_204,sv2v_dc_205,sv2v_dc_206,
  sv2v_dc_207,sv2v_dc_208,sv2v_dc_209,sv2v_dc_210,sv2v_dc_211,sv2v_dc_212,sv2v_dc_213,
  sv2v_dc_214,sv2v_dc_215,sv2v_dc_216,sv2v_dc_217,sv2v_dc_218,sv2v_dc_219,sv2v_dc_220,
  sv2v_dc_221,sv2v_dc_222,sv2v_dc_223,sv2v_dc_224,sv2v_dc_225,sv2v_dc_226,
  sv2v_dc_227,sv2v_dc_228,sv2v_dc_229,sv2v_dc_230,sv2v_dc_231,sv2v_dc_232,sv2v_dc_233,
  sv2v_dc_234,sv2v_dc_235,sv2v_dc_236,sv2v_dc_237,sv2v_dc_238,sv2v_dc_239,sv2v_dc_240,
  sv2v_dc_241,sv2v_dc_242,sv2v_dc_243,sv2v_dc_244,sv2v_dc_245,sv2v_dc_246,
  sv2v_dc_247,sv2v_dc_248,sv2v_dc_249,sv2v_dc_250,sv2v_dc_251,sv2v_dc_252,sv2v_dc_253,
  sv2v_dc_254,sv2v_dc_255,sv2v_dc_256,sv2v_dc_257,sv2v_dc_258,sv2v_dc_259,sv2v_dc_260,
  sv2v_dc_261,sv2v_dc_262,sv2v_dc_263,sv2v_dc_264,sv2v_dc_265,sv2v_dc_266,
  sv2v_dc_267,sv2v_dc_268,sv2v_dc_269,sv2v_dc_270,sv2v_dc_271,sv2v_dc_272,sv2v_dc_273,
  sv2v_dc_274,sv2v_dc_275,sv2v_dc_276,sv2v_dc_277,sv2v_dc_278,sv2v_dc_279,sv2v_dc_280,
  sv2v_dc_281,sv2v_dc_282,sv2v_dc_283,sv2v_dc_284,sv2v_dc_285,sv2v_dc_286,
  sv2v_dc_287,sv2v_dc_288,sv2v_dc_289,sv2v_dc_290,sv2v_dc_291,sv2v_dc_292,sv2v_dc_293,
  sv2v_dc_294,sv2v_dc_295,sv2v_dc_296,sv2v_dc_297,sv2v_dc_298,sv2v_dc_299,sv2v_dc_300,
  sv2v_dc_301,sv2v_dc_302,sv2v_dc_303,sv2v_dc_304,sv2v_dc_305,sv2v_dc_306,
  sv2v_dc_307,sv2v_dc_308,sv2v_dc_309,sv2v_dc_310,sv2v_dc_311,sv2v_dc_312,sv2v_dc_313,
  sv2v_dc_314,sv2v_dc_315,sv2v_dc_316,sv2v_dc_317,sv2v_dc_318,sv2v_dc_319,sv2v_dc_320,
  sv2v_dc_321,sv2v_dc_322,sv2v_dc_323,sv2v_dc_324,sv2v_dc_325,sv2v_dc_326,
  sv2v_dc_327,sv2v_dc_328,sv2v_dc_329,sv2v_dc_330,sv2v_dc_331,sv2v_dc_332,sv2v_dc_333,
  sv2v_dc_334,sv2v_dc_335,sv2v_dc_336,sv2v_dc_337,sv2v_dc_338,sv2v_dc_339,sv2v_dc_340,
  sv2v_dc_341,sv2v_dc_342,sv2v_dc_343,sv2v_dc_344,sv2v_dc_345,sv2v_dc_346,
  sv2v_dc_347,sv2v_dc_348,sv2v_dc_349,sv2v_dc_350,sv2v_dc_351,sv2v_dc_352,sv2v_dc_353,
  sv2v_dc_354,sv2v_dc_355,sv2v_dc_356,sv2v_dc_357,sv2v_dc_358,sv2v_dc_359,sv2v_dc_360,
  sv2v_dc_361,sv2v_dc_362,sv2v_dc_363,sv2v_dc_364,sv2v_dc_365,sv2v_dc_366,
  sv2v_dc_367,sv2v_dc_368,sv2v_dc_369,sv2v_dc_370,sv2v_dc_371,sv2v_dc_372,sv2v_dc_373,
  sv2v_dc_374,sv2v_dc_375,sv2v_dc_376,sv2v_dc_377,sv2v_dc_378,sv2v_dc_379,sv2v_dc_380,
  sv2v_dc_381,sv2v_dc_382;

  reverse_width25
  reverse
  (
    .in(reverseOut),
    .out(out)
  );

  assign { sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36, sv2v_dc_37, sv2v_dc_38, sv2v_dc_39, sv2v_dc_40, sv2v_dc_41, sv2v_dc_42, sv2v_dc_43, sv2v_dc_44, sv2v_dc_45, sv2v_dc_46, sv2v_dc_47, sv2v_dc_48, sv2v_dc_49, sv2v_dc_50, sv2v_dc_51, sv2v_dc_52, sv2v_dc_53, sv2v_dc_54, sv2v_dc_55, sv2v_dc_56, sv2v_dc_57, sv2v_dc_58, sv2v_dc_59, sv2v_dc_60, sv2v_dc_61, sv2v_dc_62, sv2v_dc_63, sv2v_dc_64, sv2v_dc_65, sv2v_dc_66, sv2v_dc_67, sv2v_dc_68, sv2v_dc_69, sv2v_dc_70, sv2v_dc_71, sv2v_dc_72, sv2v_dc_73, sv2v_dc_74, sv2v_dc_75, sv2v_dc_76, sv2v_dc_77, sv2v_dc_78, sv2v_dc_79, sv2v_dc_80, sv2v_dc_81, sv2v_dc_82, sv2v_dc_83, sv2v_dc_84, sv2v_dc_85, sv2v_dc_86, sv2v_dc_87, sv2v_dc_88, sv2v_dc_89, sv2v_dc_90, sv2v_dc_91, sv2v_dc_92, sv2v_dc_93, sv2v_dc_94, sv2v_dc_95, sv2v_dc_96, sv2v_dc_97, sv2v_dc_98, sv2v_dc_99, sv2v_dc_100, sv2v_dc_101, sv2v_dc_102, sv2v_dc_103, sv2v_dc_104, sv2v_dc_105, sv2v_dc_106, sv2v_dc_107, sv2v_dc_108, sv2v_dc_109, sv2v_dc_110, sv2v_dc_111, sv2v_dc_112, sv2v_dc_113, sv2v_dc_114, sv2v_dc_115, sv2v_dc_116, sv2v_dc_117, sv2v_dc_118, sv2v_dc_119, sv2v_dc_120, sv2v_dc_121, sv2v_dc_122, sv2v_dc_123, sv2v_dc_124, sv2v_dc_125, sv2v_dc_126, sv2v_dc_127, sv2v_dc_128, sv2v_dc_129, sv2v_dc_130, sv2v_dc_131, sv2v_dc_132, sv2v_dc_133, sv2v_dc_134, sv2v_dc_135, sv2v_dc_136, sv2v_dc_137, sv2v_dc_138, sv2v_dc_139, sv2v_dc_140, sv2v_dc_141, sv2v_dc_142, sv2v_dc_143, sv2v_dc_144, sv2v_dc_145, sv2v_dc_146, sv2v_dc_147, sv2v_dc_148, sv2v_dc_149, sv2v_dc_150, sv2v_dc_151, sv2v_dc_152, sv2v_dc_153, sv2v_dc_154, sv2v_dc_155, sv2v_dc_156, sv2v_dc_157, sv2v_dc_158, sv2v_dc_159, sv2v_dc_160, sv2v_dc_161, sv2v_dc_162, sv2v_dc_163, sv2v_dc_164, sv2v_dc_165, sv2v_dc_166, sv2v_dc_167, sv2v_dc_168, sv2v_dc_169, sv2v_dc_170, sv2v_dc_171, sv2v_dc_172, sv2v_dc_173, sv2v_dc_174, sv2v_dc_175, sv2v_dc_176, sv2v_dc_177, sv2v_dc_178, sv2v_dc_179, sv2v_dc_180, sv2v_dc_181, sv2v_dc_182, sv2v_dc_183, sv2v_dc_184, sv2v_dc_185, sv2v_dc_186, sv2v_dc_187, sv2v_dc_188, sv2v_dc_189, sv2v_dc_190, sv2v_dc_191, sv2v_dc_192, sv2v_dc_193, sv2v_dc_194, sv2v_dc_195, sv2v_dc_196, sv2v_dc_197, sv2v_dc_198, sv2v_dc_199, sv2v_dc_200, sv2v_dc_201, sv2v_dc_202, sv2v_dc_203, sv2v_dc_204, sv2v_dc_205, sv2v_dc_206, sv2v_dc_207, sv2v_dc_208, sv2v_dc_209, sv2v_dc_210, sv2v_dc_211, sv2v_dc_212, sv2v_dc_213, sv2v_dc_214, sv2v_dc_215, sv2v_dc_216, sv2v_dc_217, sv2v_dc_218, sv2v_dc_219, sv2v_dc_220, sv2v_dc_221, sv2v_dc_222, sv2v_dc_223, sv2v_dc_224, sv2v_dc_225, sv2v_dc_226, sv2v_dc_227, sv2v_dc_228, sv2v_dc_229, sv2v_dc_230, sv2v_dc_231, sv2v_dc_232, sv2v_dc_233, sv2v_dc_234, sv2v_dc_235, sv2v_dc_236, sv2v_dc_237, sv2v_dc_238, sv2v_dc_239, sv2v_dc_240, sv2v_dc_241, sv2v_dc_242, sv2v_dc_243, sv2v_dc_244, sv2v_dc_245, sv2v_dc_246, sv2v_dc_247, sv2v_dc_248, sv2v_dc_249, sv2v_dc_250, sv2v_dc_251, sv2v_dc_252, sv2v_dc_253, sv2v_dc_254, sv2v_dc_255, sv2v_dc_256, sv2v_dc_257, sv2v_dc_258, sv2v_dc_259, sv2v_dc_260, sv2v_dc_261, sv2v_dc_262, sv2v_dc_263, sv2v_dc_264, sv2v_dc_265, sv2v_dc_266, sv2v_dc_267, sv2v_dc_268, sv2v_dc_269, sv2v_dc_270, sv2v_dc_271, sv2v_dc_272, sv2v_dc_273, sv2v_dc_274, sv2v_dc_275, sv2v_dc_276, sv2v_dc_277, sv2v_dc_278, sv2v_dc_279, sv2v_dc_280, sv2v_dc_281, sv2v_dc_282, sv2v_dc_283, sv2v_dc_284, sv2v_dc_285, sv2v_dc_286, sv2v_dc_287, sv2v_dc_288, sv2v_dc_289, sv2v_dc_290, sv2v_dc_291, sv2v_dc_292, sv2v_dc_293, sv2v_dc_294, sv2v_dc_295, sv2v_dc_296, sv2v_dc_297, sv2v_dc_298, sv2v_dc_299, sv2v_dc_300, sv2v_dc_301, sv2v_dc_302, sv2v_dc_303, sv2v_dc_304, sv2v_dc_305, sv2v_dc_306, sv2v_dc_307, sv2v_dc_308, sv2v_dc_309, sv2v_dc_310, sv2v_dc_311, sv2v_dc_312, sv2v_dc_313, sv2v_dc_314, sv2v_dc_315, sv2v_dc_316, sv2v_dc_317, sv2v_dc_318, sv2v_dc_319, sv2v_dc_320, sv2v_dc_321, sv2v_dc_322, sv2v_dc_323, sv2v_dc_324, sv2v_dc_325, sv2v_dc_326, sv2v_dc_327, sv2v_dc_328, sv2v_dc_329, sv2v_dc_330, sv2v_dc_331, sv2v_dc_332, sv2v_dc_333, sv2v_dc_334, sv2v_dc_335, sv2v_dc_336, sv2v_dc_337, sv2v_dc_338, sv2v_dc_339, sv2v_dc_340, sv2v_dc_341, sv2v_dc_342, sv2v_dc_343, sv2v_dc_344, sv2v_dc_345, sv2v_dc_346, sv2v_dc_347, sv2v_dc_348, sv2v_dc_349, sv2v_dc_350, sv2v_dc_351, sv2v_dc_352, sv2v_dc_353, sv2v_dc_354, sv2v_dc_355, sv2v_dc_356, sv2v_dc_357, sv2v_dc_358, sv2v_dc_359, sv2v_dc_360, sv2v_dc_361, sv2v_dc_362, sv2v_dc_363, sv2v_dc_364, sv2v_dc_365, sv2v_dc_366, sv2v_dc_367, sv2v_dc_368, sv2v_dc_369, sv2v_dc_370, sv2v_dc_371, sv2v_dc_372, sv2v_dc_373, sv2v_dc_374, sv2v_dc_375, sv2v_dc_376, sv2v_dc_377, sv2v_dc_378, sv2v_dc_379, sv2v_dc_380, sv2v_dc_381, sv2v_dc_382, reverseOut } = $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) >>> { N0, N1, N2, N3, N4, N5, N6, N7, N8 };
  assign N0 = ~in[8];
  assign N1 = ~in[7];
  assign N2 = ~in[6];
  assign N3 = ~in[5];
  assign N4 = ~in[4];
  assign N5 = ~in[3];
  assign N6 = ~in[2];
  assign N7 = ~in[1];
  assign N8 = ~in[0];

endmodule



module roundAnyRawFNToRecFN_inExpWidth11_inSigWidth55_outExpWidth8_outSigWidth24
(
  control,
  invalidExc,
  infiniteExc,
  in_isNaN,
  in_isInf,
  in_isZero,
  in_sign,
  in_sExp,
  in_sig,
  roundingMode,
  out,
  exceptionFlags
);

  input [0:0] control;
  input [12:0] in_sExp;
  input [55:0] in_sig;
  input [2:0] roundingMode;
  output [32:0] out;
  output [4:0] exceptionFlags;
  input invalidExc;
  input infiniteExc;
  input in_isNaN;
  input in_isInf;
  input in_isZero;
  input in_sign;
  wire [32:0] out;
  wire [4:0] exceptionFlags;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,exceptionFlags_4_,
  exceptionFlags_3_,roundMagUp,isNaNOut,_0_net__8_,\genblk2.roundPosBit ,\genblk2.anyRoundExtra ,
  \genblk2.anyRound ,\genblk2.roundIncr ,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,
  N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,
  N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,
  N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,
  N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,
  N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,
  N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,
  N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,
  N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,
  N167,N168,N169,N170,N171,N172,common_overflow,common_totalUnderflow,
  \genblk2.unboundedRange_roundPosBit ,\genblk2.unboundedRange_anyRound ,
  \genblk2.unboundedRange_roundIncr ,\genblk2.roundCarry ,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  common_underflow,common_inexact,notNaN_isSpecialInfOut,commonCase,
  overflow_roundMagUp,pegMinNonzeroMagOut,pegMaxFiniteMagOut,notNaN_isInfOut,N182,N183,N184,N185,
  N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,
  N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,
  N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,
  N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,
  N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,
  N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,
  N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,
  N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,
  N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,
  N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,
  N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,
  N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,
  N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,
  N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,
  N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,
  N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,
  N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,
  N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,
  N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,
  N490,N491,N492,N493;
  wire [13:0] sAdjustedExp;
  wire [0:0] adjustedSig;
  wire [24:0] \genblk2.genblk1.roundMask_main ;
  wire [2:2] \genblk2.roundMask ;
  wire [26:0] \genblk2.roundPosMask ;
  wire [25:0] \genblk2.roundedSig ;
  wire [14:0] \genblk2.sRoundedExp ;
  wire [22:0] common_fractOut;
  assign exceptionFlags_4_ = invalidExc;
  assign exceptionFlags[4] = exceptionFlags_4_;
  assign exceptionFlags_3_ = infiniteExc;
  assign exceptionFlags[3] = exceptionFlags_3_;

  lowMaskLoHi_inWidth9_topBound105_bottomBound130
  \genblk2.genblk1.lowMask_roundMask 
  (
    .in({ _0_net__8_, sAdjustedExp[7:0] }),
    .out(\genblk2.genblk1.roundMask_main )
  );

  assign common_overflow = $signed(\genblk2.sRoundedExp [14:7]) >= $signed({ 1'b0, 1'b1, 1'b1 });
  assign common_totalUnderflow = $signed(\genblk2.sRoundedExp ) < $signed({ 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1 });
  assign N174 = $signed(sAdjustedExp[13:8]) <= $signed(1'b0);
  assign N210 = ~roundingMode[2];
  assign N211 = ~roundingMode[1];
  assign N212 = N211 | N210;
  assign N213 = roundingMode[0] | N212;
  assign N214 = ~N213;
  assign N215 = roundingMode[1] | N210;
  assign N216 = roundingMode[0] | N215;
  assign N217 = ~N216;
  assign N218 = roundingMode[1] | roundingMode[2];
  assign N219 = roundingMode[0] | N218;
  assign N220 = ~N219;
  assign N221 = N211 | roundingMode[2];
  assign N222 = roundingMode[0] | N221;
  assign N223 = ~N222;
  assign N224 = ~roundingMode[0];
  assign N225 = N224 | N221;
  assign N226 = ~N225;
  assign sAdjustedExp = $signed(in_sExp) + $signed({ 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 });
  assign { N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67 } = { N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66 } + 1'b1;
  assign \genblk2.sRoundedExp  = { sAdjustedExp[13:13], sAdjustedExp } + \genblk2.roundedSig [25:24];
  assign { N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17 } = (N0)? { \genblk2.genblk1.roundMask_main [24:1], \genblk2.roundMask [2:2] } : 
                                                                                                                                           (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N15;
  assign { N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121 } = (N1)? \genblk2.roundPosMask [26:1] : 
                                                                                                                                                                          (N120)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = N119;
  assign \genblk2.roundedSig  = (N2)? { N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118 } : 
                                (N3)? { N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171 } : 1'b0;
  assign N2 = \genblk2.roundIncr ;
  assign N3 = N14;
  assign common_fractOut = (N4)? \genblk2.roundedSig [23:1] : 
                           (N5)? \genblk2.roundedSig [22:0] : 1'b0;
  assign N4 = in_sig[55];
  assign N5 = N172;
  assign \genblk2.unboundedRange_roundPosBit  = (N4)? in_sig[31] : 
                                                (N5)? in_sig[30] : 1'b0;
  assign \genblk2.roundCarry  = (N4)? \genblk2.roundedSig [25] : 
                                (N5)? \genblk2.roundedSig [24] : 1'b0;
  assign N173 = (N4)? \genblk2.genblk1.roundMask_main [1] : 
                (N5)? \genblk2.roundMask [2] : 1'b0;
  assign N177 = (N6)? N173 : 
                (N7)? 1'b0 : 1'b0;
  assign N6 = N175;
  assign N7 = N176;
  assign N178 = (N4)? \genblk2.genblk1.roundMask_main [2] : 
                (N5)? \genblk2.genblk1.roundMask_main [1] : 1'b0;
  assign N181 = (N8)? N180 : 
                (N9)? 1'b0 : 1'b0;
  assign N8 = control[0];
  assign N9 = N179;
  assign out[32] = (N10)? 1'b0 : 
                   (N11)? in_sign : 1'b0;
  assign N10 = isNaNOut;
  assign N11 = N459;
  assign N185 = (N12)? common_fractOut[22] : 
                (N184)? 1'b0 : 1'b0;
  assign N12 = N183;
  assign { N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188 } = (N13)? common_fractOut[21:0] : 
                                                                                                                                                  (N187)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = N186;
  assign roundMagUp = N227 | N229;
  assign N227 = N223 & in_sign;
  assign N229 = N226 & N228;
  assign N228 = ~in_sign;
  assign isNaNOut = exceptionFlags_4_ | N231;
  assign N231 = N230 & in_isNaN;
  assign N230 = ~exceptionFlags_3_;
  assign adjustedSig[0] = N259 | in_sig[0];
  assign N259 = N258 | in_sig[1];
  assign N258 = N257 | in_sig[2];
  assign N257 = N256 | in_sig[3];
  assign N256 = N255 | in_sig[4];
  assign N255 = N254 | in_sig[5];
  assign N254 = N253 | in_sig[6];
  assign N253 = N252 | in_sig[7];
  assign N252 = N251 | in_sig[8];
  assign N251 = N250 | in_sig[9];
  assign N250 = N249 | in_sig[10];
  assign N249 = N248 | in_sig[11];
  assign N248 = N247 | in_sig[12];
  assign N247 = N246 | in_sig[13];
  assign N246 = N245 | in_sig[14];
  assign N245 = N244 | in_sig[15];
  assign N244 = N243 | in_sig[16];
  assign N243 = N242 | in_sig[17];
  assign N242 = N241 | in_sig[18];
  assign N241 = N240 | in_sig[19];
  assign N240 = N239 | in_sig[20];
  assign N239 = N238 | in_sig[21];
  assign N238 = N237 | in_sig[22];
  assign N237 = N236 | in_sig[23];
  assign N236 = N235 | in_sig[24];
  assign N235 = N234 | in_sig[25];
  assign N234 = N233 | in_sig[26];
  assign N233 = N232 | in_sig[27];
  assign N232 = in_sig[29] | in_sig[28];
  assign _0_net__8_ = sAdjustedExp[8] | 1'b0;
  assign \genblk2.roundMask [2] = \genblk2.genblk1.roundMask_main [0] | in_sig[55];
  assign \genblk2.roundPosMask [26] = N260 & \genblk2.genblk1.roundMask_main [24];
  assign N260 = ~1'b0;
  assign \genblk2.roundPosMask [25] = N261 & \genblk2.genblk1.roundMask_main [23];
  assign N261 = ~\genblk2.genblk1.roundMask_main [24];
  assign \genblk2.roundPosMask [24] = N262 & \genblk2.genblk1.roundMask_main [22];
  assign N262 = ~\genblk2.genblk1.roundMask_main [23];
  assign \genblk2.roundPosMask [23] = N263 & \genblk2.genblk1.roundMask_main [21];
  assign N263 = ~\genblk2.genblk1.roundMask_main [22];
  assign \genblk2.roundPosMask [22] = N264 & \genblk2.genblk1.roundMask_main [20];
  assign N264 = ~\genblk2.genblk1.roundMask_main [21];
  assign \genblk2.roundPosMask [21] = N265 & \genblk2.genblk1.roundMask_main [19];
  assign N265 = ~\genblk2.genblk1.roundMask_main [20];
  assign \genblk2.roundPosMask [20] = N266 & \genblk2.genblk1.roundMask_main [18];
  assign N266 = ~\genblk2.genblk1.roundMask_main [19];
  assign \genblk2.roundPosMask [19] = N267 & \genblk2.genblk1.roundMask_main [17];
  assign N267 = ~\genblk2.genblk1.roundMask_main [18];
  assign \genblk2.roundPosMask [18] = N268 & \genblk2.genblk1.roundMask_main [16];
  assign N268 = ~\genblk2.genblk1.roundMask_main [17];
  assign \genblk2.roundPosMask [17] = N269 & \genblk2.genblk1.roundMask_main [15];
  assign N269 = ~\genblk2.genblk1.roundMask_main [16];
  assign \genblk2.roundPosMask [16] = N270 & \genblk2.genblk1.roundMask_main [14];
  assign N270 = ~\genblk2.genblk1.roundMask_main [15];
  assign \genblk2.roundPosMask [15] = N271 & \genblk2.genblk1.roundMask_main [13];
  assign N271 = ~\genblk2.genblk1.roundMask_main [14];
  assign \genblk2.roundPosMask [14] = N272 & \genblk2.genblk1.roundMask_main [12];
  assign N272 = ~\genblk2.genblk1.roundMask_main [13];
  assign \genblk2.roundPosMask [13] = N273 & \genblk2.genblk1.roundMask_main [11];
  assign N273 = ~\genblk2.genblk1.roundMask_main [12];
  assign \genblk2.roundPosMask [12] = N274 & \genblk2.genblk1.roundMask_main [10];
  assign N274 = ~\genblk2.genblk1.roundMask_main [11];
  assign \genblk2.roundPosMask [11] = N275 & \genblk2.genblk1.roundMask_main [9];
  assign N275 = ~\genblk2.genblk1.roundMask_main [10];
  assign \genblk2.roundPosMask [10] = N276 & \genblk2.genblk1.roundMask_main [8];
  assign N276 = ~\genblk2.genblk1.roundMask_main [9];
  assign \genblk2.roundPosMask [9] = N277 & \genblk2.genblk1.roundMask_main [7];
  assign N277 = ~\genblk2.genblk1.roundMask_main [8];
  assign \genblk2.roundPosMask [8] = N278 & \genblk2.genblk1.roundMask_main [6];
  assign N278 = ~\genblk2.genblk1.roundMask_main [7];
  assign \genblk2.roundPosMask [7] = N279 & \genblk2.genblk1.roundMask_main [5];
  assign N279 = ~\genblk2.genblk1.roundMask_main [6];
  assign \genblk2.roundPosMask [6] = N280 & \genblk2.genblk1.roundMask_main [4];
  assign N280 = ~\genblk2.genblk1.roundMask_main [5];
  assign \genblk2.roundPosMask [5] = N281 & \genblk2.genblk1.roundMask_main [3];
  assign N281 = ~\genblk2.genblk1.roundMask_main [4];
  assign \genblk2.roundPosMask [4] = N282 & \genblk2.genblk1.roundMask_main [2];
  assign N282 = ~\genblk2.genblk1.roundMask_main [3];
  assign \genblk2.roundPosMask [3] = N283 & \genblk2.genblk1.roundMask_main [1];
  assign N283 = ~\genblk2.genblk1.roundMask_main [2];
  assign \genblk2.roundPosMask [2] = N284 & \genblk2.roundMask [2];
  assign N284 = ~\genblk2.genblk1.roundMask_main [1];
  assign \genblk2.roundPosMask [1] = N285 & 1'b1;
  assign N285 = ~\genblk2.roundMask [2];
  assign \genblk2.roundPosMask [0] = N286 & 1'b1;
  assign N286 = ~1'b1;
  assign \genblk2.roundPosBit  = N333 | N339;
  assign N333 = N331 | N332;
  assign N331 = N329 | N330;
  assign N329 = N327 | N328;
  assign N327 = N325 | N326;
  assign N325 = N323 | N324;
  assign N323 = N321 | N322;
  assign N321 = N319 | N320;
  assign N319 = N317 | N318;
  assign N317 = N315 | N316;
  assign N315 = N313 | N314;
  assign N313 = N311 | N312;
  assign N311 = N309 | N310;
  assign N309 = N307 | N308;
  assign N307 = N305 | N306;
  assign N305 = N303 | N304;
  assign N303 = N301 | N302;
  assign N301 = N299 | N300;
  assign N299 = N297 | N298;
  assign N297 = N295 | N296;
  assign N295 = N293 | N294;
  assign N293 = N291 | N292;
  assign N291 = N289 | N290;
  assign N289 = N287 | N288;
  assign N287 = in_sig[55] & \genblk2.roundPosMask [26];
  assign N288 = in_sig[54] & \genblk2.roundPosMask [25];
  assign N290 = in_sig[53] & \genblk2.roundPosMask [24];
  assign N292 = in_sig[52] & \genblk2.roundPosMask [23];
  assign N294 = in_sig[51] & \genblk2.roundPosMask [22];
  assign N296 = in_sig[50] & \genblk2.roundPosMask [21];
  assign N298 = in_sig[49] & \genblk2.roundPosMask [20];
  assign N300 = in_sig[48] & \genblk2.roundPosMask [19];
  assign N302 = in_sig[47] & \genblk2.roundPosMask [18];
  assign N304 = in_sig[46] & \genblk2.roundPosMask [17];
  assign N306 = in_sig[45] & \genblk2.roundPosMask [16];
  assign N308 = in_sig[44] & \genblk2.roundPosMask [15];
  assign N310 = in_sig[43] & \genblk2.roundPosMask [14];
  assign N312 = in_sig[42] & \genblk2.roundPosMask [13];
  assign N314 = in_sig[41] & \genblk2.roundPosMask [12];
  assign N316 = in_sig[40] & \genblk2.roundPosMask [11];
  assign N318 = in_sig[39] & \genblk2.roundPosMask [10];
  assign N320 = in_sig[38] & \genblk2.roundPosMask [9];
  assign N322 = in_sig[37] & \genblk2.roundPosMask [8];
  assign N324 = in_sig[36] & \genblk2.roundPosMask [7];
  assign N326 = in_sig[35] & \genblk2.roundPosMask [6];
  assign N328 = in_sig[34] & \genblk2.roundPosMask [5];
  assign N330 = in_sig[33] & \genblk2.roundPosMask [4];
  assign N332 = in_sig[32] & \genblk2.roundPosMask [3];
  assign N339 = N338 & N260;
  assign N338 = N336 | N337;
  assign N336 = N334 | N335;
  assign N334 = in_sig[31] & \genblk2.roundPosMask [2];
  assign N335 = in_sig[30] & \genblk2.roundPosMask [1];
  assign N337 = adjustedSig[0] & \genblk2.roundPosMask [0];
  assign \genblk2.anyRoundExtra  = N386 | N392;
  assign N386 = N384 | N385;
  assign N384 = N382 | N383;
  assign N382 = N380 | N381;
  assign N380 = N378 | N379;
  assign N378 = N376 | N377;
  assign N376 = N374 | N375;
  assign N374 = N372 | N373;
  assign N372 = N370 | N371;
  assign N370 = N368 | N369;
  assign N368 = N366 | N367;
  assign N366 = N364 | N365;
  assign N364 = N362 | N363;
  assign N362 = N360 | N361;
  assign N360 = N358 | N359;
  assign N358 = N356 | N357;
  assign N356 = N354 | N355;
  assign N354 = N352 | N353;
  assign N352 = N350 | N351;
  assign N350 = N348 | N349;
  assign N348 = N346 | N347;
  assign N346 = N344 | N345;
  assign N344 = N342 | N343;
  assign N342 = N340 | N341;
  assign N340 = in_sig[55] & 1'b0;
  assign N341 = in_sig[54] & \genblk2.genblk1.roundMask_main [24];
  assign N343 = in_sig[53] & \genblk2.genblk1.roundMask_main [23];
  assign N345 = in_sig[52] & \genblk2.genblk1.roundMask_main [22];
  assign N347 = in_sig[51] & \genblk2.genblk1.roundMask_main [21];
  assign N349 = in_sig[50] & \genblk2.genblk1.roundMask_main [20];
  assign N351 = in_sig[49] & \genblk2.genblk1.roundMask_main [19];
  assign N353 = in_sig[48] & \genblk2.genblk1.roundMask_main [18];
  assign N355 = in_sig[47] & \genblk2.genblk1.roundMask_main [17];
  assign N357 = in_sig[46] & \genblk2.genblk1.roundMask_main [16];
  assign N359 = in_sig[45] & \genblk2.genblk1.roundMask_main [15];
  assign N361 = in_sig[44] & \genblk2.genblk1.roundMask_main [14];
  assign N363 = in_sig[43] & \genblk2.genblk1.roundMask_main [13];
  assign N365 = in_sig[42] & \genblk2.genblk1.roundMask_main [12];
  assign N367 = in_sig[41] & \genblk2.genblk1.roundMask_main [11];
  assign N369 = in_sig[40] & \genblk2.genblk1.roundMask_main [10];
  assign N371 = in_sig[39] & \genblk2.genblk1.roundMask_main [9];
  assign N373 = in_sig[38] & \genblk2.genblk1.roundMask_main [8];
  assign N375 = in_sig[37] & \genblk2.genblk1.roundMask_main [7];
  assign N377 = in_sig[36] & \genblk2.genblk1.roundMask_main [6];
  assign N379 = in_sig[35] & \genblk2.genblk1.roundMask_main [5];
  assign N381 = in_sig[34] & \genblk2.genblk1.roundMask_main [4];
  assign N383 = in_sig[33] & \genblk2.genblk1.roundMask_main [3];
  assign N385 = in_sig[32] & \genblk2.genblk1.roundMask_main [2];
  assign N392 = N391 & N260;
  assign N391 = N389 | N390;
  assign N389 = N387 | N388;
  assign N387 = in_sig[31] & \genblk2.genblk1.roundMask_main [1];
  assign N388 = in_sig[30] & \genblk2.roundMask [2];
  assign N390 = adjustedSig[0] & 1'b1;
  assign \genblk2.anyRound  = \genblk2.roundPosBit  | \genblk2.anyRoundExtra ;
  assign \genblk2.roundIncr  = N394 | N395;
  assign N394 = N393 & \genblk2.roundPosBit ;
  assign N393 = N220 | N217;
  assign N395 = roundMagUp & \genblk2.anyRound ;
  assign N14 = ~\genblk2.roundIncr ;
  assign N15 = N396 & N397;
  assign N396 = N220 & \genblk2.roundPosBit ;
  assign N397 = ~\genblk2.anyRoundExtra ;
  assign N16 = ~N15;
  assign N42 = in_sig[55] | \genblk2.genblk1.roundMask_main [24];
  assign N43 = in_sig[54] | \genblk2.genblk1.roundMask_main [23];
  assign N44 = in_sig[53] | \genblk2.genblk1.roundMask_main [22];
  assign N45 = in_sig[52] | \genblk2.genblk1.roundMask_main [21];
  assign N46 = in_sig[51] | \genblk2.genblk1.roundMask_main [20];
  assign N47 = in_sig[50] | \genblk2.genblk1.roundMask_main [19];
  assign N48 = in_sig[49] | \genblk2.genblk1.roundMask_main [18];
  assign N49 = in_sig[48] | \genblk2.genblk1.roundMask_main [17];
  assign N50 = in_sig[47] | \genblk2.genblk1.roundMask_main [16];
  assign N51 = in_sig[46] | \genblk2.genblk1.roundMask_main [15];
  assign N52 = in_sig[45] | \genblk2.genblk1.roundMask_main [14];
  assign N53 = in_sig[44] | \genblk2.genblk1.roundMask_main [13];
  assign N54 = in_sig[43] | \genblk2.genblk1.roundMask_main [12];
  assign N55 = in_sig[42] | \genblk2.genblk1.roundMask_main [11];
  assign N56 = in_sig[41] | \genblk2.genblk1.roundMask_main [10];
  assign N57 = in_sig[40] | \genblk2.genblk1.roundMask_main [9];
  assign N58 = in_sig[39] | \genblk2.genblk1.roundMask_main [8];
  assign N59 = in_sig[38] | \genblk2.genblk1.roundMask_main [7];
  assign N60 = in_sig[37] | \genblk2.genblk1.roundMask_main [6];
  assign N61 = in_sig[36] | \genblk2.genblk1.roundMask_main [5];
  assign N62 = in_sig[35] | \genblk2.genblk1.roundMask_main [4];
  assign N63 = in_sig[34] | \genblk2.genblk1.roundMask_main [3];
  assign N64 = in_sig[33] | \genblk2.genblk1.roundMask_main [2];
  assign N65 = in_sig[32] | \genblk2.genblk1.roundMask_main [1];
  assign N66 = in_sig[31] | \genblk2.roundMask [2];
  assign N93 = N92 & N398;
  assign N398 = ~N41;
  assign N94 = N91 & N399;
  assign N399 = ~N40;
  assign N95 = N90 & N400;
  assign N400 = ~N39;
  assign N96 = N89 & N401;
  assign N401 = ~N38;
  assign N97 = N88 & N402;
  assign N402 = ~N37;
  assign N98 = N87 & N403;
  assign N403 = ~N36;
  assign N99 = N86 & N404;
  assign N404 = ~N35;
  assign N100 = N85 & N405;
  assign N405 = ~N34;
  assign N101 = N84 & N406;
  assign N406 = ~N33;
  assign N102 = N83 & N407;
  assign N407 = ~N32;
  assign N103 = N82 & N408;
  assign N408 = ~N31;
  assign N104 = N81 & N409;
  assign N409 = ~N30;
  assign N105 = N80 & N410;
  assign N410 = ~N29;
  assign N106 = N79 & N411;
  assign N411 = ~N28;
  assign N107 = N78 & N412;
  assign N412 = ~N27;
  assign N108 = N77 & N413;
  assign N413 = ~N26;
  assign N109 = N76 & N414;
  assign N414 = ~N25;
  assign N110 = N75 & N415;
  assign N415 = ~N24;
  assign N111 = N74 & N416;
  assign N416 = ~N23;
  assign N112 = N73 & N417;
  assign N417 = ~N22;
  assign N113 = N72 & N418;
  assign N418 = ~N21;
  assign N114 = N71 & N419;
  assign N419 = ~N20;
  assign N115 = N70 & N420;
  assign N420 = ~N19;
  assign N116 = N69 & N421;
  assign N421 = ~N18;
  assign N117 = N68 & N422;
  assign N422 = ~N17;
  assign N118 = N67 & N423;
  assign N423 = ~N15;
  assign N119 = N214 & \genblk2.anyRound ;
  assign N120 = ~N119;
  assign N147 = N424 | N145;
  assign N424 = in_sig[55] & N261;
  assign N148 = N425 | N144;
  assign N425 = in_sig[54] & N262;
  assign N149 = N426 | N143;
  assign N426 = in_sig[53] & N263;
  assign N150 = N427 | N142;
  assign N427 = in_sig[52] & N264;
  assign N151 = N428 | N141;
  assign N428 = in_sig[51] & N265;
  assign N152 = N429 | N140;
  assign N429 = in_sig[50] & N266;
  assign N153 = N430 | N139;
  assign N430 = in_sig[49] & N267;
  assign N154 = N431 | N138;
  assign N431 = in_sig[48] & N268;
  assign N155 = N432 | N137;
  assign N432 = in_sig[47] & N269;
  assign N156 = N433 | N136;
  assign N433 = in_sig[46] & N270;
  assign N157 = N434 | N135;
  assign N434 = in_sig[45] & N271;
  assign N158 = N435 | N134;
  assign N435 = in_sig[44] & N272;
  assign N159 = N436 | N133;
  assign N436 = in_sig[43] & N273;
  assign N160 = N437 | N132;
  assign N437 = in_sig[42] & N274;
  assign N161 = N438 | N131;
  assign N438 = in_sig[41] & N275;
  assign N162 = N439 | N130;
  assign N439 = in_sig[40] & N276;
  assign N163 = N440 | N129;
  assign N440 = in_sig[39] & N277;
  assign N164 = N441 | N128;
  assign N441 = in_sig[38] & N278;
  assign N165 = N442 | N127;
  assign N442 = in_sig[37] & N279;
  assign N166 = N443 | N126;
  assign N443 = in_sig[36] & N280;
  assign N167 = N444 | N125;
  assign N444 = in_sig[35] & N281;
  assign N168 = N445 | N124;
  assign N445 = in_sig[34] & N282;
  assign N169 = N446 | N123;
  assign N446 = in_sig[33] & N283;
  assign N170 = N447 | N122;
  assign N447 = in_sig[32] & N284;
  assign N171 = N448 | N121;
  assign N448 = in_sig[31] & N285;
  assign N172 = ~in_sig[55];
  assign \genblk2.unboundedRange_anyRound  = N449 | N450;
  assign N449 = in_sig[55] & in_sig[31];
  assign N450 = in_sig[30] | adjustedSig[0];
  assign \genblk2.unboundedRange_roundIncr  = N452 | N453;
  assign N452 = N451 & \genblk2.unboundedRange_roundPosBit ;
  assign N451 = N220 | N217;
  assign N453 = roundMagUp & \genblk2.unboundedRange_anyRound ;
  assign N175 = \genblk2.anyRound  & N174;
  assign N176 = ~N175;
  assign N179 = ~control[0];
  assign N180 = ~N178;
  assign common_underflow = common_totalUnderflow | N458;
  assign N458 = N177 & N457;
  assign N457 = ~N456;
  assign N456 = N455 & \genblk2.unboundedRange_roundIncr ;
  assign N455 = N454 & \genblk2.roundPosBit ;
  assign N454 = N181 & \genblk2.roundCarry ;
  assign common_inexact = common_totalUnderflow | \genblk2.anyRound ;
  assign notNaN_isSpecialInfOut = exceptionFlags_3_ | in_isInf;
  assign commonCase = N461 & N462;
  assign N461 = N459 & N460;
  assign N459 = ~isNaNOut;
  assign N460 = ~notNaN_isSpecialInfOut;
  assign N462 = ~in_isZero;
  assign exceptionFlags[2] = commonCase & common_overflow;
  assign exceptionFlags[1] = commonCase & common_underflow;
  assign exceptionFlags[0] = exceptionFlags[2] | N463;
  assign N463 = commonCase & common_inexact;
  assign overflow_roundMagUp = N464 | roundMagUp;
  assign N464 = N220 | N217;
  assign pegMinNonzeroMagOut = N465 & N466;
  assign N465 = commonCase & common_totalUnderflow;
  assign N466 = roundMagUp | N214;
  assign pegMaxFiniteMagOut = exceptionFlags[2] & N467;
  assign N467 = ~overflow_roundMagUp;
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | N468;
  assign N468 = exceptionFlags[2] & overflow_roundMagUp;
  assign N182 = in_isZero | common_totalUnderflow;
  assign out[31] = N474 | isNaNOut;
  assign N474 = N473 | notNaN_isInfOut;
  assign N473 = N472 | pegMaxFiniteMagOut;
  assign N472 = N470 & N471;
  assign N470 = \genblk2.sRoundedExp [8] & N469;
  assign N469 = ~N182;
  assign N471 = ~pegMinNonzeroMagOut;
  assign out[30] = N479 | isNaNOut;
  assign N479 = N478 | notNaN_isInfOut;
  assign N478 = N476 & N477;
  assign N476 = N475 & N471;
  assign N475 = \genblk2.sRoundedExp [7] & N469;
  assign N477 = ~pegMaxFiniteMagOut;
  assign out[29] = N484 | isNaNOut;
  assign N484 = N483 | pegMaxFiniteMagOut;
  assign N483 = N482 | pegMinNonzeroMagOut;
  assign N482 = N480 & N481;
  assign N480 = \genblk2.sRoundedExp [6] & N469;
  assign N481 = ~notNaN_isInfOut;
  assign out[28] = N485 | pegMaxFiniteMagOut;
  assign N485 = \genblk2.sRoundedExp [5] | pegMinNonzeroMagOut;
  assign out[27] = N486 | pegMaxFiniteMagOut;
  assign N486 = \genblk2.sRoundedExp [4] & N471;
  assign out[26] = N487 | pegMaxFiniteMagOut;
  assign N487 = \genblk2.sRoundedExp [3] | pegMinNonzeroMagOut;
  assign out[25] = N488 | pegMaxFiniteMagOut;
  assign N488 = \genblk2.sRoundedExp [2] & N471;
  assign out[24] = N489 | pegMaxFiniteMagOut;
  assign N489 = \genblk2.sRoundedExp [1] | pegMinNonzeroMagOut;
  assign out[23] = N490 | pegMaxFiniteMagOut;
  assign N490 = \genblk2.sRoundedExp [0] | pegMinNonzeroMagOut;
  assign N183 = N462 & N491;
  assign N491 = ~common_totalUnderflow;
  assign N184 = ~N183;
  assign N186 = N492 & N491;
  assign N492 = N459 & N462;
  assign N187 = ~N186;
  assign out[22] = N493 | pegMaxFiniteMagOut;
  assign N493 = isNaNOut | N185;
  assign out[21] = N209 | pegMaxFiniteMagOut;
  assign out[20] = N208 | pegMaxFiniteMagOut;
  assign out[19] = N207 | pegMaxFiniteMagOut;
  assign out[18] = N206 | pegMaxFiniteMagOut;
  assign out[17] = N205 | pegMaxFiniteMagOut;
  assign out[16] = N204 | pegMaxFiniteMagOut;
  assign out[15] = N203 | pegMaxFiniteMagOut;
  assign out[14] = N202 | pegMaxFiniteMagOut;
  assign out[13] = N201 | pegMaxFiniteMagOut;
  assign out[12] = N200 | pegMaxFiniteMagOut;
  assign out[11] = N199 | pegMaxFiniteMagOut;
  assign out[10] = N198 | pegMaxFiniteMagOut;
  assign out[9] = N197 | pegMaxFiniteMagOut;
  assign out[8] = N196 | pegMaxFiniteMagOut;
  assign out[7] = N195 | pegMaxFiniteMagOut;
  assign out[6] = N194 | pegMaxFiniteMagOut;
  assign out[5] = N193 | pegMaxFiniteMagOut;
  assign out[4] = N192 | pegMaxFiniteMagOut;
  assign out[3] = N191 | pegMaxFiniteMagOut;
  assign out[2] = N190 | pegMaxFiniteMagOut;
  assign out[1] = N189 | pegMaxFiniteMagOut;
  assign out[0] = N188 | pegMaxFiniteMagOut;

endmodule



module recFNToRecFN_unsafe_inExpWidth8_inSigWidth24_outExpWidth11_outSigWidth53
(
  in,
  out
);

  input [32:0] in;
  output [64:0] out;
  wire [64:0] out;
  wire N0,N1,N2,N3,isNaN,isInf,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45;
  assign out[0] = 1'b0;
  assign out[1] = 1'b0;
  assign out[2] = 1'b0;
  assign out[3] = 1'b0;
  assign out[4] = 1'b0;
  assign out[5] = 1'b0;
  assign out[6] = 1'b0;
  assign out[7] = 1'b0;
  assign out[8] = 1'b0;
  assign out[9] = 1'b0;
  assign out[10] = 1'b0;
  assign out[11] = 1'b0;
  assign out[12] = 1'b0;
  assign out[13] = 1'b0;
  assign out[14] = 1'b0;
  assign out[15] = 1'b0;
  assign out[16] = 1'b0;
  assign out[17] = 1'b0;
  assign out[18] = 1'b0;
  assign out[19] = 1'b0;
  assign out[20] = 1'b0;
  assign out[21] = 1'b0;
  assign out[22] = 1'b0;
  assign out[23] = 1'b0;
  assign out[24] = 1'b0;
  assign out[25] = 1'b0;
  assign out[26] = 1'b0;
  assign out[27] = 1'b0;
  assign out[28] = 1'b0;
  assign N41 = in[30] | in[31];
  assign N42 = in[29] | N41;
  assign N43 = ~N42;
  assign N44 = in[30] & in[31];
  assign { N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15 } = in[31:23] + { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign out[51:29] = (N0)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                      (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                      (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                      (N6)? in[22:0] : 1'b0;
  assign N0 = isNaN;
  assign { N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27 } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N2)? { N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15 } : 1'b0;
  assign N1 = N43;
  assign N2 = N42;
  assign out[63:52] = (N0)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                      (N39)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                      (N13)? { N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27 } : 1'b0;
  assign out[64] = (N0)? 1'b0 : 
                   (N3)? in[32] : 1'b0;
  assign N3 = N40;
  assign isNaN = N44 & in[29];
  assign isInf = N44 & N45;
  assign N45 = ~in[29];
  assign N4 = isInf | isNaN;
  assign N5 = N43 | N4;
  assign N6 = ~N5;
  assign N7 = ~isNaN;
  assign N8 = isInf & N7;
  assign N9 = ~isInf;
  assign N10 = N7 & N9;
  assign N11 = N43 & N10;
  assign N12 = isInf | isNaN;
  assign N13 = ~N12;
  assign N14 = N13;
  assign N39 = isInf & N7;
  assign N40 = ~isNaN;

endmodule



module roundRawFNtoRecFN_mixed_fullExpWidth11_fullSigWidth53_midExpWidth8_midSigWidth24_outExpWidth11_outSigWidth53
(
  control,
  invalidExc,
  infiniteExc,
  in_isNaN,
  in_isInf,
  in_isZero,
  in_sign,
  in_sExp,
  in_sig,
  roundingMode,
  fullOut,
  fullExceptionFlags,
  midOut,
  midExceptionFlags
);

  input [0:0] control;
  input [12:0] in_sExp;
  input [55:0] in_sig;
  input [2:0] roundingMode;
  output [64:0] fullOut;
  output [4:0] fullExceptionFlags;
  output [64:0] midOut;
  output [4:0] midExceptionFlags;
  input invalidExc;
  input infiniteExc;
  input in_isNaN;
  input in_isInf;
  input in_isZero;
  input in_sign;
  wire [64:0] fullOut,midOut;
  wire [4:0] fullExceptionFlags,midExceptionFlags;
  wire [32:0] midResult;

  roundAnyRawFNToRecFN_inExpWidth11_inSigWidth55_outExpWidth11_outSigWidth53
  round64
  (
    .control(control[0]),
    .invalidExc(invalidExc),
    .infiniteExc(infiniteExc),
    .in_isNaN(in_isNaN),
    .in_isInf(in_isInf),
    .in_isZero(in_isZero),
    .in_sign(in_sign),
    .in_sExp(in_sExp),
    .in_sig(in_sig),
    .roundingMode(roundingMode),
    .out(fullOut),
    .exceptionFlags(fullExceptionFlags)
  );


  roundAnyRawFNToRecFN_inExpWidth11_inSigWidth55_outExpWidth8_outSigWidth24
  round32
  (
    .control(control[0]),
    .invalidExc(invalidExc),
    .infiniteExc(infiniteExc),
    .in_isNaN(in_isNaN),
    .in_isInf(in_isInf),
    .in_isZero(in_isZero),
    .in_sign(in_sign),
    .in_sExp(in_sExp),
    .in_sig(in_sig),
    .roundingMode(roundingMode),
    .out(midResult),
    .exceptionFlags(midExceptionFlags)
  );


  recFNToRecFN_unsafe_inExpWidth8_inSigWidth24_outExpWidth11_outSigWidth53
  recover
  (
    .in(midResult),
    .out(midOut)
  );


endmodule



module bp_be_fp_rebox_00
(
  raw_i,
  tag_i,
  frm_i,
  invalid_exc_i,
  infinite_exc_i,
  reg_o,
  fflags_o
);

  input [74:0] raw_i;
  input [0:0] tag_i;
  input [2:0] frm_i;
  output [65:0] reg_o;
  output [4:0] fflags_o;
  input invalid_exc_i;
  input infinite_exc_i;
  wire [65:0] reg_o;
  wire [4:0] fflags_o;
  wire N0,N1,fflags_dp_nv_,fflags_dp_dz_,fflags_dp_of_,fflags_dp_uf_,fflags_dp_nx_,
  fflags_sp_nv_,fflags_sp_dz_,fflags_sp_of_,fflags_sp_uf_,fflags_sp_nx_,N2;
  wire [64:0] result_dp,result_sp;

  roundRawFNtoRecFN_mixed_fullExpWidth11_fullSigWidth53_midExpWidth8_midSigWidth24_outExpWidth11_outSigWidth53
  round_mixed
  (
    .control(1'b1),
    .invalidExc(invalid_exc_i),
    .infiniteExc(infinite_exc_i),
    .in_isNaN(raw_i[74]),
    .in_isInf(raw_i[73]),
    .in_isZero(raw_i[72]),
    .in_sign(raw_i[69]),
    .in_sExp(raw_i[68:56]),
    .in_sig(raw_i[55:0]),
    .roundingMode(frm_i),
    .fullOut(result_dp),
    .fullExceptionFlags({ fflags_dp_nv_, fflags_dp_dz_, fflags_dp_of_, fflags_dp_uf_, fflags_dp_nx_ }),
    .midOut(result_sp),
    .midExceptionFlags({ fflags_sp_nv_, fflags_sp_dz_, fflags_sp_of_, fflags_sp_uf_, fflags_sp_nx_ })
  );

  assign reg_o[64:0] = (N0)? result_sp : 
                       (N1)? result_dp : 1'b0;
  assign N0 = reg_o[65];
  assign N1 = N2;
  assign fflags_o = (N0)? { fflags_sp_nv_, fflags_sp_dz_, fflags_sp_of_, fflags_sp_uf_, fflags_sp_nx_ } : 
                    (N1)? { fflags_dp_nv_, fflags_dp_dz_, fflags_dp_of_, fflags_dp_uf_, fflags_dp_nx_ } : 1'b0;
  assign N2 = ~tag_i[0];
  assign reg_o[65] = tag_i[0];

endmodule



module bsg_dff_width_p72
(
  clk_i,
  data_i,
  data_o
);

  input [71:0] data_i;
  output [71:0] data_o;
  input clk_i;
  wire [71:0] data_o;
  reg data_o_71_sv2v_reg,data_o_70_sv2v_reg,data_o_69_sv2v_reg,data_o_68_sv2v_reg,
  data_o_67_sv2v_reg,data_o_66_sv2v_reg,data_o_65_sv2v_reg,data_o_64_sv2v_reg,
  data_o_63_sv2v_reg,data_o_62_sv2v_reg,data_o_61_sv2v_reg,data_o_60_sv2v_reg,
  data_o_59_sv2v_reg,data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,
  data_o_55_sv2v_reg,data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,data_o_51_sv2v_reg,
  data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,data_o_47_sv2v_reg,
  data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,data_o_43_sv2v_reg,
  data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,
  data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,
  data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,
  data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,
  data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,
  data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,
  data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,
  data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_chain_width_p72_num_stages_p1
(
  clk_i,
  data_i,
  data_o
);

  input [71:0] data_i;
  output [71:0] data_o;
  input clk_i;
  wire [71:0] data_o;

  bsg_dff_width_p72
  \chained.genblk1_1_.ch_reg 
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .data_o(data_o)
  );


endmodule



module bp_be_pipe_aux_00
(
  clk_i,
  reset_i,
  reservation_i,
  flush_i,
  frm_dyn_i,
  data_o,
  v_o,
  fflags_o_nv_,
  fflags_o_dz_,
  fflags_o_of_,
  fflags_o_uf_,
  fflags_o_nx_
);

  input [520:0] reservation_i;
  input [2:0] frm_dyn_i;
  output [65:0] data_o;
  input clk_i;
  input reset_i;
  input flush_i;
  output v_o;
  output fflags_o_nv_;
  output fflags_o_dz_;
  output fflags_o_of_;
  output fflags_o_uf_;
  output fflags_o_nx_;
  wire [65:0] data_o,ieee_data_lo,rebox_data_lo,frd_data_lo,ird_data_lo,aux_result;
  wire v_o,fflags_o_nv_,fflags_o_dz_,fflags_o_of_,fflags_o_uf_,fflags_o_nx_,N0,N1,N2,
  N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,
  N25,N26,N27,N28,fclass_result_q_nan_,fclass_result_s_nan_,fclass_result_p_inf_,
  fclass_result_p_norm_,fclass_result_p_sub_,fclass_result_p_zero_,
  fclass_result_n_zero_,fclass_result_n_sub_,fclass_result_n_norm_,fclass_result_n_inf_,N29,N30,
  N31,N32,N33,N34,irs1_unsigned,_2_net_,i2f_fflags_nv_,i2f_fflags_dz_,i2f_fflags_of_,
  i2f_fflags_uf_,i2f_fflags_nx_,i2f_result_is_nan_,i2f_result_is_inf_,
  i2f_result_is_zero_,i2f_result_sign_,i2f_result_sexp__12_,i2f_result_sexp__11_,
  i2f_result_sexp__10_,i2f_result_sexp__9_,i2f_result_sexp__8_,i2f_result_sexp__7_,
  i2f_result_sexp__6_,i2f_result_sexp__5_,i2f_result_sexp__4_,i2f_result_sexp__3_,
  i2f_result_sexp__2_,i2f_result_sexp__1_,i2f_result_sexp__0_,N35,N36,N37,N38,N39,N40,
  signed_f2i,f2dw_iflags_nv_,f2dw_iflags_of_,f2dw_iflags_nx_,dword_fflags_nv_,
  f2w_iflags_nv_,f2w_iflags_of_,f2w_iflags_nx_,word_fflags_nv_,f2i_fflags_nv_,f2i_fflags_nx_,
  invbox_frs1,invbox_frs2,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,
  N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,
  N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,
  N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,
  N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,
  N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,
  N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,
  N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,
  N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,
  N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,
  N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,
  N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,
  N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,
  N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,
  N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,
  N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,
  N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,
  N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,
  N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
  N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,
  N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,
  N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,
  N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,
  N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,
  N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,
  N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,
  N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,
  N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,
  N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,
  N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,
  N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,
  N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,
  N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,
  N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,
  N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,
  N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,
  N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,
  N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,
  N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,
  N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,
  N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
  N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,
  N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,
  N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,
  N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,
  N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,
  N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,
  N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,
  N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,
  N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,
  N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,
  N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,
  N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,
  N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,
  N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,
  N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,
  N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,
  N960,N961,N962,N963,N964,N965,signaling_li,flt_lo,feq_lo,fgt_lo,unordered_lo,
  fcmp_fflags_nv_,fcmp_fflags_dz_,fcmp_fflags_of_,fcmp_fflags_uf_,fcmp_fflags_nx_,
  fcmp_out,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,
  N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,
  N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,
  N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,
  N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,
  N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,
  N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,
  N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,
  N1077,N1078,N1079,raw_fflags_nv_,raw_fflags_dz_,raw_fflags_of_,raw_fflags_uf_,
  raw_fflags_nx_,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,
  N1158,N1159,rebox_fflags_nv_,rebox_fflags_dz_,rebox_fflags_of_,rebox_fflags_uf_,
  rebox_fflags_nx_,N1160,frd_fflags_nv_,frd_fflags_dz_,frd_fflags_of_,
  frd_fflags_uf_,frd_fflags_nx_,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,
  N1198,N1199,N1200,ird_fflags_nv_,ird_fflags_dz_,ird_fflags_of_,ird_fflags_uf_,
  ird_fflags_nx_,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,N1211,
  N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,N1238,
  N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,N1251,
  N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,aux_v_li,N1271,N1272,N1273,N1274,N1275,N1276,
  N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,
  N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
  N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,
  N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,
  N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,
  N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,
  N1397,N1398,N1399,N1400,N1401,N1402;
  wire [2:0] frm_li;
  wire [74:0] frs1_raw,frs2_raw,fminmax_result,raw_result;
  wire [64:0] i2f_rec;
  wire [53:0] i2f_sig;
  wire [63:0] f2dw_out,f2i_result,imvf_result,fsgnj_a,fsgnj_b,fsgnj_result,ieee_result,
  iaux_result;
  wire [31:0] f2w_out;
  wire [4:0] aux_fflags;

  bp_be_rec_to_raw_00
  frs1_to_raw
  (
    .rec_i(reservation_i[194:130]),
    .tag_i(reservation_i[412]),
    .raw_o(frs1_raw)
  );


  bp_be_rec_to_raw_00
  frs2_to_raw
  (
    .rec_i(reservation_i[129:65]),
    .tag_i(reservation_i[411]),
    .raw_o(frs2_raw)
  );

  assign N29 = ~reservation_i[406];
  assign N30 = reservation_i[408] | reservation_i[409];
  assign N31 = reservation_i[407] | N30;
  assign N32 = N29 | N31;
  assign N33 = reservation_i[405] | N32;
  assign N34 = reservation_i[404] | N33;
  assign irs1_unsigned = ~N34;

  iNToRecFN_intWidth64_expWidth11_sigWidth53
  i2f
  (
    .control(1'b1),
    .signedIn(_2_net_),
    .in(reservation_i[388:325]),
    .roundingMode(frm_li),
    .out(i2f_rec),
    .exceptionFlags({ i2f_fflags_nv_, i2f_fflags_dz_, i2f_fflags_of_, i2f_fflags_uf_, i2f_fflags_nx_ })
  );


  recFNToRawFN_expWidth11_sigWidth53
  i2f_rec_to_raw
  (
    .in(i2f_rec),
    .isNaN(i2f_result_is_nan_),
    .isInf(i2f_result_is_inf_),
    .isZero(i2f_result_is_zero_),
    .sign(i2f_result_sign_),
    .sExp({ i2f_result_sexp__12_, i2f_result_sexp__11_, i2f_result_sexp__10_, i2f_result_sexp__9_, i2f_result_sexp__8_, i2f_result_sexp__7_, i2f_result_sexp__6_, i2f_result_sexp__5_, i2f_result_sexp__4_, i2f_result_sexp__3_, i2f_result_sexp__2_, i2f_result_sexp__1_, i2f_result_sexp__0_ }),
    .sig(i2f_sig)
  );

  assign N35 = ~reservation_i[404];
  assign N36 = reservation_i[408] | reservation_i[409];
  assign N37 = reservation_i[407] | N36;
  assign N38 = reservation_i[406] | N37;
  assign N39 = reservation_i[405] | N38;
  assign N40 = N35 | N39;
  assign signed_f2i = ~N40;

  recFNToIN_expWidth11_sigWidth53_intWidth64
  f2dw
  (
    .control(1'b1),
    .in(reservation_i[194:130]),
    .roundingMode(frm_li),
    .signedOut(signed_f2i),
    .out(f2dw_out),
    .intExceptionFlags({ f2dw_iflags_nv_, f2dw_iflags_of_, f2dw_iflags_nx_ })
  );


  recFNToIN_expWidth11_sigWidth53_intWidth32
  f2w
  (
    .control(1'b1),
    .in(reservation_i[194:130]),
    .roundingMode(frm_li),
    .signedOut(signed_f2i),
    .out(f2w_out),
    .intExceptionFlags({ f2w_iflags_nv_, f2w_iflags_of_, f2w_iflags_nx_ })
  );

  assign N43 = reservation_i[409] | reservation_i[408];
  assign N44 = N1273 | reservation_i[406];
  assign N45 = reservation_i[405] | reservation_i[404];
  assign N46 = N43 | N44;
  assign N47 = N46 | N45;
  assign N49 = reservation_i[409] | reservation_i[408];
  assign N50 = N1273 | reservation_i[406];
  assign N51 = reservation_i[405] | N35;
  assign N52 = N49 | N50;
  assign N53 = N52 | N51;
  assign N55 = reservation_i[409] | reservation_i[408];
  assign N56 = reservation_i[407] | N29;
  assign N57 = N1274 | N35;
  assign N58 = N55 | N56;
  assign N59 = N58 | N57;
  assign N194 = (N130)? fsgnj_b[0] : 
                (N132)? fsgnj_b[1] : 
                (N134)? fsgnj_b[2] : 
                (N136)? fsgnj_b[3] : 
                (N138)? fsgnj_b[4] : 
                (N140)? fsgnj_b[5] : 
                (N142)? fsgnj_b[6] : 
                (N144)? fsgnj_b[7] : 
                (N146)? fsgnj_b[8] : 
                (N148)? fsgnj_b[9] : 
                (N150)? fsgnj_b[10] : 
                (N152)? fsgnj_b[11] : 
                (N154)? fsgnj_b[12] : 
                (N156)? fsgnj_b[13] : 
                (N158)? fsgnj_b[14] : 
                (N160)? fsgnj_b[15] : 
                (N162)? fsgnj_b[16] : 
                (N164)? fsgnj_b[17] : 
                (N166)? fsgnj_b[18] : 
                (N168)? fsgnj_b[19] : 
                (N170)? fsgnj_b[20] : 
                (N172)? fsgnj_b[21] : 
                (N174)? fsgnj_b[22] : 
                (N176)? fsgnj_b[23] : 
                (N178)? fsgnj_b[24] : 
                (N180)? fsgnj_b[25] : 
                (N182)? fsgnj_b[26] : 
                (N184)? fsgnj_b[27] : 
                (N186)? fsgnj_b[28] : 
                (N188)? fsgnj_b[29] : 
                (N190)? fsgnj_b[30] : 
                (N192)? fsgnj_b[31] : 
                (N131)? fsgnj_b[32] : 
                (N133)? fsgnj_b[33] : 
                (N135)? fsgnj_b[34] : 
                (N137)? fsgnj_b[35] : 
                (N139)? fsgnj_b[36] : 
                (N141)? fsgnj_b[37] : 
                (N143)? fsgnj_b[38] : 
                (N145)? fsgnj_b[39] : 
                (N147)? fsgnj_b[40] : 
                (N149)? fsgnj_b[41] : 
                (N151)? fsgnj_b[42] : 
                (N153)? fsgnj_b[43] : 
                (N155)? fsgnj_b[44] : 
                (N157)? fsgnj_b[45] : 
                (N159)? fsgnj_b[46] : 
                (N161)? fsgnj_b[47] : 
                (N163)? fsgnj_b[48] : 
                (N165)? fsgnj_b[49] : 
                (N167)? fsgnj_b[50] : 
                (N169)? fsgnj_b[51] : 
                (N171)? fsgnj_b[52] : 
                (N173)? fsgnj_b[53] : 
                (N175)? fsgnj_b[54] : 
                (N177)? fsgnj_b[55] : 
                (N179)? fsgnj_b[56] : 
                (N181)? fsgnj_b[57] : 
                (N183)? fsgnj_b[58] : 
                (N185)? fsgnj_b[59] : 
                (N187)? fsgnj_b[60] : 
                (N189)? fsgnj_b[61] : 
                (N191)? fsgnj_b[62] : 
                (N193)? fsgnj_b[63] : 1'b0;
  assign N452 = (N388)? fsgnj_b[0] : 
                (N390)? fsgnj_b[1] : 
                (N392)? fsgnj_b[2] : 
                (N394)? fsgnj_b[3] : 
                (N396)? fsgnj_b[4] : 
                (N398)? fsgnj_b[5] : 
                (N400)? fsgnj_b[6] : 
                (N402)? fsgnj_b[7] : 
                (N404)? fsgnj_b[8] : 
                (N406)? fsgnj_b[9] : 
                (N408)? fsgnj_b[10] : 
                (N410)? fsgnj_b[11] : 
                (N412)? fsgnj_b[12] : 
                (N414)? fsgnj_b[13] : 
                (N416)? fsgnj_b[14] : 
                (N418)? fsgnj_b[15] : 
                (N420)? fsgnj_b[16] : 
                (N422)? fsgnj_b[17] : 
                (N424)? fsgnj_b[18] : 
                (N426)? fsgnj_b[19] : 
                (N428)? fsgnj_b[20] : 
                (N430)? fsgnj_b[21] : 
                (N432)? fsgnj_b[22] : 
                (N434)? fsgnj_b[23] : 
                (N436)? fsgnj_b[24] : 
                (N438)? fsgnj_b[25] : 
                (N440)? fsgnj_b[26] : 
                (N442)? fsgnj_b[27] : 
                (N444)? fsgnj_b[28] : 
                (N446)? fsgnj_b[29] : 
                (N448)? fsgnj_b[30] : 
                (N450)? fsgnj_b[31] : 
                (N389)? fsgnj_b[32] : 
                (N391)? fsgnj_b[33] : 
                (N393)? fsgnj_b[34] : 
                (N395)? fsgnj_b[35] : 
                (N397)? fsgnj_b[36] : 
                (N399)? fsgnj_b[37] : 
                (N401)? fsgnj_b[38] : 
                (N403)? fsgnj_b[39] : 
                (N405)? fsgnj_b[40] : 
                (N407)? fsgnj_b[41] : 
                (N409)? fsgnj_b[42] : 
                (N411)? fsgnj_b[43] : 
                (N413)? fsgnj_b[44] : 
                (N415)? fsgnj_b[45] : 
                (N417)? fsgnj_b[46] : 
                (N419)? fsgnj_b[47] : 
                (N421)? fsgnj_b[48] : 
                (N423)? fsgnj_b[49] : 
                (N425)? fsgnj_b[50] : 
                (N427)? fsgnj_b[51] : 
                (N429)? fsgnj_b[52] : 
                (N431)? fsgnj_b[53] : 
                (N433)? fsgnj_b[54] : 
                (N435)? fsgnj_b[55] : 
                (N437)? fsgnj_b[56] : 
                (N439)? fsgnj_b[57] : 
                (N441)? fsgnj_b[58] : 
                (N443)? fsgnj_b[59] : 
                (N445)? fsgnj_b[60] : 
                (N447)? fsgnj_b[61] : 
                (N449)? fsgnj_b[62] : 
                (N451)? fsgnj_b[63] : 1'b0;
  assign N582 = (N518)? fsgnj_a[0] : 
                (N520)? fsgnj_a[1] : 
                (N522)? fsgnj_a[2] : 
                (N524)? fsgnj_a[3] : 
                (N526)? fsgnj_a[4] : 
                (N528)? fsgnj_a[5] : 
                (N530)? fsgnj_a[6] : 
                (N532)? fsgnj_a[7] : 
                (N534)? fsgnj_a[8] : 
                (N536)? fsgnj_a[9] : 
                (N538)? fsgnj_a[10] : 
                (N540)? fsgnj_a[11] : 
                (N542)? fsgnj_a[12] : 
                (N544)? fsgnj_a[13] : 
                (N546)? fsgnj_a[14] : 
                (N548)? fsgnj_a[15] : 
                (N550)? fsgnj_a[16] : 
                (N552)? fsgnj_a[17] : 
                (N554)? fsgnj_a[18] : 
                (N556)? fsgnj_a[19] : 
                (N558)? fsgnj_a[20] : 
                (N560)? fsgnj_a[21] : 
                (N562)? fsgnj_a[22] : 
                (N564)? fsgnj_a[23] : 
                (N566)? fsgnj_a[24] : 
                (N568)? fsgnj_a[25] : 
                (N570)? fsgnj_a[26] : 
                (N572)? fsgnj_a[27] : 
                (N574)? fsgnj_a[28] : 
                (N576)? fsgnj_a[29] : 
                (N578)? fsgnj_a[30] : 
                (N580)? fsgnj_a[31] : 
                (N519)? fsgnj_a[32] : 
                (N521)? fsgnj_a[33] : 
                (N523)? fsgnj_a[34] : 
                (N525)? fsgnj_a[35] : 
                (N527)? fsgnj_a[36] : 
                (N529)? fsgnj_a[37] : 
                (N531)? fsgnj_a[38] : 
                (N533)? fsgnj_a[39] : 
                (N535)? fsgnj_a[40] : 
                (N537)? fsgnj_a[41] : 
                (N539)? fsgnj_a[42] : 
                (N541)? fsgnj_a[43] : 
                (N543)? fsgnj_a[44] : 
                (N545)? fsgnj_a[45] : 
                (N547)? fsgnj_a[46] : 
                (N549)? fsgnj_a[47] : 
                (N551)? fsgnj_a[48] : 
                (N553)? fsgnj_a[49] : 
                (N555)? fsgnj_a[50] : 
                (N557)? fsgnj_a[51] : 
                (N559)? fsgnj_a[52] : 
                (N561)? fsgnj_a[53] : 
                (N563)? fsgnj_a[54] : 
                (N565)? fsgnj_a[55] : 
                (N567)? fsgnj_a[56] : 
                (N569)? fsgnj_a[57] : 
                (N571)? fsgnj_a[58] : 
                (N573)? fsgnj_a[59] : 
                (N575)? fsgnj_a[60] : 
                (N577)? fsgnj_a[61] : 
                (N579)? fsgnj_a[62] : 
                (N581)? fsgnj_a[63] : 1'b0;
  assign N839 = (N775)? fsgnj_b[0] : 
                (N777)? fsgnj_b[1] : 
                (N779)? fsgnj_b[2] : 
                (N781)? fsgnj_b[3] : 
                (N783)? fsgnj_b[4] : 
                (N785)? fsgnj_b[5] : 
                (N787)? fsgnj_b[6] : 
                (N789)? fsgnj_b[7] : 
                (N791)? fsgnj_b[8] : 
                (N793)? fsgnj_b[9] : 
                (N795)? fsgnj_b[10] : 
                (N797)? fsgnj_b[11] : 
                (N799)? fsgnj_b[12] : 
                (N801)? fsgnj_b[13] : 
                (N803)? fsgnj_b[14] : 
                (N805)? fsgnj_b[15] : 
                (N807)? fsgnj_b[16] : 
                (N809)? fsgnj_b[17] : 
                (N811)? fsgnj_b[18] : 
                (N813)? fsgnj_b[19] : 
                (N815)? fsgnj_b[20] : 
                (N817)? fsgnj_b[21] : 
                (N819)? fsgnj_b[22] : 
                (N821)? fsgnj_b[23] : 
                (N823)? fsgnj_b[24] : 
                (N825)? fsgnj_b[25] : 
                (N827)? fsgnj_b[26] : 
                (N829)? fsgnj_b[27] : 
                (N831)? fsgnj_b[28] : 
                (N833)? fsgnj_b[29] : 
                (N835)? fsgnj_b[30] : 
                (N837)? fsgnj_b[31] : 
                (N776)? fsgnj_b[32] : 
                (N778)? fsgnj_b[33] : 
                (N780)? fsgnj_b[34] : 
                (N782)? fsgnj_b[35] : 
                (N784)? fsgnj_b[36] : 
                (N786)? fsgnj_b[37] : 
                (N788)? fsgnj_b[38] : 
                (N790)? fsgnj_b[39] : 
                (N792)? fsgnj_b[40] : 
                (N794)? fsgnj_b[41] : 
                (N796)? fsgnj_b[42] : 
                (N798)? fsgnj_b[43] : 
                (N800)? fsgnj_b[44] : 
                (N802)? fsgnj_b[45] : 
                (N804)? fsgnj_b[46] : 
                (N806)? fsgnj_b[47] : 
                (N808)? fsgnj_b[48] : 
                (N810)? fsgnj_b[49] : 
                (N812)? fsgnj_b[50] : 
                (N814)? fsgnj_b[51] : 
                (N816)? fsgnj_b[52] : 
                (N818)? fsgnj_b[53] : 
                (N820)? fsgnj_b[54] : 
                (N822)? fsgnj_b[55] : 
                (N824)? fsgnj_b[56] : 
                (N826)? fsgnj_b[57] : 
                (N828)? fsgnj_b[58] : 
                (N830)? fsgnj_b[59] : 
                (N832)? fsgnj_b[60] : 
                (N834)? fsgnj_b[61] : 
                (N836)? fsgnj_b[62] : 
                (N838)? fsgnj_b[63] : 1'b0;

  compareRecFN_expWidth11_sigWidth53
  fcmp
  (
    .a(reservation_i[194:130]),
    .b(reservation_i[129:65]),
    .signaling(signaling_li),
    .lt(flt_lo),
    .eq(feq_lo),
    .gt(fgt_lo),
    .unordered(unordered_lo),
    .exceptionFlags({ fcmp_fflags_nv_, fcmp_fflags_dz_, fcmp_fflags_of_, fcmp_fflags_uf_, fcmp_fflags_nx_ })
  );

  assign N1063 = reservation_i[409] | reservation_i[408];
  assign N1064 = reservation_i[407] | N29;
  assign N1065 = reservation_i[405] | N35;
  assign N1066 = N1063 | N1064;
  assign N1067 = N1066 | N1065;

  bp_be_fp_box_00
  fp_box
  (
    .ieee_i(ieee_result),
    .tag_i(reservation_i[403]),
    .reg_o(ieee_data_lo)
  );

  assign N1071 = N1069 & N1070;
  assign N1072 = N1273 & N35;
  assign N1073 = N1071 & N1072;
  assign N1075 = reservation_i[406] | N1274;
  assign N1076 = N29 | reservation_i[405];
  assign N1078 = N29 & N1274;
  assign N1079 = reservation_i[406] & reservation_i[405];

  bp_be_fp_rebox_00
  rebox
  (
    .raw_i(raw_result),
    .tag_i(reservation_i[403]),
    .frm_i(frm_li),
    .invalid_exc_i(1'b0),
    .infinite_exc_i(1'b0),
    .reg_o(rebox_data_lo),
    .fflags_o({ rebox_fflags_nv_, rebox_fflags_dz_, rebox_fflags_of_, rebox_fflags_uf_, rebox_fflags_nx_ })
  );

  assign N1166 = N1069 & N1070;
  assign N1168 = reservation_i[407] | N29;
  assign N1169 = N1274 | reservation_i[404];
  assign N1170 = N1168 | N1169;
  assign N1172 = reservation_i[407] | reservation_i[406];
  assign N1173 = reservation_i[405] | N35;
  assign N1174 = N1172 | N1173;
  assign N1175 = reservation_i[407] | reservation_i[406];
  assign N1176 = N1274 | N35;
  assign N1177 = N1175 | N1176;
  assign N1179 = N1273 | reservation_i[406];
  assign N1180 = N1274 | reservation_i[404];
  assign N1181 = N1179 | N1180;
  assign N1182 = N1273 | reservation_i[406];
  assign N1183 = N1274 | N35;
  assign N1184 = N1182 | N1183;
  assign N1185 = N1273 | N29;
  assign N1186 = reservation_i[405] | reservation_i[404];
  assign N1187 = N1185 | N1186;
  assign N1189 = reservation_i[406] & reservation_i[404];
  assign N1190 = reservation_i[407] & N1274;
  assign N1191 = N1190 & reservation_i[404];
  assign N1192 = reservation_i[407] & reservation_i[406];
  assign N1193 = N1192 & reservation_i[405];
  assign N1194 = N1273 & N29;
  assign N1195 = N1194 & N35;
  assign N1196 = N1273 & N1274;
  assign N1197 = N1196 & N35;
  assign N1198 = N29 & N1274;
  assign N1199 = N1198 & N35;

  bp_be_int_box_00
  int_box
  (
    .raw_i(iaux_result),
    .tag_i(reservation_i[402:401]),
    .unsigned_i(1'b0),
    .reg_o(ird_data_lo)
  );


  bsg_dff_chain_width_p72_num_stages_p1
  retiming_chain
  (
    .clk_i(clk_i),
    .data_i({ aux_fflags, aux_result, aux_v_li }),
    .data_o({ fflags_o_nv_, fflags_o_dz_, fflags_o_of_, fflags_o_uf_, fflags_o_nx_, data_o, v_o })
  );

  assign N1271 = reservation_i[462] & reservation_i[463];
  assign N1272 = reservation_i[461] & N1271;
  assign N1273 = ~reservation_i[407];
  assign N1274 = ~reservation_i[405];
  assign N1275 = reservation_i[408] | reservation_i[409];
  assign N1276 = N1273 | N1275;
  assign N1277 = reservation_i[406] | N1276;
  assign N1278 = N1274 | N1277;
  assign N1279 = reservation_i[404] | N1278;
  assign N1280 = ~N1279;
  assign N1281 = reservation_i[408] | reservation_i[409];
  assign N1282 = N1273 | N1281;
  assign N1283 = reservation_i[406] | N1282;
  assign N1284 = N1274 | N1283;
  assign N1285 = N35 | N1284;
  assign N1286 = ~N1285;
  assign N1287 = reservation_i[408] | reservation_i[409];
  assign N1288 = N1273 | N1287;
  assign N1289 = N29 | N1288;
  assign N1290 = reservation_i[405] | N1289;
  assign N1291 = reservation_i[404] | N1290;
  assign N1292 = ~N1291;
  assign N1293 = ~reservation_i[401];
  assign N1294 = N1293 | reservation_i[402];
  assign N1295 = ~N1294;
  assign N1296 = reservation_i[408] | reservation_i[409];
  assign N1297 = N1273 | N1296;
  assign N1298 = N29 | N1297;
  assign N1299 = N1274 | N1298;
  assign N1300 = reservation_i[404] | N1299;
  assign N1301 = ~N1300;
  assign N1302 = reservation_i[408] | reservation_i[409];
  assign N1303 = N1273 | N1302;
  assign N1304 = N29 | N1303;
  assign N1305 = reservation_i[405] | N1304;
  assign N1306 = N35 | N1305;
  assign N1307 = ~N1306;
  assign N1308 = ~reservation_i[403];
  assign N195 = ~N1308;
  assign frm_li = (N0)? frm_dyn_i : 
                  (N28)? reservation_i[463:461] : 1'b0;
  assign N0 = N1272;
  assign f2i_result = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, f2w_out } : 
                      (N2)? f2dw_out : 1'b0;
  assign N1 = N1295;
  assign N2 = N1294;
  assign { f2i_fflags_nv_, f2i_fflags_nx_ } = (N1)? { word_fflags_nv_, f2w_iflags_nx_ } : 
                                              (N2)? { dword_fflags_nv_, f2dw_iflags_nx_ } : 1'b0;
  assign fsgnj_a = (N3)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                   (N4)? reservation_i[193:130] : 1'b0;
  assign N3 = invbox_frs1;
  assign N4 = N41;
  assign fsgnj_b = (N5)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                   (N6)? reservation_i[128:65] : 1'b0;
  assign N5 = invbox_frs2;
  assign N6 = N42;
  assign N198 = (N7)? N196 : 
                (N197)? fsgnj_a[0] : 1'b0;
  assign N7 = 1'b0;
  assign N200 = (N7)? N196 : 
                (N199)? fsgnj_a[1] : 1'b0;
  assign N202 = (N7)? N196 : 
                (N201)? fsgnj_a[2] : 1'b0;
  assign N204 = (N7)? N196 : 
                (N203)? fsgnj_a[3] : 1'b0;
  assign N206 = (N7)? N196 : 
                (N205)? fsgnj_a[4] : 1'b0;
  assign N208 = (N7)? N196 : 
                (N207)? fsgnj_a[5] : 1'b0;
  assign N210 = (N7)? N196 : 
                (N209)? fsgnj_a[6] : 1'b0;
  assign N212 = (N7)? N196 : 
                (N211)? fsgnj_a[7] : 1'b0;
  assign N214 = (N7)? N196 : 
                (N213)? fsgnj_a[8] : 1'b0;
  assign N216 = (N7)? N196 : 
                (N215)? fsgnj_a[9] : 1'b0;
  assign N218 = (N7)? N196 : 
                (N217)? fsgnj_a[10] : 1'b0;
  assign N220 = (N7)? N196 : 
                (N219)? fsgnj_a[11] : 1'b0;
  assign N222 = (N7)? N196 : 
                (N221)? fsgnj_a[12] : 1'b0;
  assign N224 = (N7)? N196 : 
                (N223)? fsgnj_a[13] : 1'b0;
  assign N226 = (N7)? N196 : 
                (N225)? fsgnj_a[14] : 1'b0;
  assign N228 = (N7)? N196 : 
                (N227)? fsgnj_a[15] : 1'b0;
  assign N230 = (N7)? N196 : 
                (N229)? fsgnj_a[16] : 1'b0;
  assign N232 = (N7)? N196 : 
                (N231)? fsgnj_a[17] : 1'b0;
  assign N234 = (N7)? N196 : 
                (N233)? fsgnj_a[18] : 1'b0;
  assign N236 = (N7)? N196 : 
                (N235)? fsgnj_a[19] : 1'b0;
  assign N238 = (N7)? N196 : 
                (N237)? fsgnj_a[20] : 1'b0;
  assign N240 = (N7)? N196 : 
                (N239)? fsgnj_a[21] : 1'b0;
  assign N242 = (N7)? N196 : 
                (N241)? fsgnj_a[22] : 1'b0;
  assign N244 = (N7)? N196 : 
                (N243)? fsgnj_a[23] : 1'b0;
  assign N246 = (N7)? N196 : 
                (N245)? fsgnj_a[24] : 1'b0;
  assign N248 = (N7)? N196 : 
                (N247)? fsgnj_a[25] : 1'b0;
  assign N250 = (N7)? N196 : 
                (N249)? fsgnj_a[26] : 1'b0;
  assign N252 = (N7)? N196 : 
                (N251)? fsgnj_a[27] : 1'b0;
  assign N254 = (N7)? N196 : 
                (N253)? fsgnj_a[28] : 1'b0;
  assign N256 = (N7)? N196 : 
                (N255)? fsgnj_a[29] : 1'b0;
  assign N258 = (N7)? N196 : 
                (N257)? fsgnj_a[30] : 1'b0;
  assign N259 = (N8)? N196 : 
                (N9)? fsgnj_a[31] : 1'b0;
  assign N8 = N195;
  assign N9 = N1308;
  assign N261 = (N7)? N196 : 
                (N260)? fsgnj_a[32] : 1'b0;
  assign N263 = (N7)? N196 : 
                (N262)? fsgnj_a[33] : 1'b0;
  assign N265 = (N7)? N196 : 
                (N264)? fsgnj_a[34] : 1'b0;
  assign N267 = (N7)? N196 : 
                (N266)? fsgnj_a[35] : 1'b0;
  assign N269 = (N7)? N196 : 
                (N268)? fsgnj_a[36] : 1'b0;
  assign N271 = (N7)? N196 : 
                (N270)? fsgnj_a[37] : 1'b0;
  assign N273 = (N7)? N196 : 
                (N272)? fsgnj_a[38] : 1'b0;
  assign N275 = (N7)? N196 : 
                (N274)? fsgnj_a[39] : 1'b0;
  assign N277 = (N7)? N196 : 
                (N276)? fsgnj_a[40] : 1'b0;
  assign N279 = (N7)? N196 : 
                (N278)? fsgnj_a[41] : 1'b0;
  assign N281 = (N7)? N196 : 
                (N280)? fsgnj_a[42] : 1'b0;
  assign N283 = (N7)? N196 : 
                (N282)? fsgnj_a[43] : 1'b0;
  assign N285 = (N7)? N196 : 
                (N284)? fsgnj_a[44] : 1'b0;
  assign N287 = (N7)? N196 : 
                (N286)? fsgnj_a[45] : 1'b0;
  assign N289 = (N7)? N196 : 
                (N288)? fsgnj_a[46] : 1'b0;
  assign N291 = (N7)? N196 : 
                (N290)? fsgnj_a[47] : 1'b0;
  assign N293 = (N7)? N196 : 
                (N292)? fsgnj_a[48] : 1'b0;
  assign N295 = (N7)? N196 : 
                (N294)? fsgnj_a[49] : 1'b0;
  assign N297 = (N7)? N196 : 
                (N296)? fsgnj_a[50] : 1'b0;
  assign N299 = (N7)? N196 : 
                (N298)? fsgnj_a[51] : 1'b0;
  assign N301 = (N7)? N196 : 
                (N300)? fsgnj_a[52] : 1'b0;
  assign N303 = (N7)? N196 : 
                (N302)? fsgnj_a[53] : 1'b0;
  assign N305 = (N7)? N196 : 
                (N304)? fsgnj_a[54] : 1'b0;
  assign N307 = (N7)? N196 : 
                (N306)? fsgnj_a[55] : 1'b0;
  assign N309 = (N7)? N196 : 
                (N308)? fsgnj_a[56] : 1'b0;
  assign N311 = (N7)? N196 : 
                (N310)? fsgnj_a[57] : 1'b0;
  assign N313 = (N7)? N196 : 
                (N312)? fsgnj_a[58] : 1'b0;
  assign N315 = (N7)? N196 : 
                (N314)? fsgnj_a[59] : 1'b0;
  assign N317 = (N7)? N196 : 
                (N316)? fsgnj_a[60] : 1'b0;
  assign N319 = (N7)? N196 : 
                (N318)? fsgnj_a[61] : 1'b0;
  assign N321 = (N7)? N196 : 
                (N320)? fsgnj_a[62] : 1'b0;
  assign N322 = (N9)? N196 : 
                (N129)? fsgnj_a[63] : 1'b0;
  assign N585 = (N7)? N583 : 
                (N584)? fsgnj_a[0] : 1'b0;
  assign N587 = (N7)? N583 : 
                (N586)? fsgnj_a[1] : 1'b0;
  assign N589 = (N7)? N583 : 
                (N588)? fsgnj_a[2] : 1'b0;
  assign N591 = (N7)? N583 : 
                (N590)? fsgnj_a[3] : 1'b0;
  assign N593 = (N7)? N583 : 
                (N592)? fsgnj_a[4] : 1'b0;
  assign N595 = (N7)? N583 : 
                (N594)? fsgnj_a[5] : 1'b0;
  assign N597 = (N7)? N583 : 
                (N596)? fsgnj_a[6] : 1'b0;
  assign N599 = (N7)? N583 : 
                (N598)? fsgnj_a[7] : 1'b0;
  assign N601 = (N7)? N583 : 
                (N600)? fsgnj_a[8] : 1'b0;
  assign N603 = (N7)? N583 : 
                (N602)? fsgnj_a[9] : 1'b0;
  assign N605 = (N7)? N583 : 
                (N604)? fsgnj_a[10] : 1'b0;
  assign N607 = (N7)? N583 : 
                (N606)? fsgnj_a[11] : 1'b0;
  assign N609 = (N7)? N583 : 
                (N608)? fsgnj_a[12] : 1'b0;
  assign N611 = (N7)? N583 : 
                (N610)? fsgnj_a[13] : 1'b0;
  assign N613 = (N7)? N583 : 
                (N612)? fsgnj_a[14] : 1'b0;
  assign N615 = (N7)? N583 : 
                (N614)? fsgnj_a[15] : 1'b0;
  assign N617 = (N7)? N583 : 
                (N616)? fsgnj_a[16] : 1'b0;
  assign N619 = (N7)? N583 : 
                (N618)? fsgnj_a[17] : 1'b0;
  assign N621 = (N7)? N583 : 
                (N620)? fsgnj_a[18] : 1'b0;
  assign N623 = (N7)? N583 : 
                (N622)? fsgnj_a[19] : 1'b0;
  assign N625 = (N7)? N583 : 
                (N624)? fsgnj_a[20] : 1'b0;
  assign N627 = (N7)? N583 : 
                (N626)? fsgnj_a[21] : 1'b0;
  assign N629 = (N7)? N583 : 
                (N628)? fsgnj_a[22] : 1'b0;
  assign N631 = (N7)? N583 : 
                (N630)? fsgnj_a[23] : 1'b0;
  assign N633 = (N7)? N583 : 
                (N632)? fsgnj_a[24] : 1'b0;
  assign N635 = (N7)? N583 : 
                (N634)? fsgnj_a[25] : 1'b0;
  assign N637 = (N7)? N583 : 
                (N636)? fsgnj_a[26] : 1'b0;
  assign N639 = (N7)? N583 : 
                (N638)? fsgnj_a[27] : 1'b0;
  assign N641 = (N7)? N583 : 
                (N640)? fsgnj_a[28] : 1'b0;
  assign N643 = (N7)? N583 : 
                (N642)? fsgnj_a[29] : 1'b0;
  assign N645 = (N7)? N583 : 
                (N644)? fsgnj_a[30] : 1'b0;
  assign N646 = (N8)? N583 : 
                (N9)? fsgnj_a[31] : 1'b0;
  assign N648 = (N7)? N583 : 
                (N647)? fsgnj_a[32] : 1'b0;
  assign N650 = (N7)? N583 : 
                (N649)? fsgnj_a[33] : 1'b0;
  assign N652 = (N7)? N583 : 
                (N651)? fsgnj_a[34] : 1'b0;
  assign N654 = (N7)? N583 : 
                (N653)? fsgnj_a[35] : 1'b0;
  assign N656 = (N7)? N583 : 
                (N655)? fsgnj_a[36] : 1'b0;
  assign N658 = (N7)? N583 : 
                (N657)? fsgnj_a[37] : 1'b0;
  assign N660 = (N7)? N583 : 
                (N659)? fsgnj_a[38] : 1'b0;
  assign N662 = (N7)? N583 : 
                (N661)? fsgnj_a[39] : 1'b0;
  assign N664 = (N7)? N583 : 
                (N663)? fsgnj_a[40] : 1'b0;
  assign N666 = (N7)? N583 : 
                (N665)? fsgnj_a[41] : 1'b0;
  assign N668 = (N7)? N583 : 
                (N667)? fsgnj_a[42] : 1'b0;
  assign N670 = (N7)? N583 : 
                (N669)? fsgnj_a[43] : 1'b0;
  assign N672 = (N7)? N583 : 
                (N671)? fsgnj_a[44] : 1'b0;
  assign N674 = (N7)? N583 : 
                (N673)? fsgnj_a[45] : 1'b0;
  assign N676 = (N7)? N583 : 
                (N675)? fsgnj_a[46] : 1'b0;
  assign N678 = (N7)? N583 : 
                (N677)? fsgnj_a[47] : 1'b0;
  assign N680 = (N7)? N583 : 
                (N679)? fsgnj_a[48] : 1'b0;
  assign N682 = (N7)? N583 : 
                (N681)? fsgnj_a[49] : 1'b0;
  assign N684 = (N7)? N583 : 
                (N683)? fsgnj_a[50] : 1'b0;
  assign N686 = (N7)? N583 : 
                (N685)? fsgnj_a[51] : 1'b0;
  assign N688 = (N7)? N583 : 
                (N687)? fsgnj_a[52] : 1'b0;
  assign N690 = (N7)? N583 : 
                (N689)? fsgnj_a[53] : 1'b0;
  assign N692 = (N7)? N583 : 
                (N691)? fsgnj_a[54] : 1'b0;
  assign N694 = (N7)? N583 : 
                (N693)? fsgnj_a[55] : 1'b0;
  assign N696 = (N7)? N583 : 
                (N695)? fsgnj_a[56] : 1'b0;
  assign N698 = (N7)? N583 : 
                (N697)? fsgnj_a[57] : 1'b0;
  assign N700 = (N7)? N583 : 
                (N699)? fsgnj_a[58] : 1'b0;
  assign N702 = (N7)? N583 : 
                (N701)? fsgnj_a[59] : 1'b0;
  assign N704 = (N7)? N583 : 
                (N703)? fsgnj_a[60] : 1'b0;
  assign N706 = (N7)? N583 : 
                (N705)? fsgnj_a[61] : 1'b0;
  assign N708 = (N7)? N583 : 
                (N707)? fsgnj_a[62] : 1'b0;
  assign N709 = (N9)? N583 : 
                (N129)? fsgnj_a[63] : 1'b0;
  assign N841 = (N7)? N839 : 
                (N840)? fsgnj_a[0] : 1'b0;
  assign N843 = (N7)? N839 : 
                (N842)? fsgnj_a[1] : 1'b0;
  assign N845 = (N7)? N839 : 
                (N844)? fsgnj_a[2] : 1'b0;
  assign N847 = (N7)? N839 : 
                (N846)? fsgnj_a[3] : 1'b0;
  assign N849 = (N7)? N839 : 
                (N848)? fsgnj_a[4] : 1'b0;
  assign N851 = (N7)? N839 : 
                (N850)? fsgnj_a[5] : 1'b0;
  assign N853 = (N7)? N839 : 
                (N852)? fsgnj_a[6] : 1'b0;
  assign N855 = (N7)? N839 : 
                (N854)? fsgnj_a[7] : 1'b0;
  assign N857 = (N7)? N839 : 
                (N856)? fsgnj_a[8] : 1'b0;
  assign N859 = (N7)? N839 : 
                (N858)? fsgnj_a[9] : 1'b0;
  assign N861 = (N7)? N839 : 
                (N860)? fsgnj_a[10] : 1'b0;
  assign N863 = (N7)? N839 : 
                (N862)? fsgnj_a[11] : 1'b0;
  assign N865 = (N7)? N839 : 
                (N864)? fsgnj_a[12] : 1'b0;
  assign N867 = (N7)? N839 : 
                (N866)? fsgnj_a[13] : 1'b0;
  assign N869 = (N7)? N839 : 
                (N868)? fsgnj_a[14] : 1'b0;
  assign N871 = (N7)? N839 : 
                (N870)? fsgnj_a[15] : 1'b0;
  assign N873 = (N7)? N839 : 
                (N872)? fsgnj_a[16] : 1'b0;
  assign N875 = (N7)? N839 : 
                (N874)? fsgnj_a[17] : 1'b0;
  assign N877 = (N7)? N839 : 
                (N876)? fsgnj_a[18] : 1'b0;
  assign N879 = (N7)? N839 : 
                (N878)? fsgnj_a[19] : 1'b0;
  assign N881 = (N7)? N839 : 
                (N880)? fsgnj_a[20] : 1'b0;
  assign N883 = (N7)? N839 : 
                (N882)? fsgnj_a[21] : 1'b0;
  assign N885 = (N7)? N839 : 
                (N884)? fsgnj_a[22] : 1'b0;
  assign N887 = (N7)? N839 : 
                (N886)? fsgnj_a[23] : 1'b0;
  assign N889 = (N7)? N839 : 
                (N888)? fsgnj_a[24] : 1'b0;
  assign N891 = (N7)? N839 : 
                (N890)? fsgnj_a[25] : 1'b0;
  assign N893 = (N7)? N839 : 
                (N892)? fsgnj_a[26] : 1'b0;
  assign N895 = (N7)? N839 : 
                (N894)? fsgnj_a[27] : 1'b0;
  assign N897 = (N7)? N839 : 
                (N896)? fsgnj_a[28] : 1'b0;
  assign N899 = (N7)? N839 : 
                (N898)? fsgnj_a[29] : 1'b0;
  assign N901 = (N7)? N839 : 
                (N900)? fsgnj_a[30] : 1'b0;
  assign N902 = (N8)? N839 : 
                (N9)? fsgnj_a[31] : 1'b0;
  assign N904 = (N7)? N839 : 
                (N903)? fsgnj_a[32] : 1'b0;
  assign N906 = (N7)? N839 : 
                (N905)? fsgnj_a[33] : 1'b0;
  assign N908 = (N7)? N839 : 
                (N907)? fsgnj_a[34] : 1'b0;
  assign N910 = (N7)? N839 : 
                (N909)? fsgnj_a[35] : 1'b0;
  assign N912 = (N7)? N839 : 
                (N911)? fsgnj_a[36] : 1'b0;
  assign N914 = (N7)? N839 : 
                (N913)? fsgnj_a[37] : 1'b0;
  assign N916 = (N7)? N839 : 
                (N915)? fsgnj_a[38] : 1'b0;
  assign N918 = (N7)? N839 : 
                (N917)? fsgnj_a[39] : 1'b0;
  assign N920 = (N7)? N839 : 
                (N919)? fsgnj_a[40] : 1'b0;
  assign N922 = (N7)? N839 : 
                (N921)? fsgnj_a[41] : 1'b0;
  assign N924 = (N7)? N839 : 
                (N923)? fsgnj_a[42] : 1'b0;
  assign N926 = (N7)? N839 : 
                (N925)? fsgnj_a[43] : 1'b0;
  assign N928 = (N7)? N839 : 
                (N927)? fsgnj_a[44] : 1'b0;
  assign N930 = (N7)? N839 : 
                (N929)? fsgnj_a[45] : 1'b0;
  assign N932 = (N7)? N839 : 
                (N931)? fsgnj_a[46] : 1'b0;
  assign N934 = (N7)? N839 : 
                (N933)? fsgnj_a[47] : 1'b0;
  assign N936 = (N7)? N839 : 
                (N935)? fsgnj_a[48] : 1'b0;
  assign N938 = (N7)? N839 : 
                (N937)? fsgnj_a[49] : 1'b0;
  assign N940 = (N7)? N839 : 
                (N939)? fsgnj_a[50] : 1'b0;
  assign N942 = (N7)? N839 : 
                (N941)? fsgnj_a[51] : 1'b0;
  assign N944 = (N7)? N839 : 
                (N943)? fsgnj_a[52] : 1'b0;
  assign N946 = (N7)? N839 : 
                (N945)? fsgnj_a[53] : 1'b0;
  assign N948 = (N7)? N839 : 
                (N947)? fsgnj_a[54] : 1'b0;
  assign N950 = (N7)? N839 : 
                (N949)? fsgnj_a[55] : 1'b0;
  assign N952 = (N7)? N839 : 
                (N951)? fsgnj_a[56] : 1'b0;
  assign N954 = (N7)? N839 : 
                (N953)? fsgnj_a[57] : 1'b0;
  assign N956 = (N7)? N839 : 
                (N955)? fsgnj_a[58] : 1'b0;
  assign N958 = (N7)? N839 : 
                (N957)? fsgnj_a[59] : 1'b0;
  assign N960 = (N7)? N839 : 
                (N959)? fsgnj_a[60] : 1'b0;
  assign N962 = (N7)? N839 : 
                (N961)? fsgnj_a[61] : 1'b0;
  assign N964 = (N7)? N839 : 
                (N963)? fsgnj_a[62] : 1'b0;
  assign N965 = (N9)? N839 : 
                (N129)? fsgnj_a[63] : 1'b0;
  assign fsgnj_result = (N10)? { N322, N321, N319, N317, N315, N313, N311, N309, N307, N305, N303, N301, N299, N297, N295, N293, N291, N289, N287, N285, N283, N281, N279, N277, N275, N273, N271, N269, N267, N265, N263, N261, N259, N258, N256, N254, N252, N250, N248, N246, N244, N242, N240, N238, N236, N234, N232, N230, N228, N226, N224, N222, N220, N218, N216, N214, N212, N210, N208, N206, N204, N202, N200, N198 } : 
                        (N11)? { N709, N708, N706, N704, N702, N700, N698, N696, N694, N692, N690, N688, N686, N684, N682, N680, N678, N676, N674, N672, N670, N668, N666, N664, N662, N660, N658, N656, N654, N652, N650, N648, N646, N645, N643, N641, N639, N637, N635, N633, N631, N629, N627, N625, N623, N621, N619, N617, N615, N613, N611, N609, N607, N605, N603, N601, N599, N597, N595, N593, N591, N589, N587, N585 } : 
                        (N12)? { N965, N964, N962, N960, N958, N956, N954, N952, N950, N948, N946, N944, N942, N940, N938, N936, N934, N932, N930, N928, N926, N924, N922, N920, N918, N916, N914, N912, N910, N908, N906, N904, N902, N901, N899, N897, N895, N893, N891, N889, N887, N885, N883, N881, N879, N877, N875, N873, N871, N869, N867, N865, N863, N861, N859, N857, N855, N853, N851, N849, N847, N845, N843, N841 } : 
                        (N63)? fsgnj_a : 1'b0;
  assign N10 = N48;
  assign N11 = N54;
  assign N12 = N60;
  assign { N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977 } = (N13)? frs2_raw : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N976)? frs1_raw : 1'b0;
  assign N13 = N975;
  assign fminmax_result = (N14)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                          (N1053)? frs2_raw : 
                          (N1056)? frs1_raw : 
                          (N1059)? { N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977 } : 
                          (N1062)? frs1_raw : 
                          (N974)? frs2_raw : 1'b0;
  assign N14 = N966;
  assign ieee_result = (N15)? imvf_result : 
                       (N16)? fsgnj_result : 1'b0;
  assign N15 = N1068;
  assign N16 = N1067;
  assign { N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080 } = (N17)? { i2f_result_is_nan_, i2f_result_is_inf_, i2f_result_is_zero_, 1'b0, 1'b0, i2f_result_sign_, i2f_result_sexp__12_, i2f_result_sexp__11_, i2f_result_sexp__10_, i2f_result_sexp__9_, i2f_result_sexp__8_, i2f_result_sexp__7_, i2f_result_sexp__6_, i2f_result_sexp__5_, i2f_result_sexp__4_, i2f_result_sexp__3_, i2f_result_sexp__2_, i2f_result_sexp__1_, i2f_result_sexp__0_, i2f_sig, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           (N18)? frs1_raw : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           (N19)? fminmax_result : 1'b0;
  assign N17 = N1077;
  assign N18 = N1078;
  assign N19 = N1079;
  assign { N1159, N1158, N1157, N1156, N1155 } = (N17)? { i2f_fflags_nv_, i2f_fflags_dz_, i2f_fflags_of_, i2f_fflags_uf_, i2f_fflags_nx_ } : 
                                                 (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                 (N19)? { fcmp_fflags_nv_, fcmp_fflags_dz_, fcmp_fflags_of_, fcmp_fflags_uf_, fcmp_fflags_nx_ } : 1'b0;
  assign raw_result = (N20)? { N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080 } : 
                      (N1074)? fminmax_result : 1'b0;
  assign N20 = N1073;
  assign { raw_fflags_nv_, raw_fflags_dz_, raw_fflags_of_, raw_fflags_uf_, raw_fflags_nx_ } = (N20)? { N1159, N1158, N1157, N1156, N1155 } : 
                                                                                              (N1074)? { fcmp_fflags_nv_, fcmp_fflags_dz_, fcmp_fflags_of_, fcmp_fflags_uf_, fcmp_fflags_nx_ } : 1'b0;
  assign frd_data_lo = (N21)? ieee_data_lo : 
                       (N1160)? rebox_data_lo : 1'b0;
  assign N21 = reservation_i[420];
  assign { frd_fflags_nv_, frd_fflags_dz_, frd_fflags_of_, frd_fflags_uf_, frd_fflags_nx_ } = (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                              (N1160)? { N1161, N1162, N1163, N1164, N1165 } : 1'b0;
  assign { N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201 } = (N22)? reservation_i[193:130] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N23)? f2i_result : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fcmp_out } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fclass_result_q_nan_, fclass_result_s_nan_, fclass_result_p_inf_, fclass_result_p_norm_, fclass_result_p_sub_, fclass_result_p_zero_, fclass_result_n_zero_, fclass_result_n_sub_, fclass_result_n_norm_, fclass_result_n_inf_ } : 1'b0;
  assign N22 = N1171;
  assign N23 = N1178;
  assign N24 = N1188;
  assign N25 = N1200;
  assign { N1269, N1268, N1267, N1266, N1265 } = (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                 (N23)? { f2i_fflags_nv_, 1'b0, 1'b0, 1'b0, f2i_fflags_nx_ } : 
                                                 (N24)? { fcmp_fflags_nv_, fcmp_fflags_dz_, fcmp_fflags_of_, fcmp_fflags_uf_, fcmp_fflags_nx_ } : 
                                                 (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign iaux_result = (N26)? { N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201 } : 
                       (N1167)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fclass_result_q_nan_, fclass_result_s_nan_, fclass_result_p_inf_, fclass_result_p_norm_, fclass_result_p_sub_, fclass_result_p_zero_, fclass_result_n_zero_, fclass_result_n_sub_, fclass_result_n_norm_, fclass_result_n_inf_ } : 1'b0;
  assign N26 = N1166;
  assign { ird_fflags_nv_, ird_fflags_dz_, ird_fflags_of_, ird_fflags_uf_, ird_fflags_nx_ } = (N26)? { N1269, N1268, N1267, N1266, N1265 } : 
                                                                                              (N1167)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign aux_result = (N27)? ird_data_lo : 
                      (N1270)? frd_data_lo : 1'b0;
  assign N27 = reservation_i[435];
  assign aux_fflags = (N27)? { ird_fflags_nv_, ird_fflags_dz_, ird_fflags_of_, ird_fflags_uf_, ird_fflags_nx_ } : 
                      (N1270)? { frd_fflags_nv_, frd_fflags_dz_, frd_fflags_of_, frd_fflags_uf_, frd_fflags_nx_ } : 1'b0;
  assign N28 = ~N1272;
  assign fclass_result_q_nan_ = frs1_raw[74] & N1309;
  assign N1309 = ~frs1_raw[71];
  assign fclass_result_s_nan_ = frs1_raw[74] & frs1_raw[71];
  assign fclass_result_p_inf_ = N1310 & frs1_raw[73];
  assign N1310 = ~frs1_raw[69];
  assign fclass_result_p_norm_ = N1316 & N1317;
  assign N1316 = N1314 & N1315;
  assign N1314 = N1312 & N1313;
  assign N1312 = N1310 & N1311;
  assign N1311 = ~frs1_raw[70];
  assign N1313 = ~frs1_raw[72];
  assign N1315 = ~frs1_raw[73];
  assign N1317 = ~frs1_raw[74];
  assign fclass_result_p_sub_ = N1310 & frs1_raw[70];
  assign fclass_result_p_zero_ = N1310 & frs1_raw[72];
  assign fclass_result_n_zero_ = frs1_raw[69] & frs1_raw[72];
  assign fclass_result_n_sub_ = frs1_raw[69] & frs1_raw[70];
  assign fclass_result_n_norm_ = N1320 & N1317;
  assign N1320 = N1319 & N1315;
  assign N1319 = N1318 & N1313;
  assign N1318 = frs1_raw[69] & N1311;
  assign fclass_result_n_inf_ = frs1_raw[69] & frs1_raw[73];
  assign _2_net_ = ~irs1_unsigned;
  assign dword_fflags_nv_ = f2dw_iflags_nv_ | f2dw_iflags_of_;
  assign word_fflags_nv_ = f2w_iflags_nv_ | f2w_iflags_of_;
  assign imvf_result[63] = reservation_i[388] | N1295;
  assign imvf_result[62] = reservation_i[387] | N1295;
  assign imvf_result[61] = reservation_i[386] | N1295;
  assign imvf_result[60] = reservation_i[385] | N1295;
  assign imvf_result[59] = reservation_i[384] | N1295;
  assign imvf_result[58] = reservation_i[383] | N1295;
  assign imvf_result[57] = reservation_i[382] | N1295;
  assign imvf_result[56] = reservation_i[381] | N1295;
  assign imvf_result[55] = reservation_i[380] | N1295;
  assign imvf_result[54] = reservation_i[379] | N1295;
  assign imvf_result[53] = reservation_i[378] | N1295;
  assign imvf_result[52] = reservation_i[377] | N1295;
  assign imvf_result[51] = reservation_i[376] | N1295;
  assign imvf_result[50] = reservation_i[375] | N1295;
  assign imvf_result[49] = reservation_i[374] | N1295;
  assign imvf_result[48] = reservation_i[373] | N1295;
  assign imvf_result[47] = reservation_i[372] | N1295;
  assign imvf_result[46] = reservation_i[371] | N1295;
  assign imvf_result[45] = reservation_i[370] | N1295;
  assign imvf_result[44] = reservation_i[369] | N1295;
  assign imvf_result[43] = reservation_i[368] | N1295;
  assign imvf_result[42] = reservation_i[367] | N1295;
  assign imvf_result[41] = reservation_i[366] | N1295;
  assign imvf_result[40] = reservation_i[365] | N1295;
  assign imvf_result[39] = reservation_i[364] | N1295;
  assign imvf_result[38] = reservation_i[363] | N1295;
  assign imvf_result[37] = reservation_i[362] | N1295;
  assign imvf_result[36] = reservation_i[361] | N1295;
  assign imvf_result[35] = reservation_i[360] | N1295;
  assign imvf_result[34] = reservation_i[359] | N1295;
  assign imvf_result[33] = reservation_i[358] | N1295;
  assign imvf_result[32] = reservation_i[357] | N1295;
  assign imvf_result[31] = reservation_i[356] | 1'b0;
  assign imvf_result[30] = reservation_i[355] | 1'b0;
  assign imvf_result[29] = reservation_i[354] | 1'b0;
  assign imvf_result[28] = reservation_i[353] | 1'b0;
  assign imvf_result[27] = reservation_i[352] | 1'b0;
  assign imvf_result[26] = reservation_i[351] | 1'b0;
  assign imvf_result[25] = reservation_i[350] | 1'b0;
  assign imvf_result[24] = reservation_i[349] | 1'b0;
  assign imvf_result[23] = reservation_i[348] | 1'b0;
  assign imvf_result[22] = reservation_i[347] | 1'b0;
  assign imvf_result[21] = reservation_i[346] | 1'b0;
  assign imvf_result[20] = reservation_i[345] | 1'b0;
  assign imvf_result[19] = reservation_i[344] | 1'b0;
  assign imvf_result[18] = reservation_i[343] | 1'b0;
  assign imvf_result[17] = reservation_i[342] | 1'b0;
  assign imvf_result[16] = reservation_i[341] | 1'b0;
  assign imvf_result[15] = reservation_i[340] | 1'b0;
  assign imvf_result[14] = reservation_i[339] | 1'b0;
  assign imvf_result[13] = reservation_i[338] | 1'b0;
  assign imvf_result[12] = reservation_i[337] | 1'b0;
  assign imvf_result[11] = reservation_i[336] | 1'b0;
  assign imvf_result[10] = reservation_i[335] | 1'b0;
  assign imvf_result[9] = reservation_i[334] | 1'b0;
  assign imvf_result[8] = reservation_i[333] | 1'b0;
  assign imvf_result[7] = reservation_i[332] | 1'b0;
  assign imvf_result[6] = reservation_i[331] | 1'b0;
  assign imvf_result[5] = reservation_i[330] | 1'b0;
  assign imvf_result[4] = reservation_i[329] | 1'b0;
  assign imvf_result[3] = reservation_i[328] | 1'b0;
  assign imvf_result[2] = reservation_i[327] | 1'b0;
  assign imvf_result[1] = reservation_i[326] | 1'b0;
  assign imvf_result[0] = reservation_i[325] | 1'b0;
  assign invbox_frs1 = reservation_i[403] & N1352;
  assign N1352 = ~N1351;
  assign N1351 = N1350 & reservation_i[162];
  assign N1350 = N1349 & reservation_i[163];
  assign N1349 = N1348 & reservation_i[164];
  assign N1348 = N1347 & reservation_i[165];
  assign N1347 = N1346 & reservation_i[166];
  assign N1346 = N1345 & reservation_i[167];
  assign N1345 = N1344 & reservation_i[168];
  assign N1344 = N1343 & reservation_i[169];
  assign N1343 = N1342 & reservation_i[170];
  assign N1342 = N1341 & reservation_i[171];
  assign N1341 = N1340 & reservation_i[172];
  assign N1340 = N1339 & reservation_i[173];
  assign N1339 = N1338 & reservation_i[174];
  assign N1338 = N1337 & reservation_i[175];
  assign N1337 = N1336 & reservation_i[176];
  assign N1336 = N1335 & reservation_i[177];
  assign N1335 = N1334 & reservation_i[178];
  assign N1334 = N1333 & reservation_i[179];
  assign N1333 = N1332 & reservation_i[180];
  assign N1332 = N1331 & reservation_i[181];
  assign N1331 = N1330 & reservation_i[182];
  assign N1330 = N1329 & reservation_i[183];
  assign N1329 = N1328 & reservation_i[184];
  assign N1328 = N1327 & reservation_i[185];
  assign N1327 = N1326 & reservation_i[186];
  assign N1326 = N1325 & reservation_i[187];
  assign N1325 = N1324 & reservation_i[188];
  assign N1324 = N1323 & reservation_i[189];
  assign N1323 = N1322 & reservation_i[190];
  assign N1322 = N1321 & reservation_i[191];
  assign N1321 = reservation_i[193] & reservation_i[192];
  assign invbox_frs2 = reservation_i[403] & N1384;
  assign N1384 = ~N1383;
  assign N1383 = N1382 & reservation_i[97];
  assign N1382 = N1381 & reservation_i[98];
  assign N1381 = N1380 & reservation_i[99];
  assign N1380 = N1379 & reservation_i[100];
  assign N1379 = N1378 & reservation_i[101];
  assign N1378 = N1377 & reservation_i[102];
  assign N1377 = N1376 & reservation_i[103];
  assign N1376 = N1375 & reservation_i[104];
  assign N1375 = N1374 & reservation_i[105];
  assign N1374 = N1373 & reservation_i[106];
  assign N1373 = N1372 & reservation_i[107];
  assign N1372 = N1371 & reservation_i[108];
  assign N1371 = N1370 & reservation_i[109];
  assign N1370 = N1369 & reservation_i[110];
  assign N1369 = N1368 & reservation_i[111];
  assign N1368 = N1367 & reservation_i[112];
  assign N1367 = N1366 & reservation_i[113];
  assign N1366 = N1365 & reservation_i[114];
  assign N1365 = N1364 & reservation_i[115];
  assign N1364 = N1363 & reservation_i[116];
  assign N1363 = N1362 & reservation_i[117];
  assign N1362 = N1361 & reservation_i[118];
  assign N1361 = N1360 & reservation_i[119];
  assign N1360 = N1359 & reservation_i[120];
  assign N1359 = N1358 & reservation_i[121];
  assign N1358 = N1357 & reservation_i[122];
  assign N1357 = N1356 & reservation_i[123];
  assign N1356 = N1355 & reservation_i[124];
  assign N1355 = N1354 & reservation_i[125];
  assign N1354 = N1353 & reservation_i[126];
  assign N1353 = reservation_i[128] & reservation_i[127];
  assign N41 = ~invbox_frs1;
  assign N42 = ~invbox_frs2;
  assign N48 = ~N47;
  assign N54 = ~N53;
  assign N60 = ~N59;
  assign N61 = N54 | N48;
  assign N62 = N60 | N61;
  assign N63 = ~N62;
  assign N64 = ~1'b1;
  assign N65 = ~1'b1;
  assign N66 = N64 & N65;
  assign N67 = N64 & 1'b1;
  assign N68 = 1'b1 & N65;
  assign N69 = 1'b1 & 1'b1;
  assign N70 = ~1'b1;
  assign N71 = N66 & N70;
  assign N72 = N66 & 1'b1;
  assign N73 = N68 & N70;
  assign N74 = N68 & 1'b1;
  assign N75 = N67 & N70;
  assign N76 = N67 & 1'b1;
  assign N77 = N69 & N70;
  assign N78 = N69 & 1'b1;
  assign N79 = ~1'b1;
  assign N80 = N71 & N79;
  assign N81 = N71 & 1'b1;
  assign N82 = N73 & N79;
  assign N83 = N73 & 1'b1;
  assign N84 = N75 & N79;
  assign N85 = N75 & 1'b1;
  assign N86 = N77 & N79;
  assign N87 = N77 & 1'b1;
  assign N88 = N72 & N79;
  assign N89 = N72 & 1'b1;
  assign N90 = N74 & N79;
  assign N91 = N74 & 1'b1;
  assign N92 = N76 & N79;
  assign N93 = N76 & 1'b1;
  assign N94 = N78 & N79;
  assign N95 = N78 & 1'b1;
  assign N96 = ~1'b1;
  assign N97 = N80 & N96;
  assign N98 = N80 & 1'b1;
  assign N99 = N82 & N96;
  assign N100 = N82 & 1'b1;
  assign N101 = N84 & N96;
  assign N102 = N84 & 1'b1;
  assign N103 = N86 & N96;
  assign N104 = N86 & 1'b1;
  assign N105 = N88 & N96;
  assign N106 = N88 & 1'b1;
  assign N107 = N90 & N96;
  assign N108 = N90 & 1'b1;
  assign N109 = N92 & N96;
  assign N110 = N92 & 1'b1;
  assign N111 = N94 & N96;
  assign N112 = N94 & 1'b1;
  assign N113 = N81 & N96;
  assign N114 = N81 & 1'b1;
  assign N115 = N83 & N96;
  assign N116 = N83 & 1'b1;
  assign N117 = N85 & N96;
  assign N118 = N85 & 1'b1;
  assign N119 = N87 & N96;
  assign N120 = N87 & 1'b1;
  assign N121 = N89 & N96;
  assign N122 = N89 & 1'b1;
  assign N123 = N91 & N96;
  assign N124 = N91 & 1'b1;
  assign N125 = N93 & N96;
  assign N126 = N93 & 1'b1;
  assign N127 = N95 & N96;
  assign N128 = N95 & 1'b1;
  assign N129 = ~N1308;
  assign N130 = N97 & N129;
  assign N131 = N97 & N1308;
  assign N132 = N99 & N129;
  assign N133 = N99 & N1308;
  assign N134 = N101 & N129;
  assign N135 = N101 & N1308;
  assign N136 = N103 & N129;
  assign N137 = N103 & N1308;
  assign N138 = N105 & N129;
  assign N139 = N105 & N1308;
  assign N140 = N107 & N129;
  assign N141 = N107 & N1308;
  assign N142 = N109 & N129;
  assign N143 = N109 & N1308;
  assign N144 = N111 & N129;
  assign N145 = N111 & N1308;
  assign N146 = N113 & N129;
  assign N147 = N113 & N1308;
  assign N148 = N115 & N129;
  assign N149 = N115 & N1308;
  assign N150 = N117 & N129;
  assign N151 = N117 & N1308;
  assign N152 = N119 & N129;
  assign N153 = N119 & N1308;
  assign N154 = N121 & N129;
  assign N155 = N121 & N1308;
  assign N156 = N123 & N129;
  assign N157 = N123 & N1308;
  assign N158 = N125 & N129;
  assign N159 = N125 & N1308;
  assign N160 = N127 & N129;
  assign N161 = N127 & N1308;
  assign N162 = N98 & N129;
  assign N163 = N98 & N1308;
  assign N164 = N100 & N129;
  assign N165 = N100 & N1308;
  assign N166 = N102 & N129;
  assign N167 = N102 & N1308;
  assign N168 = N104 & N129;
  assign N169 = N104 & N1308;
  assign N170 = N106 & N129;
  assign N171 = N106 & N1308;
  assign N172 = N108 & N129;
  assign N173 = N108 & N1308;
  assign N174 = N110 & N129;
  assign N175 = N110 & N1308;
  assign N176 = N112 & N129;
  assign N177 = N112 & N1308;
  assign N178 = N114 & N129;
  assign N179 = N114 & N1308;
  assign N180 = N116 & N129;
  assign N181 = N116 & N1308;
  assign N182 = N118 & N129;
  assign N183 = N118 & N1308;
  assign N184 = N120 & N129;
  assign N185 = N120 & N1308;
  assign N186 = N122 & N129;
  assign N187 = N122 & N1308;
  assign N188 = N124 & N129;
  assign N189 = N124 & N1308;
  assign N190 = N126 & N129;
  assign N191 = N126 & N1308;
  assign N192 = N128 & N129;
  assign N193 = N128 & N1308;
  assign N196 = ~N194;
  assign N197 = ~1'b0;
  assign N199 = ~1'b0;
  assign N201 = ~1'b0;
  assign N203 = ~1'b0;
  assign N205 = ~1'b0;
  assign N207 = ~1'b0;
  assign N209 = ~1'b0;
  assign N211 = ~1'b0;
  assign N213 = ~1'b0;
  assign N215 = ~1'b0;
  assign N217 = ~1'b0;
  assign N219 = ~1'b0;
  assign N221 = ~1'b0;
  assign N223 = ~1'b0;
  assign N225 = ~1'b0;
  assign N227 = ~1'b0;
  assign N229 = ~1'b0;
  assign N231 = ~1'b0;
  assign N233 = ~1'b0;
  assign N235 = ~1'b0;
  assign N237 = ~1'b0;
  assign N239 = ~1'b0;
  assign N241 = ~1'b0;
  assign N243 = ~1'b0;
  assign N245 = ~1'b0;
  assign N247 = ~1'b0;
  assign N249 = ~1'b0;
  assign N251 = ~1'b0;
  assign N253 = ~1'b0;
  assign N255 = ~1'b0;
  assign N257 = ~1'b0;
  assign N260 = ~1'b0;
  assign N262 = ~1'b0;
  assign N264 = ~1'b0;
  assign N266 = ~1'b0;
  assign N268 = ~1'b0;
  assign N270 = ~1'b0;
  assign N272 = ~1'b0;
  assign N274 = ~1'b0;
  assign N276 = ~1'b0;
  assign N278 = ~1'b0;
  assign N280 = ~1'b0;
  assign N282 = ~1'b0;
  assign N284 = ~1'b0;
  assign N286 = ~1'b0;
  assign N288 = ~1'b0;
  assign N290 = ~1'b0;
  assign N292 = ~1'b0;
  assign N294 = ~1'b0;
  assign N296 = ~1'b0;
  assign N298 = ~1'b0;
  assign N300 = ~1'b0;
  assign N302 = ~1'b0;
  assign N304 = ~1'b0;
  assign N306 = ~1'b0;
  assign N308 = ~1'b0;
  assign N310 = ~1'b0;
  assign N312 = ~1'b0;
  assign N314 = ~1'b0;
  assign N316 = ~1'b0;
  assign N318 = ~1'b0;
  assign N320 = ~1'b0;
  assign N323 = ~1'b1;
  assign N324 = ~1'b1;
  assign N325 = N323 & N324;
  assign N326 = N323 & 1'b1;
  assign N327 = 1'b1 & N324;
  assign N328 = 1'b1 & 1'b1;
  assign N329 = ~1'b1;
  assign N330 = N325 & N329;
  assign N331 = N325 & 1'b1;
  assign N332 = N327 & N329;
  assign N333 = N327 & 1'b1;
  assign N334 = N326 & N329;
  assign N335 = N326 & 1'b1;
  assign N336 = N328 & N329;
  assign N337 = N328 & 1'b1;
  assign N338 = ~1'b1;
  assign N339 = N330 & N338;
  assign N340 = N330 & 1'b1;
  assign N341 = N332 & N338;
  assign N342 = N332 & 1'b1;
  assign N343 = N334 & N338;
  assign N344 = N334 & 1'b1;
  assign N345 = N336 & N338;
  assign N346 = N336 & 1'b1;
  assign N347 = N331 & N338;
  assign N348 = N331 & 1'b1;
  assign N349 = N333 & N338;
  assign N350 = N333 & 1'b1;
  assign N351 = N335 & N338;
  assign N352 = N335 & 1'b1;
  assign N353 = N337 & N338;
  assign N354 = N337 & 1'b1;
  assign N355 = ~1'b1;
  assign N356 = N339 & N355;
  assign N357 = N339 & 1'b1;
  assign N358 = N341 & N355;
  assign N359 = N341 & 1'b1;
  assign N360 = N343 & N355;
  assign N361 = N343 & 1'b1;
  assign N362 = N345 & N355;
  assign N363 = N345 & 1'b1;
  assign N364 = N347 & N355;
  assign N365 = N347 & 1'b1;
  assign N366 = N349 & N355;
  assign N367 = N349 & 1'b1;
  assign N368 = N351 & N355;
  assign N369 = N351 & 1'b1;
  assign N370 = N353 & N355;
  assign N371 = N353 & 1'b1;
  assign N372 = N340 & N355;
  assign N373 = N340 & 1'b1;
  assign N374 = N342 & N355;
  assign N375 = N342 & 1'b1;
  assign N376 = N344 & N355;
  assign N377 = N344 & 1'b1;
  assign N378 = N346 & N355;
  assign N379 = N346 & 1'b1;
  assign N380 = N348 & N355;
  assign N381 = N348 & 1'b1;
  assign N382 = N350 & N355;
  assign N383 = N350 & 1'b1;
  assign N384 = N352 & N355;
  assign N385 = N352 & 1'b1;
  assign N386 = N354 & N355;
  assign N387 = N354 & 1'b1;
  assign N388 = N356 & N129;
  assign N389 = N356 & N1308;
  assign N390 = N358 & N129;
  assign N391 = N358 & N1308;
  assign N392 = N360 & N129;
  assign N393 = N360 & N1308;
  assign N394 = N362 & N129;
  assign N395 = N362 & N1308;
  assign N396 = N364 & N129;
  assign N397 = N364 & N1308;
  assign N398 = N366 & N129;
  assign N399 = N366 & N1308;
  assign N400 = N368 & N129;
  assign N401 = N368 & N1308;
  assign N402 = N370 & N129;
  assign N403 = N370 & N1308;
  assign N404 = N372 & N129;
  assign N405 = N372 & N1308;
  assign N406 = N374 & N129;
  assign N407 = N374 & N1308;
  assign N408 = N376 & N129;
  assign N409 = N376 & N1308;
  assign N410 = N378 & N129;
  assign N411 = N378 & N1308;
  assign N412 = N380 & N129;
  assign N413 = N380 & N1308;
  assign N414 = N382 & N129;
  assign N415 = N382 & N1308;
  assign N416 = N384 & N129;
  assign N417 = N384 & N1308;
  assign N418 = N386 & N129;
  assign N419 = N386 & N1308;
  assign N420 = N357 & N129;
  assign N421 = N357 & N1308;
  assign N422 = N359 & N129;
  assign N423 = N359 & N1308;
  assign N424 = N361 & N129;
  assign N425 = N361 & N1308;
  assign N426 = N363 & N129;
  assign N427 = N363 & N1308;
  assign N428 = N365 & N129;
  assign N429 = N365 & N1308;
  assign N430 = N367 & N129;
  assign N431 = N367 & N1308;
  assign N432 = N369 & N129;
  assign N433 = N369 & N1308;
  assign N434 = N371 & N129;
  assign N435 = N371 & N1308;
  assign N436 = N373 & N129;
  assign N437 = N373 & N1308;
  assign N438 = N375 & N129;
  assign N439 = N375 & N1308;
  assign N440 = N377 & N129;
  assign N441 = N377 & N1308;
  assign N442 = N379 & N129;
  assign N443 = N379 & N1308;
  assign N444 = N381 & N129;
  assign N445 = N381 & N1308;
  assign N446 = N383 & N129;
  assign N447 = N383 & N1308;
  assign N448 = N385 & N129;
  assign N449 = N385 & N1308;
  assign N450 = N387 & N129;
  assign N451 = N387 & N1308;
  assign N453 = ~1'b1;
  assign N454 = ~1'b1;
  assign N455 = N453 & N454;
  assign N456 = N453 & 1'b1;
  assign N457 = 1'b1 & N454;
  assign N458 = 1'b1 & 1'b1;
  assign N459 = ~1'b1;
  assign N460 = N455 & N459;
  assign N461 = N455 & 1'b1;
  assign N462 = N457 & N459;
  assign N463 = N457 & 1'b1;
  assign N464 = N456 & N459;
  assign N465 = N456 & 1'b1;
  assign N466 = N458 & N459;
  assign N467 = N458 & 1'b1;
  assign N468 = ~1'b1;
  assign N469 = N460 & N468;
  assign N470 = N460 & 1'b1;
  assign N471 = N462 & N468;
  assign N472 = N462 & 1'b1;
  assign N473 = N464 & N468;
  assign N474 = N464 & 1'b1;
  assign N475 = N466 & N468;
  assign N476 = N466 & 1'b1;
  assign N477 = N461 & N468;
  assign N478 = N461 & 1'b1;
  assign N479 = N463 & N468;
  assign N480 = N463 & 1'b1;
  assign N481 = N465 & N468;
  assign N482 = N465 & 1'b1;
  assign N483 = N467 & N468;
  assign N484 = N467 & 1'b1;
  assign N485 = ~1'b1;
  assign N486 = N469 & N485;
  assign N487 = N469 & 1'b1;
  assign N488 = N471 & N485;
  assign N489 = N471 & 1'b1;
  assign N490 = N473 & N485;
  assign N491 = N473 & 1'b1;
  assign N492 = N475 & N485;
  assign N493 = N475 & 1'b1;
  assign N494 = N477 & N485;
  assign N495 = N477 & 1'b1;
  assign N496 = N479 & N485;
  assign N497 = N479 & 1'b1;
  assign N498 = N481 & N485;
  assign N499 = N481 & 1'b1;
  assign N500 = N483 & N485;
  assign N501 = N483 & 1'b1;
  assign N502 = N470 & N485;
  assign N503 = N470 & 1'b1;
  assign N504 = N472 & N485;
  assign N505 = N472 & 1'b1;
  assign N506 = N474 & N485;
  assign N507 = N474 & 1'b1;
  assign N508 = N476 & N485;
  assign N509 = N476 & 1'b1;
  assign N510 = N478 & N485;
  assign N511 = N478 & 1'b1;
  assign N512 = N480 & N485;
  assign N513 = N480 & 1'b1;
  assign N514 = N482 & N485;
  assign N515 = N482 & 1'b1;
  assign N516 = N484 & N485;
  assign N517 = N484 & 1'b1;
  assign N518 = N486 & N129;
  assign N519 = N486 & N1308;
  assign N520 = N488 & N129;
  assign N521 = N488 & N1308;
  assign N522 = N490 & N129;
  assign N523 = N490 & N1308;
  assign N524 = N492 & N129;
  assign N525 = N492 & N1308;
  assign N526 = N494 & N129;
  assign N527 = N494 & N1308;
  assign N528 = N496 & N129;
  assign N529 = N496 & N1308;
  assign N530 = N498 & N129;
  assign N531 = N498 & N1308;
  assign N532 = N500 & N129;
  assign N533 = N500 & N1308;
  assign N534 = N502 & N129;
  assign N535 = N502 & N1308;
  assign N536 = N504 & N129;
  assign N537 = N504 & N1308;
  assign N538 = N506 & N129;
  assign N539 = N506 & N1308;
  assign N540 = N508 & N129;
  assign N541 = N508 & N1308;
  assign N542 = N510 & N129;
  assign N543 = N510 & N1308;
  assign N544 = N512 & N129;
  assign N545 = N512 & N1308;
  assign N546 = N514 & N129;
  assign N547 = N514 & N1308;
  assign N548 = N516 & N129;
  assign N549 = N516 & N1308;
  assign N550 = N487 & N129;
  assign N551 = N487 & N1308;
  assign N552 = N489 & N129;
  assign N553 = N489 & N1308;
  assign N554 = N491 & N129;
  assign N555 = N491 & N1308;
  assign N556 = N493 & N129;
  assign N557 = N493 & N1308;
  assign N558 = N495 & N129;
  assign N559 = N495 & N1308;
  assign N560 = N497 & N129;
  assign N561 = N497 & N1308;
  assign N562 = N499 & N129;
  assign N563 = N499 & N1308;
  assign N564 = N501 & N129;
  assign N565 = N501 & N1308;
  assign N566 = N503 & N129;
  assign N567 = N503 & N1308;
  assign N568 = N505 & N129;
  assign N569 = N505 & N1308;
  assign N570 = N507 & N129;
  assign N571 = N507 & N1308;
  assign N572 = N509 & N129;
  assign N573 = N509 & N1308;
  assign N574 = N511 & N129;
  assign N575 = N511 & N1308;
  assign N576 = N513 & N129;
  assign N577 = N513 & N1308;
  assign N578 = N515 & N129;
  assign N579 = N515 & N1308;
  assign N580 = N517 & N129;
  assign N581 = N517 & N1308;
  assign N583 = N452 ^ N582;
  assign N584 = ~1'b0;
  assign N586 = ~1'b0;
  assign N588 = ~1'b0;
  assign N590 = ~1'b0;
  assign N592 = ~1'b0;
  assign N594 = ~1'b0;
  assign N596 = ~1'b0;
  assign N598 = ~1'b0;
  assign N600 = ~1'b0;
  assign N602 = ~1'b0;
  assign N604 = ~1'b0;
  assign N606 = ~1'b0;
  assign N608 = ~1'b0;
  assign N610 = ~1'b0;
  assign N612 = ~1'b0;
  assign N614 = ~1'b0;
  assign N616 = ~1'b0;
  assign N618 = ~1'b0;
  assign N620 = ~1'b0;
  assign N622 = ~1'b0;
  assign N624 = ~1'b0;
  assign N626 = ~1'b0;
  assign N628 = ~1'b0;
  assign N630 = ~1'b0;
  assign N632 = ~1'b0;
  assign N634 = ~1'b0;
  assign N636 = ~1'b0;
  assign N638 = ~1'b0;
  assign N640 = ~1'b0;
  assign N642 = ~1'b0;
  assign N644 = ~1'b0;
  assign N647 = ~1'b0;
  assign N649 = ~1'b0;
  assign N651 = ~1'b0;
  assign N653 = ~1'b0;
  assign N655 = ~1'b0;
  assign N657 = ~1'b0;
  assign N659 = ~1'b0;
  assign N661 = ~1'b0;
  assign N663 = ~1'b0;
  assign N665 = ~1'b0;
  assign N667 = ~1'b0;
  assign N669 = ~1'b0;
  assign N671 = ~1'b0;
  assign N673 = ~1'b0;
  assign N675 = ~1'b0;
  assign N677 = ~1'b0;
  assign N679 = ~1'b0;
  assign N681 = ~1'b0;
  assign N683 = ~1'b0;
  assign N685 = ~1'b0;
  assign N687 = ~1'b0;
  assign N689 = ~1'b0;
  assign N691 = ~1'b0;
  assign N693 = ~1'b0;
  assign N695 = ~1'b0;
  assign N697 = ~1'b0;
  assign N699 = ~1'b0;
  assign N701 = ~1'b0;
  assign N703 = ~1'b0;
  assign N705 = ~1'b0;
  assign N707 = ~1'b0;
  assign N710 = ~1'b1;
  assign N711 = ~1'b1;
  assign N712 = N710 & N711;
  assign N713 = N710 & 1'b1;
  assign N714 = 1'b1 & N711;
  assign N715 = 1'b1 & 1'b1;
  assign N716 = ~1'b1;
  assign N717 = N712 & N716;
  assign N718 = N712 & 1'b1;
  assign N719 = N714 & N716;
  assign N720 = N714 & 1'b1;
  assign N721 = N713 & N716;
  assign N722 = N713 & 1'b1;
  assign N723 = N715 & N716;
  assign N724 = N715 & 1'b1;
  assign N725 = ~1'b1;
  assign N726 = N717 & N725;
  assign N727 = N717 & 1'b1;
  assign N728 = N719 & N725;
  assign N729 = N719 & 1'b1;
  assign N730 = N721 & N725;
  assign N731 = N721 & 1'b1;
  assign N732 = N723 & N725;
  assign N733 = N723 & 1'b1;
  assign N734 = N718 & N725;
  assign N735 = N718 & 1'b1;
  assign N736 = N720 & N725;
  assign N737 = N720 & 1'b1;
  assign N738 = N722 & N725;
  assign N739 = N722 & 1'b1;
  assign N740 = N724 & N725;
  assign N741 = N724 & 1'b1;
  assign N742 = ~1'b1;
  assign N743 = N726 & N742;
  assign N744 = N726 & 1'b1;
  assign N745 = N728 & N742;
  assign N746 = N728 & 1'b1;
  assign N747 = N730 & N742;
  assign N748 = N730 & 1'b1;
  assign N749 = N732 & N742;
  assign N750 = N732 & 1'b1;
  assign N751 = N734 & N742;
  assign N752 = N734 & 1'b1;
  assign N753 = N736 & N742;
  assign N754 = N736 & 1'b1;
  assign N755 = N738 & N742;
  assign N756 = N738 & 1'b1;
  assign N757 = N740 & N742;
  assign N758 = N740 & 1'b1;
  assign N759 = N727 & N742;
  assign N760 = N727 & 1'b1;
  assign N761 = N729 & N742;
  assign N762 = N729 & 1'b1;
  assign N763 = N731 & N742;
  assign N764 = N731 & 1'b1;
  assign N765 = N733 & N742;
  assign N766 = N733 & 1'b1;
  assign N767 = N735 & N742;
  assign N768 = N735 & 1'b1;
  assign N769 = N737 & N742;
  assign N770 = N737 & 1'b1;
  assign N771 = N739 & N742;
  assign N772 = N739 & 1'b1;
  assign N773 = N741 & N742;
  assign N774 = N741 & 1'b1;
  assign N775 = N743 & N129;
  assign N776 = N743 & N1308;
  assign N777 = N745 & N129;
  assign N778 = N745 & N1308;
  assign N779 = N747 & N129;
  assign N780 = N747 & N1308;
  assign N781 = N749 & N129;
  assign N782 = N749 & N1308;
  assign N783 = N751 & N129;
  assign N784 = N751 & N1308;
  assign N785 = N753 & N129;
  assign N786 = N753 & N1308;
  assign N787 = N755 & N129;
  assign N788 = N755 & N1308;
  assign N789 = N757 & N129;
  assign N790 = N757 & N1308;
  assign N791 = N759 & N129;
  assign N792 = N759 & N1308;
  assign N793 = N761 & N129;
  assign N794 = N761 & N1308;
  assign N795 = N763 & N129;
  assign N796 = N763 & N1308;
  assign N797 = N765 & N129;
  assign N798 = N765 & N1308;
  assign N799 = N767 & N129;
  assign N800 = N767 & N1308;
  assign N801 = N769 & N129;
  assign N802 = N769 & N1308;
  assign N803 = N771 & N129;
  assign N804 = N771 & N1308;
  assign N805 = N773 & N129;
  assign N806 = N773 & N1308;
  assign N807 = N744 & N129;
  assign N808 = N744 & N1308;
  assign N809 = N746 & N129;
  assign N810 = N746 & N1308;
  assign N811 = N748 & N129;
  assign N812 = N748 & N1308;
  assign N813 = N750 & N129;
  assign N814 = N750 & N1308;
  assign N815 = N752 & N129;
  assign N816 = N752 & N1308;
  assign N817 = N754 & N129;
  assign N818 = N754 & N1308;
  assign N819 = N756 & N129;
  assign N820 = N756 & N1308;
  assign N821 = N758 & N129;
  assign N822 = N758 & N1308;
  assign N823 = N760 & N129;
  assign N824 = N760 & N1308;
  assign N825 = N762 & N129;
  assign N826 = N762 & N1308;
  assign N827 = N764 & N129;
  assign N828 = N764 & N1308;
  assign N829 = N766 & N129;
  assign N830 = N766 & N1308;
  assign N831 = N768 & N129;
  assign N832 = N768 & N1308;
  assign N833 = N770 & N129;
  assign N834 = N770 & N1308;
  assign N835 = N772 & N129;
  assign N836 = N772 & N1308;
  assign N837 = N774 & N129;
  assign N838 = N774 & N1308;
  assign N840 = ~1'b0;
  assign N842 = ~1'b0;
  assign N844 = ~1'b0;
  assign N846 = ~1'b0;
  assign N848 = ~1'b0;
  assign N850 = ~1'b0;
  assign N852 = ~1'b0;
  assign N854 = ~1'b0;
  assign N856 = ~1'b0;
  assign N858 = ~1'b0;
  assign N860 = ~1'b0;
  assign N862 = ~1'b0;
  assign N864 = ~1'b0;
  assign N866 = ~1'b0;
  assign N868 = ~1'b0;
  assign N870 = ~1'b0;
  assign N872 = ~1'b0;
  assign N874 = ~1'b0;
  assign N876 = ~1'b0;
  assign N878 = ~1'b0;
  assign N880 = ~1'b0;
  assign N882 = ~1'b0;
  assign N884 = ~1'b0;
  assign N886 = ~1'b0;
  assign N888 = ~1'b0;
  assign N890 = ~1'b0;
  assign N892 = ~1'b0;
  assign N894 = ~1'b0;
  assign N896 = ~1'b0;
  assign N898 = ~1'b0;
  assign N900 = ~1'b0;
  assign N903 = ~1'b0;
  assign N905 = ~1'b0;
  assign N907 = ~1'b0;
  assign N909 = ~1'b0;
  assign N911 = ~1'b0;
  assign N913 = ~1'b0;
  assign N915 = ~1'b0;
  assign N917 = ~1'b0;
  assign N919 = ~1'b0;
  assign N921 = ~1'b0;
  assign N923 = ~1'b0;
  assign N925 = ~1'b0;
  assign N927 = ~1'b0;
  assign N929 = ~1'b0;
  assign N931 = ~1'b0;
  assign N933 = ~1'b0;
  assign N935 = ~1'b0;
  assign N937 = ~1'b0;
  assign N939 = ~1'b0;
  assign N941 = ~1'b0;
  assign N943 = ~1'b0;
  assign N945 = ~1'b0;
  assign N947 = ~1'b0;
  assign N949 = ~1'b0;
  assign N951 = ~1'b0;
  assign N953 = ~1'b0;
  assign N955 = ~1'b0;
  assign N957 = ~1'b0;
  assign N959 = ~1'b0;
  assign N961 = ~1'b0;
  assign N963 = ~1'b0;
  assign signaling_li = N1286 | N1292;
  assign fcmp_out = N1387 | N1389;
  assign N1387 = N1385 | N1386;
  assign N1385 = N1280 & feq_lo;
  assign N1386 = N1286 & flt_lo;
  assign N1389 = N1292 & N1388;
  assign N1388 = flt_lo | feq_lo;
  assign N966 = frs1_raw[74] & frs2_raw[74];
  assign N967 = frs1_raw[74] & N1390;
  assign N1390 = ~frs2_raw[74];
  assign N968 = N1317 & frs2_raw[74];
  assign N969 = N1307 ^ flt_lo;
  assign N970 = N967 | N966;
  assign N971 = N968 | N970;
  assign N972 = feq_lo | N971;
  assign N973 = N969 | N972;
  assign N974 = ~N973;
  assign N975 = N1301 ^ frs1_raw[69];
  assign N976 = ~N975;
  assign N1052 = ~N966;
  assign N1053 = N967 & N1052;
  assign N1054 = ~N967;
  assign N1055 = N1052 & N1054;
  assign N1056 = N968 & N1055;
  assign N1057 = ~N968;
  assign N1058 = N1055 & N1057;
  assign N1059 = feq_lo & N1058;
  assign N1060 = ~feq_lo;
  assign N1061 = N1058 & N1060;
  assign N1062 = N969 & N1061;
  assign N1068 = ~N1067;
  assign N1069 = ~reservation_i[409];
  assign N1070 = ~reservation_i[408];
  assign N1074 = ~N1073;
  assign N1077 = N1391 | N1392;
  assign N1391 = ~N1075;
  assign N1392 = ~N1076;
  assign N1160 = ~reservation_i[420];
  assign N1161 = raw_fflags_nv_ | rebox_fflags_nv_;
  assign N1162 = raw_fflags_dz_ | rebox_fflags_dz_;
  assign N1163 = raw_fflags_of_ | rebox_fflags_of_;
  assign N1164 = raw_fflags_uf_ | rebox_fflags_uf_;
  assign N1165 = raw_fflags_nx_ | rebox_fflags_nx_;
  assign N1167 = ~N1166;
  assign N1171 = ~N1170;
  assign N1178 = N1393 | N1394;
  assign N1393 = ~N1174;
  assign N1394 = ~N1177;
  assign N1188 = N1397 | N1398;
  assign N1397 = N1395 | N1396;
  assign N1395 = ~N1181;
  assign N1396 = ~N1184;
  assign N1398 = ~N1187;
  assign N1200 = N1189 | N1402;
  assign N1402 = N1191 | N1401;
  assign N1401 = N1193 | N1400;
  assign N1400 = N1195 | N1399;
  assign N1399 = N1197 | N1199;
  assign N1270 = ~reservation_i[435];
  assign aux_v_li = reservation_i[520] & reservation_i[446];

endmodule



module bsg_dff_width_p1
(
  clk_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  wire [0:0] data_o;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_chain_width_p1_num_stages_p2
(
  clk_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  wire [0:0] data_o;
  wire \chained.data_delayed_1__0_ ;

  bsg_dff_width_p1
  \chained.genblk1_1_.ch_reg 
  (
    .clk_i(clk_i),
    .data_i(data_i[0]),
    .data_o(\chained.data_delayed_1__0_ )
  );


  bsg_dff_width_p1
  \chained.genblk1_2_.ch_reg 
  (
    .clk_i(clk_i),
    .data_i(\chained.data_delayed_1__0_ ),
    .data_o(data_o[0])
  );


endmodule



module bsg_dff_reset_en_width_p59
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [58:0] data_i;
  output [58:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [58:0] data_o;
  wire N0,N1,N2;
  reg data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,data_o_55_sv2v_reg,
  data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,data_o_51_sv2v_reg,
  data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,data_o_47_sv2v_reg,
  data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,data_o_43_sv2v_reg,
  data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,
  data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,
  data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,
  data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,
  data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,
  data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,
  data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,
  data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,
  data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_58_sv2v_reg <= 1'b0;
      data_o_57_sv2v_reg <= 1'b0;
      data_o_56_sv2v_reg <= 1'b0;
      data_o_55_sv2v_reg <= 1'b0;
      data_o_54_sv2v_reg <= 1'b0;
      data_o_53_sv2v_reg <= 1'b0;
      data_o_52_sv2v_reg <= 1'b0;
      data_o_51_sv2v_reg <= 1'b0;
      data_o_50_sv2v_reg <= 1'b0;
      data_o_49_sv2v_reg <= 1'b0;
      data_o_48_sv2v_reg <= 1'b0;
      data_o_47_sv2v_reg <= 1'b0;
      data_o_46_sv2v_reg <= 1'b0;
      data_o_45_sv2v_reg <= 1'b0;
      data_o_44_sv2v_reg <= 1'b0;
      data_o_43_sv2v_reg <= 1'b0;
      data_o_42_sv2v_reg <= 1'b0;
      data_o_41_sv2v_reg <= 1'b0;
      data_o_40_sv2v_reg <= 1'b0;
      data_o_39_sv2v_reg <= 1'b0;
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_rotate_left_width_p36
(
  data_i,
  rot_i,
  o
);

  input [35:0] data_i;
  input [5:0] rot_i;
  output [35:0] o;
  wire [35:0] o;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,
  sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,
  sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,sv2v_dc_21,sv2v_dc_22,
  sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,sv2v_dc_27,sv2v_dc_28,sv2v_dc_29,
  sv2v_dc_30,sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,sv2v_dc_34,sv2v_dc_35,sv2v_dc_36;
  assign { o, sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36 } = { data_i, data_i } << rot_i;

endmodule



module bsg_dff_en_0000001b
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [26:0] data_i;
  output [26:0] data_o;
  input clk_i;
  input en_i;
  wire [26:0] data_o;
  reg data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,
  data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,
  data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,
  data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_en_width_p1
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [0:0] data_o;
  wire N0,N1,N2;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_cam_1r1w_tag_array_0000001b_00000008
(
  clk_i,
  reset_i,
  w_v_i,
  w_set_not_clear_i,
  w_tag_i,
  w_empty_o,
  r_v_i,
  r_tag_i,
  r_match_o
);

  input [7:0] w_v_i;
  input [26:0] w_tag_i;
  output [7:0] w_empty_o;
  input [26:0] r_tag_i;
  output [7:0] r_match_o;
  input clk_i;
  input reset_i;
  input w_set_not_clear_i;
  input r_v_i;
  wire [7:0] w_empty_o,r_match_o,v_r;
  wire _0_net_,N0,_1_net_,N1,_2_net_,N2,_3_net_,N3,_4_net_,N4,_5_net_,N5,_6_net_,N6,
  _7_net_,N7,N8,N9,N10,N11,N12,N13,N14,N15;
  wire [215:0] tag_r;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_0_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[0]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[0])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_0_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_0_net_),
    .data_o(tag_r[26:0])
  );

  assign N0 = tag_r[26:0] == r_tag_i;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_1_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[1]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[1])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_1_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_1_net_),
    .data_o(tag_r[53:27])
  );

  assign N1 = tag_r[53:27] == r_tag_i;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_2_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[2]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[2])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_2_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_2_net_),
    .data_o(tag_r[80:54])
  );

  assign N2 = tag_r[80:54] == r_tag_i;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_3_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[3]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[3])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_3_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_3_net_),
    .data_o(tag_r[107:81])
  );

  assign N3 = tag_r[107:81] == r_tag_i;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_4_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[4]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[4])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_4_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_4_net_),
    .data_o(tag_r[134:108])
  );

  assign N4 = tag_r[134:108] == r_tag_i;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_5_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[5]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[5])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_5_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_5_net_),
    .data_o(tag_r[161:135])
  );

  assign N5 = tag_r[161:135] == r_tag_i;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_6_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[6]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[6])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_6_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_6_net_),
    .data_o(tag_r[188:162])
  );

  assign N6 = tag_r[188:162] == r_tag_i;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_7_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[7]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[7])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_7_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_7_net_),
    .data_o(tag_r[215:189])
  );

  assign N7 = tag_r[215:189] == r_tag_i;
  assign _0_net_ = w_v_i[0] & w_set_not_clear_i;
  assign r_match_o[0] = N8 & N0;
  assign N8 = r_v_i & v_r[0];
  assign w_empty_o[0] = ~v_r[0];
  assign _1_net_ = w_v_i[1] & w_set_not_clear_i;
  assign r_match_o[1] = N9 & N1;
  assign N9 = r_v_i & v_r[1];
  assign w_empty_o[1] = ~v_r[1];
  assign _2_net_ = w_v_i[2] & w_set_not_clear_i;
  assign r_match_o[2] = N10 & N2;
  assign N10 = r_v_i & v_r[2];
  assign w_empty_o[2] = ~v_r[2];
  assign _3_net_ = w_v_i[3] & w_set_not_clear_i;
  assign r_match_o[3] = N11 & N3;
  assign N11 = r_v_i & v_r[3];
  assign w_empty_o[3] = ~v_r[3];
  assign _4_net_ = w_v_i[4] & w_set_not_clear_i;
  assign r_match_o[4] = N12 & N4;
  assign N12 = r_v_i & v_r[4];
  assign w_empty_o[4] = ~v_r[4];
  assign _5_net_ = w_v_i[5] & w_set_not_clear_i;
  assign r_match_o[5] = N13 & N5;
  assign N13 = r_v_i & v_r[5];
  assign w_empty_o[5] = ~v_r[5];
  assign _6_net_ = w_v_i[6] & w_set_not_clear_i;
  assign r_match_o[6] = N14 & N6;
  assign N14 = r_v_i & v_r[6];
  assign w_empty_o[6] = ~v_r[6];
  assign _7_net_ = w_v_i[7] & w_set_not_clear_i;
  assign r_match_o[7] = N15 & N7;
  assign N15 = r_v_i & v_r[7];
  assign w_empty_o[7] = ~v_r[7];

endmodule



module bsg_dff_reset_en_00000007
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [6:0] data_i;
  output [6:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [6:0] data_o;
  wire N0,N1,N2;
  reg data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mux_width_p1_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [1:0] data_i;
  input [0:0] sel_i;
  output [0:0] data_o;
  wire [0:0] data_o;
  wire N0,N1;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[1] : 1'b0;
  assign N0 = sel_i[0];
  assign N1 = ~sel_i[0];

endmodule



module bsg_mux_width_p1_els_p4
(
  data_i,
  sel_i,
  data_o
);

  input [3:0] data_i;
  input [1:0] sel_i;
  output [0:0] data_o;
  wire [0:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[1] : 
                     (N3)? data_i[2] : 
                     (N5)? data_i[3] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_lru_pseudo_tree_encode_00000008
(
  lru_i,
  way_id_o
);

  input [6:0] lru_i;
  output [2:0] way_id_o;
  wire [2:0] way_id_o;
  wire way_id_o_2_;
  assign way_id_o_2_ = lru_i[0];
  assign way_id_o[2] = way_id_o_2_;

  bsg_mux_width_p1_els_p2
  \lru.rank_1_.nz.mux 
  (
    .data_i(lru_i[2:1]),
    .sel_i(way_id_o_2_),
    .data_o(way_id_o[1])
  );


  bsg_mux_width_p1_els_p4
  \lru.rank_2_.nz.mux 
  (
    .data_i(lru_i[6:3]),
    .sel_i({ way_id_o_2_, way_id_o[1:1] }),
    .data_o(way_id_o[0])
  );


endmodule



module bsg_scan_00000008_1_1
(
  i,
  o
);

  input [7:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__7_,t_1__6_,
  t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__7_ = i[0] | 1'b0;
  assign t_1__6_ = i[1] | i[0];
  assign t_1__5_ = i[2] | i[1];
  assign t_1__4_ = i[3] | i[2];
  assign t_1__3_ = i[4] | i[3];
  assign t_1__2_ = i[5] | i[4];
  assign t_1__1_ = i[6] | i[5];
  assign t_1__0_ = i[7] | i[6];
  assign t_2__7_ = t_1__7_ | 1'b0;
  assign t_2__6_ = t_1__6_ | 1'b0;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign o[0] = t_2__7_ | 1'b0;
  assign o[1] = t_2__6_ | 1'b0;
  assign o[2] = t_2__5_ | 1'b0;
  assign o[3] = t_2__4_ | 1'b0;
  assign o[4] = t_2__3_ | t_2__7_;
  assign o[5] = t_2__2_ | t_2__6_;
  assign o[6] = t_2__1_ | t_2__5_;
  assign o[7] = t_2__0_ | t_2__4_;

endmodule



module bsg_priority_encode_one_hot_out_00000008_1
(
  i,
  o,
  v_o
);

  input [7:0] i;
  output [7:0] o;
  output v_o;
  wire [7:0] o;
  wire v_o,N0,N1,N2,N3,N4,N5,N6;
  wire [6:1] scan_lo;

  bsg_scan_00000008_1_1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, scan_lo, o[0:0] })
  );

  assign o[7] = v_o & N0;
  assign N0 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N1;
  assign N1 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N2;
  assign N2 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N3;
  assign N3 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N4;
  assign N4 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N5;
  assign N5 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N6;
  assign N6 = ~o[0];

endmodule



module bsg_encode_one_hot_00000008_1
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o,v_2__0_,v_1__6_,v_1__4_,v_1__2_,v_1__0_,addr_2__4_,addr_2__0_;
  assign v_1__0_ = i[1] | i[0];
  assign v_1__2_ = i[3] | i[2];
  assign v_1__4_ = i[5] | i[4];
  assign v_1__6_ = i[7] | i[6];
  assign v_2__0_ = v_1__2_ | v_1__0_;
  assign addr_2__0_ = i[1] | i[3];
  assign addr_o[2] = v_1__6_ | v_1__4_;
  assign addr_2__4_ = i[5] | i[7];
  assign v_o = addr_o[2] | v_2__0_;
  assign addr_o[1] = v_1__2_ | v_1__6_;
  assign addr_o[0] = addr_2__0_ | addr_2__4_;

endmodule



module bsg_priority_encode_00000008_1
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [7:0] enc_lo;

  bsg_priority_encode_one_hot_out_00000008_1
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_00000008_1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o)
  );


endmodule



module bsg_decode_00000008
(
  i,
  o
);

  input [2:0] i;
  output [7:0] o;
  wire [7:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_encode_one_hot_00000008
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o,v_2__0_,v_1__6_,v_1__4_,v_1__2_,v_1__0_,addr_2__4_,addr_2__0_;
  assign v_1__0_ = i[1] | i[0];
  assign v_1__2_ = i[3] | i[2];
  assign v_1__4_ = i[5] | i[4];
  assign v_1__6_ = i[7] | i[6];
  assign v_2__0_ = v_1__2_ | v_1__0_;
  assign addr_2__0_ = i[1] | i[3];
  assign addr_o[2] = v_1__6_ | v_1__4_;
  assign addr_2__4_ = i[5] | i[7];
  assign v_o = addr_o[2] | v_2__0_;
  assign addr_o[1] = v_1__2_ | v_1__6_;
  assign addr_o[0] = addr_2__0_ | addr_2__4_;

endmodule



module bsg_lru_pseudo_tree_decode_00000008
(
  way_id_i,
  data_o,
  mask_o
);

  input [2:0] way_id_i;
  output [6:0] data_o;
  output [6:0] mask_o;
  wire [6:0] data_o,mask_o;
  wire N0,N1,N2;
  assign mask_o[0] = 1'b1;
  assign data_o[0] = 1'b1 & N0;
  assign N0 = ~way_id_i[2];
  assign mask_o[1] = 1'b1 & N0;
  assign data_o[1] = mask_o[1] & N1;
  assign N1 = ~way_id_i[1];
  assign mask_o[2] = 1'b1 & way_id_i[2];
  assign data_o[2] = mask_o[2] & N1;
  assign mask_o[3] = mask_o[1] & N1;
  assign data_o[3] = mask_o[3] & N2;
  assign N2 = ~way_id_i[0];
  assign mask_o[4] = mask_o[1] & way_id_i[1];
  assign data_o[4] = mask_o[4] & N2;
  assign mask_o[5] = mask_o[2] & N1;
  assign data_o[5] = mask_o[5] & N2;
  assign mask_o[6] = mask_o[2] & way_id_i[1];
  assign data_o[6] = mask_o[6] & N2;

endmodule



module bsg_mux_segmented_00000007_1
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [6:0] data0_i;
  input [6:0] data1_i;
  input [6:0] sel_i;
  output [6:0] data_o;
  wire [6:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;
  assign data_o[0] = (N0)? data1_i[0] : 
                     (N7)? data0_i[0] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[1] = (N1)? data1_i[1] : 
                     (N8)? data0_i[1] : 1'b0;
  assign N1 = sel_i[1];
  assign data_o[2] = (N2)? data1_i[2] : 
                     (N9)? data0_i[2] : 1'b0;
  assign N2 = sel_i[2];
  assign data_o[3] = (N3)? data1_i[3] : 
                     (N10)? data0_i[3] : 1'b0;
  assign N3 = sel_i[3];
  assign data_o[4] = (N4)? data1_i[4] : 
                     (N11)? data0_i[4] : 1'b0;
  assign N4 = sel_i[4];
  assign data_o[5] = (N5)? data1_i[5] : 
                     (N12)? data0_i[5] : 1'b0;
  assign N5 = sel_i[5];
  assign data_o[6] = (N6)? data1_i[6] : 
                     (N13)? data0_i[6] : 1'b0;
  assign N6 = sel_i[6];
  assign N7 = ~sel_i[0];
  assign N8 = ~sel_i[1];
  assign N9 = ~sel_i[2];
  assign N10 = ~sel_i[3];
  assign N11 = ~sel_i[4];
  assign N12 = ~sel_i[5];
  assign N13 = ~sel_i[6];

endmodule



module bsg_mux_bitwise_00000007
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [6:0] data0_i;
  input [6:0] data1_i;
  input [6:0] sel_i;
  output [6:0] data_o;
  wire [6:0] data_o;

  bsg_mux_segmented_00000007_1
  mux_segmented
  (
    .data0_i(data0_i),
    .data1_i(data1_i),
    .sel_i(sel_i),
    .data_o(data_o)
  );


endmodule



module bsg_cam_1r1w_replacement_00000008
(
  clk_i,
  reset_i,
  read_v_i,
  alloc_v_i,
  alloc_empty_i,
  alloc_v_o
);

  input [7:0] read_v_i;
  input [7:0] alloc_empty_i;
  output [7:0] alloc_v_o;
  input clk_i;
  input reset_i;
  input alloc_v_i;
  wire [7:0] alloc_v_o;
  wire N0,N1,\lru.read_v_li ,\lru.lru_touch_li ,\lru.empty_way_v_lo ,N2,N3,N4,N5,N6,N7,
  N8;
  wire [6:0] \lru.lru_r ,\lru.read_update_data_lo ,\lru.read_update_mask_lo ,
  \lru.read_sel_lo ,\lru.read_update_lo ,\lru.alloc_update_data_lo ,\lru.alloc_update_mask_lo ,
  \lru.alloc_sel_lo ,\lru.alloc_update_lo ;
  wire [2:0] \lru.lru_way_lo ,\lru.empty_way_lo ,\lru.way_lo ,\lru.read_way_li ;

  bsg_dff_reset_en_00000007
  \lru.lru_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(\lru.lru_touch_li ),
    .data_i(\lru.alloc_update_lo ),
    .data_o(\lru.lru_r )
  );


  bsg_lru_pseudo_tree_encode_00000008
  \lru.lru_encoder 
  (
    .lru_i(\lru.lru_r ),
    .way_id_o(\lru.lru_way_lo )
  );


  bsg_priority_encode_00000008_1
  \lru.empty_encoder 
  (
    .i(alloc_empty_i),
    .addr_o(\lru.empty_way_lo ),
    .v_o(\lru.empty_way_v_lo )
  );


  bsg_decode_00000008
  \lru.way_decoder 
  (
    .i(\lru.way_lo ),
    .o(alloc_v_o)
  );


  bsg_encode_one_hot_00000008
  \lru.read_way_encoder 
  (
    .i(read_v_i),
    .addr_o(\lru.read_way_li )
  );


  bsg_lru_pseudo_tree_decode_00000008
  \lru.read_decoder 
  (
    .way_id_i(\lru.read_way_li ),
    .data_o(\lru.read_update_data_lo ),
    .mask_o(\lru.read_update_mask_lo )
  );


  bsg_mux_bitwise_00000007
  \lru.read_update_mux 
  (
    .data0_i(\lru.lru_r ),
    .data1_i(\lru.read_update_data_lo ),
    .sel_i(\lru.read_sel_lo ),
    .data_o(\lru.read_update_lo )
  );


  bsg_lru_pseudo_tree_decode_00000008
  \lru.alloc_decoder 
  (
    .way_id_i(\lru.way_lo ),
    .data_o(\lru.alloc_update_data_lo ),
    .mask_o(\lru.alloc_update_mask_lo )
  );


  bsg_mux_bitwise_00000007
  \lru.alloc_update_mux 
  (
    .data0_i(\lru.read_update_lo ),
    .data1_i(\lru.alloc_update_data_lo ),
    .sel_i(\lru.alloc_sel_lo ),
    .data_o(\lru.alloc_update_lo )
  );

  assign \lru.way_lo  = (N0)? \lru.empty_way_lo  : 
                        (N1)? \lru.lru_way_lo  : 1'b0;
  assign N0 = \lru.empty_way_v_lo ;
  assign N1 = N2;
  assign \lru.read_v_li  = N8 | read_v_i[0];
  assign N8 = N7 | read_v_i[1];
  assign N7 = N6 | read_v_i[2];
  assign N6 = N5 | read_v_i[3];
  assign N5 = N4 | read_v_i[4];
  assign N4 = N3 | read_v_i[5];
  assign N3 = read_v_i[7] | read_v_i[6];
  assign \lru.lru_touch_li  = \lru.read_v_li  | alloc_v_i;
  assign N2 = ~\lru.empty_way_v_lo ;
  assign \lru.read_sel_lo [6] = \lru.read_update_mask_lo [6] & \lru.read_v_li ;
  assign \lru.read_sel_lo [5] = \lru.read_update_mask_lo [5] & \lru.read_v_li ;
  assign \lru.read_sel_lo [4] = \lru.read_update_mask_lo [4] & \lru.read_v_li ;
  assign \lru.read_sel_lo [3] = \lru.read_update_mask_lo [3] & \lru.read_v_li ;
  assign \lru.read_sel_lo [2] = \lru.read_update_mask_lo [2] & \lru.read_v_li ;
  assign \lru.read_sel_lo [1] = \lru.read_update_mask_lo [1] & \lru.read_v_li ;
  assign \lru.read_sel_lo [0] = \lru.read_update_mask_lo [0] & \lru.read_v_li ;
  assign \lru.alloc_sel_lo [6] = \lru.alloc_update_mask_lo [6] & alloc_v_i;
  assign \lru.alloc_sel_lo [5] = \lru.alloc_update_mask_lo [5] & alloc_v_i;
  assign \lru.alloc_sel_lo [4] = \lru.alloc_update_mask_lo [4] & alloc_v_i;
  assign \lru.alloc_sel_lo [3] = \lru.alloc_update_mask_lo [3] & alloc_v_i;
  assign \lru.alloc_sel_lo [2] = \lru.alloc_update_mask_lo [2] & alloc_v_i;
  assign \lru.alloc_sel_lo [1] = \lru.alloc_update_mask_lo [1] & alloc_v_i;
  assign \lru.alloc_sel_lo [0] = \lru.alloc_update_mask_lo [0] & alloc_v_i;

endmodule



module bsg_cam_1r1w_tag_array_0000001b_00000002
(
  clk_i,
  reset_i,
  w_v_i,
  w_set_not_clear_i,
  w_tag_i,
  w_empty_o,
  r_v_i,
  r_tag_i,
  r_match_o
);

  input [1:0] w_v_i;
  input [26:0] w_tag_i;
  output [1:0] w_empty_o;
  input [26:0] r_tag_i;
  output [1:0] r_match_o;
  input clk_i;
  input reset_i;
  input w_set_not_clear_i;
  input r_v_i;
  wire [1:0] w_empty_o,r_match_o,v_r;
  wire _0_net_,N0,_1_net_,N1,N2,N3;
  wire [53:0] tag_r;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_0_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[0]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[0])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_0_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_0_net_),
    .data_o(tag_r[26:0])
  );

  assign N0 = tag_r[26:0] == r_tag_i;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_1_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[1]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[1])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_1_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_1_net_),
    .data_o(tag_r[53:27])
  );

  assign N1 = tag_r[53:27] == r_tag_i;
  assign _0_net_ = w_v_i[0] & w_set_not_clear_i;
  assign r_match_o[0] = N2 & N0;
  assign N2 = r_v_i & v_r[0];
  assign w_empty_o[0] = ~v_r[0];
  assign _1_net_ = w_v_i[1] & w_set_not_clear_i;
  assign r_match_o[1] = N3 & N1;
  assign N3 = r_v_i & v_r[1];
  assign w_empty_o[1] = ~v_r[1];

endmodule



module bsg_lru_pseudo_tree_encode_00000002
(
  lru_i,
  way_id_o
);

  input [0:0] lru_i;
  output [0:0] way_id_o;
  wire [0:0] way_id_o;
  assign way_id_o[0] = lru_i[0];

endmodule



module bsg_scan_00000002_1_1
(
  i,
  o
);

  input [1:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o[0] = i[0] | 1'b0;
  assign o[1] = i[1] | i[0];

endmodule



module bsg_priority_encode_one_hot_out_00000002_1
(
  i,
  o,
  v_o
);

  input [1:0] i;
  output [1:0] o;
  output v_o;
  wire [1:0] o;
  wire v_o,N0;

  bsg_scan_00000002_1_1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, o[0:0] })
  );

  assign o[1] = v_o & N0;
  assign N0 = ~o[0];

endmodule



module bsg_encode_one_hot_00000002_1
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign addr_o[0] = i[1];
  assign v_o = addr_o[0] | i[0];

endmodule



module bsg_priority_encode_00000002_1
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  wire [1:0] enc_lo;

  bsg_priority_encode_one_hot_out_00000002_1
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_00000002_1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o[0])
  );


endmodule



module bsg_decode_num_out_p2
(
  i,
  o
);

  input [0:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o = { 1'b0, 1'b1 } << i[0];

endmodule



module bsg_encode_one_hot_00000002
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign addr_o[0] = i[1];
  assign v_o = addr_o[0] | i[0];

endmodule



module bsg_lru_pseudo_tree_decode_00000002
(
  way_id_i,
  data_o,
  mask_o
);

  input [0:0] way_id_i;
  output [0:0] data_o;
  output [0:0] mask_o;
  wire [0:0] data_o,mask_o;
  wire N0;
  assign mask_o[0] = 1'b1;
  assign data_o[0] = 1'b1 & N0;
  assign N0 = ~way_id_i[0];

endmodule



module bsg_mux_segmented_00000001_1
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [0:0] data0_i;
  input [0:0] data1_i;
  input [0:0] sel_i;
  output [0:0] data_o;
  wire [0:0] data_o;
  wire N0,N1;
  assign data_o[0] = (N0)? data1_i[0] : 
                     (N1)? data0_i[0] : 1'b0;
  assign N0 = sel_i[0];
  assign N1 = ~sel_i[0];

endmodule



module bsg_mux_bitwise_00000001
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [0:0] data0_i;
  input [0:0] data1_i;
  input [0:0] sel_i;
  output [0:0] data_o;
  wire [0:0] data_o;

  bsg_mux_segmented_00000001_1
  mux_segmented
  (
    .data0_i(data0_i[0]),
    .data1_i(data1_i[0]),
    .sel_i(sel_i[0]),
    .data_o(data_o[0])
  );


endmodule



module bsg_cam_1r1w_replacement_00000002
(
  clk_i,
  reset_i,
  read_v_i,
  alloc_v_i,
  alloc_empty_i,
  alloc_v_o
);

  input [1:0] read_v_i;
  input [1:0] alloc_empty_i;
  output [1:0] alloc_v_o;
  input clk_i;
  input reset_i;
  input alloc_v_i;
  wire [1:0] alloc_v_o;
  wire N0,N1,\lru.read_v_li ,\lru.lru_touch_li ,\lru.empty_way_v_lo ,N2;
  wire [0:0] \lru.lru_r ,\lru.lru_way_lo ,\lru.empty_way_lo ,\lru.way_lo ,\lru.read_way_li ,
  \lru.read_update_data_lo ,\lru.read_update_mask_lo ,\lru.read_sel_lo ,
  \lru.read_update_lo ,\lru.alloc_update_data_lo ,\lru.alloc_update_mask_lo ,
  \lru.alloc_sel_lo ,\lru.alloc_update_lo ;

  bsg_dff_reset_en_width_p1
  \lru.lru_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(\lru.lru_touch_li ),
    .data_i(\lru.alloc_update_lo [0]),
    .data_o(\lru.lru_r [0])
  );


  bsg_lru_pseudo_tree_encode_00000002
  \lru.lru_encoder 
  (
    .lru_i(\lru.lru_r [0]),
    .way_id_o(\lru.lru_way_lo [0])
  );


  bsg_priority_encode_00000002_1
  \lru.empty_encoder 
  (
    .i(alloc_empty_i),
    .addr_o(\lru.empty_way_lo [0]),
    .v_o(\lru.empty_way_v_lo )
  );


  bsg_decode_num_out_p2
  \lru.way_decoder 
  (
    .i(\lru.way_lo [0]),
    .o(alloc_v_o)
  );


  bsg_encode_one_hot_00000002
  \lru.read_way_encoder 
  (
    .i(read_v_i),
    .addr_o(\lru.read_way_li [0])
  );


  bsg_lru_pseudo_tree_decode_00000002
  \lru.read_decoder 
  (
    .way_id_i(\lru.read_way_li [0]),
    .data_o(\lru.read_update_data_lo [0]),
    .mask_o(\lru.read_update_mask_lo [0])
  );


  bsg_mux_bitwise_00000001
  \lru.read_update_mux 
  (
    .data0_i(\lru.lru_r [0]),
    .data1_i(\lru.read_update_data_lo [0]),
    .sel_i(\lru.read_sel_lo [0]),
    .data_o(\lru.read_update_lo [0])
  );


  bsg_lru_pseudo_tree_decode_00000002
  \lru.alloc_decoder 
  (
    .way_id_i(\lru.way_lo [0]),
    .data_o(\lru.alloc_update_data_lo [0]),
    .mask_o(\lru.alloc_update_mask_lo [0])
  );


  bsg_mux_bitwise_00000001
  \lru.alloc_update_mux 
  (
    .data0_i(\lru.read_update_lo [0]),
    .data1_i(\lru.alloc_update_data_lo [0]),
    .sel_i(\lru.alloc_sel_lo [0]),
    .data_o(\lru.alloc_update_lo [0])
  );

  assign \lru.way_lo [0] = (N0)? \lru.empty_way_lo [0] : 
                           (N1)? \lru.lru_way_lo [0] : 1'b0;
  assign N0 = \lru.empty_way_v_lo ;
  assign N1 = N2;
  assign \lru.read_v_li  = read_v_i[1] | read_v_i[0];
  assign \lru.lru_touch_li  = \lru.read_v_li  | alloc_v_i;
  assign N2 = ~\lru.empty_way_v_lo ;
  assign \lru.read_sel_lo [0] = \lru.read_update_mask_lo [0] & \lru.read_v_li ;
  assign \lru.alloc_sel_lo [0] = \lru.alloc_update_mask_lo [0] & alloc_v_i;

endmodule



module bsg_cam_1r1w_tag_array_0000001b_00000001
(
  clk_i,
  reset_i,
  w_v_i,
  w_set_not_clear_i,
  w_tag_i,
  w_empty_o,
  r_v_i,
  r_tag_i,
  r_match_o
);

  input [0:0] w_v_i;
  input [26:0] w_tag_i;
  output [0:0] w_empty_o;
  input [26:0] r_tag_i;
  output [0:0] r_match_o;
  input clk_i;
  input reset_i;
  input w_set_not_clear_i;
  input r_v_i;
  wire [0:0] w_empty_o,r_match_o,v_r;
  wire _0_net_,N0,N1;
  wire [26:0] tag_r;

  bsg_dff_reset_en_width_p1
  \nz.tag_array_0_.v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(w_v_i[0]),
    .data_i(w_set_not_clear_i),
    .data_o(v_r[0])
  );


  bsg_dff_en_0000001b
  \nz.tag_array_0_.tag_r_reg 
  (
    .clk_i(clk_i),
    .data_i(w_tag_i),
    .en_i(_0_net_),
    .data_o(tag_r)
  );

  assign N0 = tag_r == r_tag_i;
  assign _0_net_ = w_v_i[0] & w_set_not_clear_i;
  assign r_match_o[0] = N1 & N0;
  assign N1 = r_v_i & v_r[0];
  assign w_empty_o[0] = ~v_r[0];

endmodule



module bsg_cam_1r1w_replacement_00000001
(
  clk_i,
  reset_i,
  read_v_i,
  alloc_v_i,
  alloc_empty_i,
  alloc_v_o
);

  input [0:0] read_v_i;
  input [0:0] alloc_empty_i;
  output [0:0] alloc_v_o;
  input clk_i;
  input reset_i;
  input alloc_v_i;
  wire [0:0] alloc_v_o;
  assign alloc_v_o[0] = 1'b1;

endmodule



module bsg_dff_en_00000024
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [35:0] data_i;
  output [35:0] data_o;
  input clk_i;
  input en_i;
  wire [35:0] data_o;
  reg data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,
  data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,
  data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,
  data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_width_p18
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [17:0] data_i;
  output [17:0] data_o;
  input clk_i;
  input en_i;
  wire [17:0] data_o;
  reg data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,
  data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mux_one_hot_9_00000009
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [80:0] data_i;
  input [8:0] sel_one_hot_i;
  output [8:0] data_o;
  wire [8:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62;
  wire [80:0] data_masked;
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[1];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[1];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[1];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[1];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[1];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[1];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[1];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[1];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[1];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[2];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[2];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[2];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[2];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[2];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[2];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[2];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[2];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[2];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[3];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[3];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[3];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[3];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[3];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[3];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[3];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[3];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[3];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[4];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[4];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[4];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[4];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[4];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[4];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[4];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[4];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[4];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[5];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[5];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[5];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[5];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[5];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[5];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[5];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[5];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[5];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[6];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[6];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[6];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[6];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[6];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[6];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[6];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[6];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[6];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[7];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[7];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[7];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[7];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[7];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[7];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[7];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[7];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[7];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[8];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[8];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[8];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[8];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[8];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[8];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[8];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[8];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[8];
  assign data_o[0] = N6 | data_masked[0];
  assign N6 = N5 | data_masked[9];
  assign N5 = N4 | data_masked[18];
  assign N4 = N3 | data_masked[27];
  assign N3 = N2 | data_masked[36];
  assign N2 = N1 | data_masked[45];
  assign N1 = N0 | data_masked[54];
  assign N0 = data_masked[72] | data_masked[63];
  assign data_o[1] = N13 | data_masked[1];
  assign N13 = N12 | data_masked[10];
  assign N12 = N11 | data_masked[19];
  assign N11 = N10 | data_masked[28];
  assign N10 = N9 | data_masked[37];
  assign N9 = N8 | data_masked[46];
  assign N8 = N7 | data_masked[55];
  assign N7 = data_masked[73] | data_masked[64];
  assign data_o[2] = N20 | data_masked[2];
  assign N20 = N19 | data_masked[11];
  assign N19 = N18 | data_masked[20];
  assign N18 = N17 | data_masked[29];
  assign N17 = N16 | data_masked[38];
  assign N16 = N15 | data_masked[47];
  assign N15 = N14 | data_masked[56];
  assign N14 = data_masked[74] | data_masked[65];
  assign data_o[3] = N27 | data_masked[3];
  assign N27 = N26 | data_masked[12];
  assign N26 = N25 | data_masked[21];
  assign N25 = N24 | data_masked[30];
  assign N24 = N23 | data_masked[39];
  assign N23 = N22 | data_masked[48];
  assign N22 = N21 | data_masked[57];
  assign N21 = data_masked[75] | data_masked[66];
  assign data_o[4] = N34 | data_masked[4];
  assign N34 = N33 | data_masked[13];
  assign N33 = N32 | data_masked[22];
  assign N32 = N31 | data_masked[31];
  assign N31 = N30 | data_masked[40];
  assign N30 = N29 | data_masked[49];
  assign N29 = N28 | data_masked[58];
  assign N28 = data_masked[76] | data_masked[67];
  assign data_o[5] = N41 | data_masked[5];
  assign N41 = N40 | data_masked[14];
  assign N40 = N39 | data_masked[23];
  assign N39 = N38 | data_masked[32];
  assign N38 = N37 | data_masked[41];
  assign N37 = N36 | data_masked[50];
  assign N36 = N35 | data_masked[59];
  assign N35 = data_masked[77] | data_masked[68];
  assign data_o[6] = N48 | data_masked[6];
  assign N48 = N47 | data_masked[15];
  assign N47 = N46 | data_masked[24];
  assign N46 = N45 | data_masked[33];
  assign N45 = N44 | data_masked[42];
  assign N44 = N43 | data_masked[51];
  assign N43 = N42 | data_masked[60];
  assign N42 = data_masked[78] | data_masked[69];
  assign data_o[7] = N55 | data_masked[7];
  assign N55 = N54 | data_masked[16];
  assign N54 = N53 | data_masked[25];
  assign N53 = N52 | data_masked[34];
  assign N52 = N51 | data_masked[43];
  assign N51 = N50 | data_masked[52];
  assign N50 = N49 | data_masked[61];
  assign N49 = data_masked[79] | data_masked[70];
  assign data_o[8] = N62 | data_masked[8];
  assign N62 = N61 | data_masked[17];
  assign N61 = N60 | data_masked[26];
  assign N60 = N59 | data_masked[35];
  assign N59 = N58 | data_masked[44];
  assign N58 = N57 | data_masked[53];
  assign N57 = N56 | data_masked[62];
  assign N56 = data_masked[80] | data_masked[71];

endmodule



module bsg_mux_one_hot_9_0000000b
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [98:0] data_i;
  input [10:0] sel_one_hot_i;
  output [8:0] data_o;
  wire [8:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80;
  wire [98:0] data_masked;
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[1];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[1];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[1];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[1];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[1];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[1];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[1];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[1];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[1];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[2];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[2];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[2];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[2];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[2];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[2];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[2];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[2];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[2];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[3];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[3];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[3];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[3];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[3];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[3];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[3];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[3];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[3];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[4];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[4];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[4];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[4];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[4];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[4];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[4];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[4];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[4];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[5];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[5];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[5];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[5];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[5];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[5];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[5];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[5];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[5];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[6];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[6];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[6];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[6];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[6];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[6];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[6];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[6];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[6];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[7];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[7];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[7];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[7];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[7];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[7];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[7];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[7];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[7];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[8];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[8];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[8];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[8];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[8];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[8];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[8];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[8];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[8];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[9];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[9];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[9];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[9];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[9];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[9];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[9];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[9];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[9];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[10];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[10];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[10];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[10];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[10];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[10];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[10];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[10];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[10];
  assign data_o[0] = N8 | data_masked[0];
  assign N8 = N7 | data_masked[9];
  assign N7 = N6 | data_masked[18];
  assign N6 = N5 | data_masked[27];
  assign N5 = N4 | data_masked[36];
  assign N4 = N3 | data_masked[45];
  assign N3 = N2 | data_masked[54];
  assign N2 = N1 | data_masked[63];
  assign N1 = N0 | data_masked[72];
  assign N0 = data_masked[90] | data_masked[81];
  assign data_o[1] = N17 | data_masked[1];
  assign N17 = N16 | data_masked[10];
  assign N16 = N15 | data_masked[19];
  assign N15 = N14 | data_masked[28];
  assign N14 = N13 | data_masked[37];
  assign N13 = N12 | data_masked[46];
  assign N12 = N11 | data_masked[55];
  assign N11 = N10 | data_masked[64];
  assign N10 = N9 | data_masked[73];
  assign N9 = data_masked[91] | data_masked[82];
  assign data_o[2] = N26 | data_masked[2];
  assign N26 = N25 | data_masked[11];
  assign N25 = N24 | data_masked[20];
  assign N24 = N23 | data_masked[29];
  assign N23 = N22 | data_masked[38];
  assign N22 = N21 | data_masked[47];
  assign N21 = N20 | data_masked[56];
  assign N20 = N19 | data_masked[65];
  assign N19 = N18 | data_masked[74];
  assign N18 = data_masked[92] | data_masked[83];
  assign data_o[3] = N35 | data_masked[3];
  assign N35 = N34 | data_masked[12];
  assign N34 = N33 | data_masked[21];
  assign N33 = N32 | data_masked[30];
  assign N32 = N31 | data_masked[39];
  assign N31 = N30 | data_masked[48];
  assign N30 = N29 | data_masked[57];
  assign N29 = N28 | data_masked[66];
  assign N28 = N27 | data_masked[75];
  assign N27 = data_masked[93] | data_masked[84];
  assign data_o[4] = N44 | data_masked[4];
  assign N44 = N43 | data_masked[13];
  assign N43 = N42 | data_masked[22];
  assign N42 = N41 | data_masked[31];
  assign N41 = N40 | data_masked[40];
  assign N40 = N39 | data_masked[49];
  assign N39 = N38 | data_masked[58];
  assign N38 = N37 | data_masked[67];
  assign N37 = N36 | data_masked[76];
  assign N36 = data_masked[94] | data_masked[85];
  assign data_o[5] = N53 | data_masked[5];
  assign N53 = N52 | data_masked[14];
  assign N52 = N51 | data_masked[23];
  assign N51 = N50 | data_masked[32];
  assign N50 = N49 | data_masked[41];
  assign N49 = N48 | data_masked[50];
  assign N48 = N47 | data_masked[59];
  assign N47 = N46 | data_masked[68];
  assign N46 = N45 | data_masked[77];
  assign N45 = data_masked[95] | data_masked[86];
  assign data_o[6] = N62 | data_masked[6];
  assign N62 = N61 | data_masked[15];
  assign N61 = N60 | data_masked[24];
  assign N60 = N59 | data_masked[33];
  assign N59 = N58 | data_masked[42];
  assign N58 = N57 | data_masked[51];
  assign N57 = N56 | data_masked[60];
  assign N56 = N55 | data_masked[69];
  assign N55 = N54 | data_masked[78];
  assign N54 = data_masked[96] | data_masked[87];
  assign data_o[7] = N71 | data_masked[7];
  assign N71 = N70 | data_masked[16];
  assign N70 = N69 | data_masked[25];
  assign N69 = N68 | data_masked[34];
  assign N68 = N67 | data_masked[43];
  assign N67 = N66 | data_masked[52];
  assign N66 = N65 | data_masked[61];
  assign N65 = N64 | data_masked[70];
  assign N64 = N63 | data_masked[79];
  assign N63 = data_masked[97] | data_masked[88];
  assign data_o[8] = N80 | data_masked[8];
  assign N80 = N79 | data_masked[17];
  assign N79 = N78 | data_masked[26];
  assign N78 = N77 | data_masked[35];
  assign N77 = N76 | data_masked[44];
  assign N76 = N75 | data_masked[53];
  assign N75 = N74 | data_masked[62];
  assign N74 = N73 | data_masked[71];
  assign N73 = N72 | data_masked[80];
  assign N72 = data_masked[98] | data_masked[89];

endmodule



module bsg_mux_one_hot_18_0000000b
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [197:0] data_i;
  input [10:0] sel_one_hot_i;
  output [17:0] data_o;
  wire [17:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161;
  wire [197:0] data_masked;
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[1];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[1];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[1];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[1];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[1];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[1];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[1];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[1];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[1];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[1];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[1];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[1];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[1];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[1];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[1];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[1];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[1];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[1];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[2];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[2];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[2];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[2];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[2];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[2];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[2];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[2];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[2];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[2];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[2];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[2];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[2];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[2];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[2];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[2];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[2];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[2];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[3];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[3];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[3];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[3];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[3];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[3];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[3];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[3];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[3];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[3];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[3];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[3];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[3];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[3];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[3];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[3];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[3];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[3];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[4];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[4];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[4];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[4];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[4];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[4];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[4];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[4];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[4];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[4];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[4];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[4];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[4];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[4];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[4];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[4];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[4];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[4];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[5];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[5];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[5];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[5];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[5];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[5];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[5];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[5];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[5];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[5];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[5];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[5];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[5];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[5];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[5];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[5];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[5];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[5];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[6];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[6];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[6];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[6];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[6];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[6];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[6];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[6];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[6];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[6];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[6];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[6];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[6];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[6];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[6];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[6];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[6];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[6];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[7];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[7];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[7];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[7];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[7];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[7];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[7];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[7];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[7];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[7];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[7];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[7];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[7];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[7];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[7];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[7];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[7];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[7];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[8];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[8];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[8];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[8];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[8];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[8];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[8];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[8];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[8];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[8];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[8];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[8];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[8];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[8];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[8];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[8];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[8];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[8];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[9];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[9];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[9];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[9];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[9];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[9];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[9];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[9];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[9];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[9];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[9];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[9];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[9];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[9];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[9];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[9];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[9];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[9];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[10];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[10];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[10];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[10];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[10];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[10];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[10];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[10];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[10];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[10];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[10];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[10];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[10];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[10];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[10];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[10];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[10];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[10];
  assign data_o[0] = N8 | data_masked[0];
  assign N8 = N7 | data_masked[18];
  assign N7 = N6 | data_masked[36];
  assign N6 = N5 | data_masked[54];
  assign N5 = N4 | data_masked[72];
  assign N4 = N3 | data_masked[90];
  assign N3 = N2 | data_masked[108];
  assign N2 = N1 | data_masked[126];
  assign N1 = N0 | data_masked[144];
  assign N0 = data_masked[180] | data_masked[162];
  assign data_o[1] = N17 | data_masked[1];
  assign N17 = N16 | data_masked[19];
  assign N16 = N15 | data_masked[37];
  assign N15 = N14 | data_masked[55];
  assign N14 = N13 | data_masked[73];
  assign N13 = N12 | data_masked[91];
  assign N12 = N11 | data_masked[109];
  assign N11 = N10 | data_masked[127];
  assign N10 = N9 | data_masked[145];
  assign N9 = data_masked[181] | data_masked[163];
  assign data_o[2] = N26 | data_masked[2];
  assign N26 = N25 | data_masked[20];
  assign N25 = N24 | data_masked[38];
  assign N24 = N23 | data_masked[56];
  assign N23 = N22 | data_masked[74];
  assign N22 = N21 | data_masked[92];
  assign N21 = N20 | data_masked[110];
  assign N20 = N19 | data_masked[128];
  assign N19 = N18 | data_masked[146];
  assign N18 = data_masked[182] | data_masked[164];
  assign data_o[3] = N35 | data_masked[3];
  assign N35 = N34 | data_masked[21];
  assign N34 = N33 | data_masked[39];
  assign N33 = N32 | data_masked[57];
  assign N32 = N31 | data_masked[75];
  assign N31 = N30 | data_masked[93];
  assign N30 = N29 | data_masked[111];
  assign N29 = N28 | data_masked[129];
  assign N28 = N27 | data_masked[147];
  assign N27 = data_masked[183] | data_masked[165];
  assign data_o[4] = N44 | data_masked[4];
  assign N44 = N43 | data_masked[22];
  assign N43 = N42 | data_masked[40];
  assign N42 = N41 | data_masked[58];
  assign N41 = N40 | data_masked[76];
  assign N40 = N39 | data_masked[94];
  assign N39 = N38 | data_masked[112];
  assign N38 = N37 | data_masked[130];
  assign N37 = N36 | data_masked[148];
  assign N36 = data_masked[184] | data_masked[166];
  assign data_o[5] = N53 | data_masked[5];
  assign N53 = N52 | data_masked[23];
  assign N52 = N51 | data_masked[41];
  assign N51 = N50 | data_masked[59];
  assign N50 = N49 | data_masked[77];
  assign N49 = N48 | data_masked[95];
  assign N48 = N47 | data_masked[113];
  assign N47 = N46 | data_masked[131];
  assign N46 = N45 | data_masked[149];
  assign N45 = data_masked[185] | data_masked[167];
  assign data_o[6] = N62 | data_masked[6];
  assign N62 = N61 | data_masked[24];
  assign N61 = N60 | data_masked[42];
  assign N60 = N59 | data_masked[60];
  assign N59 = N58 | data_masked[78];
  assign N58 = N57 | data_masked[96];
  assign N57 = N56 | data_masked[114];
  assign N56 = N55 | data_masked[132];
  assign N55 = N54 | data_masked[150];
  assign N54 = data_masked[186] | data_masked[168];
  assign data_o[7] = N71 | data_masked[7];
  assign N71 = N70 | data_masked[25];
  assign N70 = N69 | data_masked[43];
  assign N69 = N68 | data_masked[61];
  assign N68 = N67 | data_masked[79];
  assign N67 = N66 | data_masked[97];
  assign N66 = N65 | data_masked[115];
  assign N65 = N64 | data_masked[133];
  assign N64 = N63 | data_masked[151];
  assign N63 = data_masked[187] | data_masked[169];
  assign data_o[8] = N80 | data_masked[8];
  assign N80 = N79 | data_masked[26];
  assign N79 = N78 | data_masked[44];
  assign N78 = N77 | data_masked[62];
  assign N77 = N76 | data_masked[80];
  assign N76 = N75 | data_masked[98];
  assign N75 = N74 | data_masked[116];
  assign N74 = N73 | data_masked[134];
  assign N73 = N72 | data_masked[152];
  assign N72 = data_masked[188] | data_masked[170];
  assign data_o[9] = N89 | data_masked[9];
  assign N89 = N88 | data_masked[27];
  assign N88 = N87 | data_masked[45];
  assign N87 = N86 | data_masked[63];
  assign N86 = N85 | data_masked[81];
  assign N85 = N84 | data_masked[99];
  assign N84 = N83 | data_masked[117];
  assign N83 = N82 | data_masked[135];
  assign N82 = N81 | data_masked[153];
  assign N81 = data_masked[189] | data_masked[171];
  assign data_o[10] = N98 | data_masked[10];
  assign N98 = N97 | data_masked[28];
  assign N97 = N96 | data_masked[46];
  assign N96 = N95 | data_masked[64];
  assign N95 = N94 | data_masked[82];
  assign N94 = N93 | data_masked[100];
  assign N93 = N92 | data_masked[118];
  assign N92 = N91 | data_masked[136];
  assign N91 = N90 | data_masked[154];
  assign N90 = data_masked[190] | data_masked[172];
  assign data_o[11] = N107 | data_masked[11];
  assign N107 = N106 | data_masked[29];
  assign N106 = N105 | data_masked[47];
  assign N105 = N104 | data_masked[65];
  assign N104 = N103 | data_masked[83];
  assign N103 = N102 | data_masked[101];
  assign N102 = N101 | data_masked[119];
  assign N101 = N100 | data_masked[137];
  assign N100 = N99 | data_masked[155];
  assign N99 = data_masked[191] | data_masked[173];
  assign data_o[12] = N116 | data_masked[12];
  assign N116 = N115 | data_masked[30];
  assign N115 = N114 | data_masked[48];
  assign N114 = N113 | data_masked[66];
  assign N113 = N112 | data_masked[84];
  assign N112 = N111 | data_masked[102];
  assign N111 = N110 | data_masked[120];
  assign N110 = N109 | data_masked[138];
  assign N109 = N108 | data_masked[156];
  assign N108 = data_masked[192] | data_masked[174];
  assign data_o[13] = N125 | data_masked[13];
  assign N125 = N124 | data_masked[31];
  assign N124 = N123 | data_masked[49];
  assign N123 = N122 | data_masked[67];
  assign N122 = N121 | data_masked[85];
  assign N121 = N120 | data_masked[103];
  assign N120 = N119 | data_masked[121];
  assign N119 = N118 | data_masked[139];
  assign N118 = N117 | data_masked[157];
  assign N117 = data_masked[193] | data_masked[175];
  assign data_o[14] = N134 | data_masked[14];
  assign N134 = N133 | data_masked[32];
  assign N133 = N132 | data_masked[50];
  assign N132 = N131 | data_masked[68];
  assign N131 = N130 | data_masked[86];
  assign N130 = N129 | data_masked[104];
  assign N129 = N128 | data_masked[122];
  assign N128 = N127 | data_masked[140];
  assign N127 = N126 | data_masked[158];
  assign N126 = data_masked[194] | data_masked[176];
  assign data_o[15] = N143 | data_masked[15];
  assign N143 = N142 | data_masked[33];
  assign N142 = N141 | data_masked[51];
  assign N141 = N140 | data_masked[69];
  assign N140 = N139 | data_masked[87];
  assign N139 = N138 | data_masked[105];
  assign N138 = N137 | data_masked[123];
  assign N137 = N136 | data_masked[141];
  assign N136 = N135 | data_masked[159];
  assign N135 = data_masked[195] | data_masked[177];
  assign data_o[16] = N152 | data_masked[16];
  assign N152 = N151 | data_masked[34];
  assign N151 = N150 | data_masked[52];
  assign N150 = N149 | data_masked[70];
  assign N149 = N148 | data_masked[88];
  assign N148 = N147 | data_masked[106];
  assign N147 = N146 | data_masked[124];
  assign N146 = N145 | data_masked[142];
  assign N145 = N144 | data_masked[160];
  assign N144 = data_masked[196] | data_masked[178];
  assign data_o[17] = N161 | data_masked[17];
  assign N161 = N160 | data_masked[35];
  assign N160 = N159 | data_masked[53];
  assign N159 = N158 | data_masked[71];
  assign N158 = N157 | data_masked[89];
  assign N157 = N156 | data_masked[107];
  assign N156 = N155 | data_masked[125];
  assign N155 = N154 | data_masked[143];
  assign N154 = N153 | data_masked[161];
  assign N153 = data_masked[197] | data_masked[179];

endmodule



module bsg_popcount_width_p3
(
  i,
  o
);

  input [2:0] i;
  output [1:0] o;
  wire [1:0] o;
  wire N0,N1,N2,N3,N4;
  assign o[0] = N0 ^ i[0];
  assign N0 = i[2] ^ i[1];
  assign o[1] = N3 | N4;
  assign N3 = N1 | N2;
  assign N1 = i[1] & i[0];
  assign N2 = i[2] & i[1];
  assign N4 = i[0] & i[2];

endmodule



module bsg_rotate_right_width_p36
(
  data_i,
  rot_i,
  o
);

  input [35:0] data_i;
  input [5:0] rot_i;
  output [35:0] o;
  wire [35:0] o;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,
  sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,
  sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,sv2v_dc_21,sv2v_dc_22,
  sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,sv2v_dc_27,sv2v_dc_28,sv2v_dc_29,
  sv2v_dc_30,sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,sv2v_dc_34,sv2v_dc_35,sv2v_dc_36;
  assign { sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36, o } = { data_i, data_i } >> rot_i;

endmodule



module bp_tlb_00_00000001_00000002_00000008
(
  clk_i,
  reset_i,
  fence_i,
  v_i,
  w_i,
  vtag_i,
  entry_i,
  v_o,
  entry_o
);

  input [26:0] vtag_i;
  input [35:0] entry_i;
  output [35:0] entry_o;
  input clk_i;
  input reset_i;
  input fence_i;
  input v_i;
  input w_i;
  output v_o;
  wire [35:0] entry_o,entry_shifted,data_2m_high_r,r_entry;
  wire v_o,w_v_li,fill_gigapage,fill_megapage,fill_kilopage,flush_4k_li,_1_net_,
  any_match_4k_lo,flush_2m_li,_3_net_,any_match_2m_lo,_5_net_,_21_net__8_,N0,N1,N3,N4,N5,
  N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26;
  wire [26:0] vtag_r;
  wire [7:0] repl_way_4k_lo,tag_4k_w_v_li,tag_empty_4k_lo,tag_r_match_4k_lo,mem_4k_w_v_li;
  wire [1:0] repl_way_2m_lo,tag_2m_w_v_li,tag_empty_2m_lo,tag_r_match_2m_lo,mem_2m_w_v_li,
  match_cnt;
  wire [0:0] repl_way_1g_lo,tag_1g_w_v_li,tag_empty_1g_lo,tag_r_match_1g_lo,mem_1g_w_v_li;
  wire [143:0] data_4k_high_r;
  wire [71:0] data_4k_med_r,data_4k_low_r;
  wire [17:0] data_2m_med_r,data_1g_high_r;

  bsg_rotate_left_width_p36
  entry_shift
  (
    .data_i(entry_i),
    .rot_i({ 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0 }),
    .o(entry_shifted)
  );


  bsg_dff_en_0000001b
  vtag_reg
  (
    .clk_i(clk_i),
    .data_i(vtag_i),
    .en_i(v_i),
    .data_o(vtag_r)
  );


  bsg_cam_1r1w_tag_array_0000001b_00000008
  tag_array_4k
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(tag_4k_w_v_li),
    .w_set_not_clear_i(_1_net_),
    .w_tag_i(vtag_i),
    .w_empty_o(tag_empty_4k_lo),
    .r_v_i(1'b1),
    .r_tag_i(vtag_r),
    .r_match_o(tag_r_match_4k_lo)
  );


  bsg_cam_1r1w_replacement_00000008
  replacement_4k
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .read_v_i(tag_r_match_4k_lo),
    .alloc_v_i(fill_kilopage),
    .alloc_empty_i(tag_empty_4k_lo),
    .alloc_v_o(repl_way_4k_lo)
  );


  bsg_cam_1r1w_tag_array_0000001b_00000002
  tag_array_2m
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(tag_2m_w_v_li),
    .w_set_not_clear_i(_3_net_),
    .w_tag_i(vtag_i),
    .w_empty_o(tag_empty_2m_lo),
    .r_v_i(1'b1),
    .r_tag_i(vtag_r),
    .r_match_o(tag_r_match_2m_lo)
  );


  bsg_cam_1r1w_replacement_00000002
  replacement_2m
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .read_v_i(tag_r_match_2m_lo),
    .alloc_v_i(fill_megapage),
    .alloc_empty_i(tag_empty_2m_lo),
    .alloc_v_o(repl_way_2m_lo)
  );


  bsg_cam_1r1w_tag_array_0000001b_00000001
  tag_array_1g
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(tag_1g_w_v_li[0]),
    .w_set_not_clear_i(_5_net_),
    .w_tag_i(vtag_i),
    .w_empty_o(tag_empty_1g_lo[0]),
    .r_v_i(1'b1),
    .r_tag_i(vtag_r),
    .r_match_o(tag_r_match_1g_lo[0])
  );


  bsg_cam_1r1w_replacement_00000001
  replacement_1g
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .read_v_i(tag_r_match_1g_lo[0]),
    .alloc_v_i(fill_gigapage),
    .alloc_empty_i(tag_empty_1g_lo[0]),
    .alloc_v_o(repl_way_1g_lo[0])
  );


  bsg_dff_en_00000024
  \mem_array_4k_0_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted),
    .en_i(mem_4k_w_v_li[0]),
    .data_o({ data_4k_high_r[17:0], data_4k_med_r[8:0], data_4k_low_r[8:0] })
  );


  bsg_dff_en_00000024
  \mem_array_4k_1_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted),
    .en_i(mem_4k_w_v_li[1]),
    .data_o({ data_4k_high_r[35:18], data_4k_med_r[17:9], data_4k_low_r[17:9] })
  );


  bsg_dff_en_00000024
  \mem_array_4k_2_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted),
    .en_i(mem_4k_w_v_li[2]),
    .data_o({ data_4k_high_r[53:36], data_4k_med_r[26:18], data_4k_low_r[26:18] })
  );


  bsg_dff_en_00000024
  \mem_array_4k_3_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted),
    .en_i(mem_4k_w_v_li[3]),
    .data_o({ data_4k_high_r[71:54], data_4k_med_r[35:27], data_4k_low_r[35:27] })
  );


  bsg_dff_en_00000024
  \mem_array_4k_4_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted),
    .en_i(mem_4k_w_v_li[4]),
    .data_o({ data_4k_high_r[89:72], data_4k_med_r[44:36], data_4k_low_r[44:36] })
  );


  bsg_dff_en_00000024
  \mem_array_4k_5_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted),
    .en_i(mem_4k_w_v_li[5]),
    .data_o({ data_4k_high_r[107:90], data_4k_med_r[53:45], data_4k_low_r[53:45] })
  );


  bsg_dff_en_00000024
  \mem_array_4k_6_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted),
    .en_i(mem_4k_w_v_li[6]),
    .data_o({ data_4k_high_r[125:108], data_4k_med_r[62:54], data_4k_low_r[62:54] })
  );


  bsg_dff_en_00000024
  \mem_array_4k_7_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted),
    .en_i(mem_4k_w_v_li[7]),
    .data_o({ data_4k_high_r[143:126], data_4k_med_r[71:63], data_4k_low_r[71:63] })
  );


  bsg_dff_en_0000001b
  \genblk2.mem_array_2m_0_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted[35:9]),
    .en_i(mem_2m_w_v_li[0]),
    .data_o({ data_2m_high_r[17:0], data_2m_med_r[8:0] })
  );


  bsg_dff_en_0000001b
  \genblk2.mem_array_2m_1_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted[35:9]),
    .en_i(mem_2m_w_v_li[1]),
    .data_o({ data_2m_high_r[35:18], data_2m_med_r[17:9] })
  );


  bsg_dff_en_width_p18
  \genblk3.mem_array_1g_0_.mem_reg 
  (
    .clk_i(clk_i),
    .data_i(entry_shifted[35:18]),
    .en_i(mem_1g_w_v_li[0]),
    .data_o(data_1g_high_r)
  );


  bsg_mux_one_hot_9_00000009
  one_hot_sel_low
  (
    .data_i({ vtag_r[8:0], data_4k_low_r }),
    .sel_one_hot_i({ _21_net__8_, tag_r_match_4k_lo }),
    .data_o(r_entry[8:0])
  );


  bsg_mux_one_hot_9_0000000b
  one_hot_sel_med
  (
    .data_i({ vtag_r[17:9], data_2m_med_r, data_4k_med_r }),
    .sel_one_hot_i({ tag_r_match_1g_lo[0:0], tag_r_match_2m_lo, tag_r_match_4k_lo }),
    .data_o(r_entry[17:9])
  );


  bsg_mux_one_hot_18_0000000b
  one_hot_sel_high
  (
    .data_i({ data_1g_high_r, data_2m_high_r, data_4k_high_r }),
    .sel_one_hot_i({ tag_r_match_1g_lo[0:0], tag_r_match_2m_lo, tag_r_match_4k_lo }),
    .data_o(r_entry[35:18])
  );


  bsg_popcount_width_p3
  mpc
  (
    .i({ tag_r_match_1g_lo[0:0], any_match_2m_lo, any_match_4k_lo }),
    .o(match_cnt)
  );


  bsg_rotate_right_width_p36
  entry_unshift
  (
    .data_i(r_entry),
    .rot_i({ 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0 }),
    .o(entry_o)
  );

  assign N0 = ~match_cnt[0];
  assign N1 = N0 | match_cnt[1];
  assign v_o = ~N1;
  assign w_v_li = v_i & w_i;
  assign fill_gigapage = w_v_li & entry_i[7];
  assign fill_megapage = w_v_li & entry_i[6];
  assign fill_kilopage = N4 & N5;
  assign N4 = w_v_li & N3;
  assign N3 = ~fill_gigapage;
  assign N5 = ~fill_megapage;
  assign tag_4k_w_v_li[7] = N6 | flush_4k_li;
  assign N6 = fill_kilopage & repl_way_4k_lo[7];
  assign tag_4k_w_v_li[6] = N7 | flush_4k_li;
  assign N7 = fill_kilopage & repl_way_4k_lo[6];
  assign tag_4k_w_v_li[5] = N8 | flush_4k_li;
  assign N8 = fill_kilopage & repl_way_4k_lo[5];
  assign tag_4k_w_v_li[4] = N9 | flush_4k_li;
  assign N9 = fill_kilopage & repl_way_4k_lo[4];
  assign tag_4k_w_v_li[3] = N10 | flush_4k_li;
  assign N10 = fill_kilopage & repl_way_4k_lo[3];
  assign tag_4k_w_v_li[2] = N11 | flush_4k_li;
  assign N11 = fill_kilopage & repl_way_4k_lo[2];
  assign tag_4k_w_v_li[1] = N12 | flush_4k_li;
  assign N12 = fill_kilopage & repl_way_4k_lo[1];
  assign tag_4k_w_v_li[0] = N13 | flush_4k_li;
  assign N13 = fill_kilopage & repl_way_4k_lo[0];
  assign _1_net_ = ~flush_4k_li;
  assign any_match_4k_lo = N19 | tag_r_match_4k_lo[0];
  assign N19 = N18 | tag_r_match_4k_lo[1];
  assign N18 = N17 | tag_r_match_4k_lo[2];
  assign N17 = N16 | tag_r_match_4k_lo[3];
  assign N16 = N15 | tag_r_match_4k_lo[4];
  assign N15 = N14 | tag_r_match_4k_lo[5];
  assign N14 = tag_r_match_4k_lo[7] | tag_r_match_4k_lo[6];
  assign tag_2m_w_v_li[1] = N20 | flush_2m_li;
  assign N20 = fill_megapage & repl_way_2m_lo[1];
  assign tag_2m_w_v_li[0] = N21 | flush_2m_li;
  assign N21 = fill_megapage & repl_way_2m_lo[0];
  assign _3_net_ = ~flush_2m_li;
  assign any_match_2m_lo = tag_r_match_2m_lo[1] | tag_r_match_2m_lo[0];
  assign tag_1g_w_v_li[0] = N22 | fence_i;
  assign N22 = fill_gigapage & repl_way_1g_lo[0];
  assign _5_net_ = ~fence_i;
  assign mem_4k_w_v_li[7] = fill_kilopage & repl_way_4k_lo[7];
  assign mem_4k_w_v_li[6] = fill_kilopage & repl_way_4k_lo[6];
  assign mem_4k_w_v_li[5] = fill_kilopage & repl_way_4k_lo[5];
  assign mem_4k_w_v_li[4] = fill_kilopage & repl_way_4k_lo[4];
  assign mem_4k_w_v_li[3] = fill_kilopage & repl_way_4k_lo[3];
  assign mem_4k_w_v_li[2] = fill_kilopage & repl_way_4k_lo[2];
  assign mem_4k_w_v_li[1] = fill_kilopage & repl_way_4k_lo[1];
  assign mem_4k_w_v_li[0] = fill_kilopage & repl_way_4k_lo[0];
  assign mem_2m_w_v_li[1] = fill_megapage & repl_way_2m_lo[1];
  assign mem_2m_w_v_li[0] = fill_megapage & repl_way_2m_lo[0];
  assign mem_1g_w_v_li[0] = fill_gigapage & repl_way_1g_lo[0];
  assign _21_net__8_ = tag_r_match_1g_lo[0] | any_match_2m_lo;
  assign flush_4k_li = N24 | N25;
  assign N24 = fence_i | N23;
  assign N23 = tag_r_match_1g_lo[0] & any_match_4k_lo;
  assign N25 = any_match_2m_lo & any_match_4k_lo;
  assign flush_2m_li = fence_i | N26;
  assign N26 = tag_r_match_1g_lo[0] & any_match_2m_lo;

endmodule



module bsg_dff_en_width_p37_harden_p0_strength_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [36:0] data_i;
  output [36:0] data_o;
  input clk_i;
  input en_i;
  wire [36:0] data_o;
  reg data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,
  data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,
  data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,
  data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,
  data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,
  data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,
  data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,
  data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_bypass_width_p37
(
  clk_i,
  en_i,
  data_i,
  data_o
);

  input [36:0] data_i;
  output [36:0] data_o;
  input clk_i;
  input en_i;
  wire [36:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_en_width_p37_harden_p0_strength_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(en_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_dff_sync_read_width_p37_bypass_p1
(
  clk_i,
  reset_i,
  v_n_i,
  data_i,
  data_o
);

  input [36:0] data_i;
  output [36:0] data_o;
  input clk_i;
  input reset_i;
  input v_n_i;
  wire [36:0] data_o;
  wire v_r;

  bsg_dff_width_p1
  v_reg
  (
    .clk_i(clk_i),
    .data_i(v_n_i),
    .data_o(v_r)
  );


  bsg_dff_en_bypass_width_p37
  \bypass.data_reg 
  (
    .clk_i(clk_i),
    .en_i(v_r),
    .data_i(data_i),
    .data_o(data_o)
  );


endmodule



module bp_pma_00
(
  clk_i,
  reset_i,
  ptag_i,
  uncached_mode_i,
  nonspec_mode_i,
  uncached_o,
  nonidem_o,
  dram_o
);

  input [27:0] ptag_i;
  input clk_i;
  input reset_i;
  input uncached_mode_i;
  input nonspec_mode_i;
  output uncached_o;
  output nonidem_o;
  output dram_o;
  wire uncached_o,nonidem_o,dram_o,is_local_addr,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,
  N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;
  assign N0 = ptag_i[26] | ptag_i[27];
  assign N1 = ptag_i[25] | N0;
  assign N2 = ptag_i[24] | N1;
  assign N3 = ptag_i[23] | N2;
  assign N4 = ptag_i[22] | N3;
  assign N5 = ptag_i[21] | N4;
  assign N6 = ptag_i[20] | N5;
  assign is_local_addr = ~N14;
  assign N14 = N13 | ptag_i[19];
  assign N13 = N12 | ptag_i[20];
  assign N12 = N11 | ptag_i[21];
  assign N11 = N10 | ptag_i[22];
  assign N10 = N9 | ptag_i[23];
  assign N9 = N8 | ptag_i[24];
  assign N8 = N7 | ptag_i[25];
  assign N7 = ptag_i[27] | ptag_i[26];
  assign uncached_o = N16 | uncached_mode_i;
  assign N16 = N15 | is_local_addr;
  assign N15 = N6 | N5;
  assign nonidem_o = N19 | nonspec_mode_i;
  assign N19 = N18 | uncached_mode_i;
  assign N18 = N17 | is_local_addr;
  assign N17 = N6 | N5;
  assign dram_o = N22 & N23;
  assign N22 = N20 & N21;
  assign N20 = ~is_local_addr;
  assign N21 = ~N5;
  assign N23 = ~N6;

endmodule



module bp_mmu_00_00000008_00000002_00000001_0
(
  clk_i,
  reset_i,
  flush_i,
  fence_i,
  priv_mode_i,
  trans_en_i,
  sum_i,
  mxr_i,
  uncached_mode_i,
  nonspec_mode_i,
  hio_mask_i,
  w_v_i,
  w_vtag_i,
  w_entry_i,
  r_v_i,
  r_instr_i,
  r_load_i,
  r_store_i,
  r_eaddr_i,
  r_size_i,
  r_cbo_i,
  r_ptw_i,
  r_v_o,
  r_ptag_o,
  r_instr_miss_o,
  r_load_miss_o,
  r_store_miss_o,
  r_uncached_o,
  r_nonidem_o,
  r_dram_o,
  r_instr_access_fault_o,
  r_load_access_fault_o,
  r_store_access_fault_o,
  r_instr_misaligned_o,
  r_load_misaligned_o,
  r_store_misaligned_o,
  r_instr_page_fault_o,
  r_load_page_fault_o,
  r_store_page_fault_o
);

  input [1:0] priv_mode_i;
  input [6:0] hio_mask_i;
  input [26:0] w_vtag_i;
  input [35:0] w_entry_i;
  input [63:0] r_eaddr_i;
  input [1:0] r_size_i;
  output [27:0] r_ptag_o;
  input clk_i;
  input reset_i;
  input flush_i;
  input fence_i;
  input trans_en_i;
  input sum_i;
  input mxr_i;
  input uncached_mode_i;
  input nonspec_mode_i;
  input w_v_i;
  input r_v_i;
  input r_instr_i;
  input r_load_i;
  input r_store_i;
  input r_cbo_i;
  input r_ptw_i;
  output r_v_o;
  output r_instr_miss_o;
  output r_load_miss_o;
  output r_store_miss_o;
  output r_uncached_o;
  output r_nonidem_o;
  output r_dram_o;
  output r_instr_access_fault_o;
  output r_load_access_fault_o;
  output r_store_access_fault_o;
  output r_instr_misaligned_o;
  output r_load_misaligned_o;
  output r_store_misaligned_o;
  output r_instr_page_fault_o;
  output r_load_page_fault_o;
  output r_store_page_fault_o;
  wire [27:0] r_ptag_o;
  wire r_v_o,r_instr_miss_o,r_load_miss_o,r_store_miss_o,r_uncached_o,r_nonidem_o,
  r_dram_o,r_instr_access_fault_o,r_load_access_fault_o,r_store_access_fault_o,
  r_instr_misaligned_o,r_load_misaligned_o,r_store_misaligned_o,r_instr_page_fault_o,
  r_load_page_fault_o,r_store_page_fault_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,
  N13,N14,N15,N16,N17,N18,N19,N20,r_misaligned,N21,N22,N23,trans_li,trans_r,
  r_misaligned_r,r_instr_r,r_load_r,r_store_r,r_cbo_r,r_ptw_r,r_v_r,tlb_r_v_li,tlb_v_li,
  N24,N25,tlb_r_v_lo,tlb_r_v_r,passthrough_entry_ptag__27_,
  passthrough_entry_ptag__26_,passthrough_entry_ptag__25_,passthrough_entry_ptag__24_,
  passthrough_entry_ptag__23_,passthrough_entry_ptag__22_,passthrough_entry_ptag__21_,
  passthrough_entry_ptag__20_,passthrough_entry_ptag__19_,passthrough_entry_ptag__18_,
  passthrough_entry_ptag__17_,passthrough_entry_ptag__16_,passthrough_entry_ptag__15_,
  passthrough_entry_ptag__14_,passthrough_entry_ptag__13_,passthrough_entry_ptag__12_,
  passthrough_entry_ptag__11_,passthrough_entry_ptag__10_,passthrough_entry_ptag__9_,
  passthrough_entry_ptag__8_,passthrough_entry_ptag__7_,passthrough_entry_ptag__6_,
  passthrough_entry_ptag__5_,passthrough_entry_ptag__4_,passthrough_entry_ptag__3_,
  passthrough_entry_ptag__2_,passthrough_entry_ptag__1_,
  passthrough_entry_ptag__0_,tlb_entry_lo_d_,tlb_entry_lo_u_,tlb_entry_lo_x_,tlb_entry_lo_w_,
  tlb_entry_lo_r_,N26,tlb_v_lo,eaddr_fault_v,cached_fault_v,hio_fault_v,instr_access_fault_v,
  load_access_fault_v,store_access_fault_v,any_access_fault_v,instr_exe_page_fault_v,
  instr_priv_page_fault_v,data_priv_page_fault,data_read_page_fault,
  data_write_page_fault,instr_page_fault_v,load_page_fault_v,store_page_fault_v,any_page_fault_v,
  any_fault_v,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,
  N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,
  N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,
  N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,
  N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,
  N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134;
  wire [51:28] r_etag_r;
  wire [26:0] tlb_vtag_li;
  wire [35:0] tlb_r_entry_lo,tlb_r_entry_r;
  assign N11 = N9 & N10;
  assign N14 = r_size_i[1] | N13;
  assign N17 = N16 | r_size_i[0];
  assign N19 = r_size_i[1] & r_size_i[0];
  assign N20 = N16 & N13;

  bsg_dff_reset_en_width_p59
  read_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(r_v_i),
    .data_i({ trans_li, r_misaligned, r_instr_i, r_load_i, r_store_i, r_cbo_i, r_ptw_i, r_eaddr_i[63:12] }),
    .data_o({ trans_r, r_misaligned_r, r_instr_r, r_load_r, r_store_r, r_cbo_r, r_ptw_r, r_etag_r, passthrough_entry_ptag__27_, passthrough_entry_ptag__26_, passthrough_entry_ptag__25_, passthrough_entry_ptag__24_, passthrough_entry_ptag__23_, passthrough_entry_ptag__22_, passthrough_entry_ptag__21_, passthrough_entry_ptag__20_, passthrough_entry_ptag__19_, passthrough_entry_ptag__18_, passthrough_entry_ptag__17_, passthrough_entry_ptag__16_, passthrough_entry_ptag__15_, passthrough_entry_ptag__14_, passthrough_entry_ptag__13_, passthrough_entry_ptag__12_, passthrough_entry_ptag__11_, passthrough_entry_ptag__10_, passthrough_entry_ptag__9_, passthrough_entry_ptag__8_, passthrough_entry_ptag__7_, passthrough_entry_ptag__6_, passthrough_entry_ptag__5_, passthrough_entry_ptag__4_, passthrough_entry_ptag__3_, passthrough_entry_ptag__2_, passthrough_entry_ptag__1_, passthrough_entry_ptag__0_ })
  );


  bsg_dff_reset_set_clear_width_p1
  r_v_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .set_i(r_v_i),
    .clear_i(1'b1),
    .data_o(r_v_r)
  );


  bp_tlb_00_00000001_00000002_00000008
  tlb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .fence_i(fence_i),
    .v_i(tlb_v_li),
    .w_i(w_v_i),
    .vtag_i(tlb_vtag_li),
    .entry_i(w_entry_i),
    .v_o(tlb_r_v_lo),
    .entry_o(tlb_r_entry_lo)
  );


  bsg_dff_sync_read_width_p37_bypass_p1
  entry_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_n_i(tlb_r_v_li),
    .data_i({ tlb_r_v_lo, tlb_r_entry_lo }),
    .data_o({ tlb_r_v_r, tlb_r_entry_r })
  );


  bp_pma_00
  pma
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ptag_i(r_ptag_o),
    .uncached_mode_i(uncached_mode_i),
    .nonspec_mode_i(nonspec_mode_i),
    .uncached_o(r_uncached_o),
    .nonidem_o(r_nonidem_o),
    .dram_o(r_dram_o)
  );

  assign N27 = r_ptag_o[26] | r_ptag_o[27];
  assign N28 = r_ptag_o[25] | N27;
  assign N29 = r_ptag_o[24] | N28;
  assign N30 = r_ptag_o[23] | N29;
  assign N31 = r_ptag_o[22] | N30;
  assign N32 = r_ptag_o[21] | N31;
  assign N33 = ~priv_mode_i[0];
  assign N34 = N33 | priv_mode_i[1];
  assign N35 = ~N34;
  assign N36 = priv_mode_i[0] | priv_mode_i[1];
  assign N37 = ~N36;
  assign N23 = (N0)? r_eaddr_i[0] : 
               (N1)? N21 : 
               (N2)? N22 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = N15;
  assign N1 = N18;
  assign N2 = N19;
  assign N3 = N20;
  assign r_misaligned = (N4)? N23 : 
                        (N12)? 1'b0 : 1'b0;
  assign N4 = N11;
  assign tlb_vtag_li = (N5)? w_vtag_i : 
                       (N6)? r_eaddr_i[38:12] : 1'b0;
  assign N5 = N25;
  assign N6 = N24;
  assign { r_ptag_o, tlb_entry_lo_d_, tlb_entry_lo_u_, tlb_entry_lo_x_, tlb_entry_lo_w_, tlb_entry_lo_r_ } = (N7)? { tlb_r_entry_r[35:8], tlb_r_entry_r[4:0] } : 
                                                                                                             (N8)? { passthrough_entry_ptag__27_, passthrough_entry_ptag__26_, passthrough_entry_ptag__25_, passthrough_entry_ptag__24_, passthrough_entry_ptag__23_, passthrough_entry_ptag__22_, passthrough_entry_ptag__21_, passthrough_entry_ptag__20_, passthrough_entry_ptag__19_, passthrough_entry_ptag__18_, passthrough_entry_ptag__17_, passthrough_entry_ptag__16_, passthrough_entry_ptag__15_, passthrough_entry_ptag__14_, passthrough_entry_ptag__13_, passthrough_entry_ptag__12_, passthrough_entry_ptag__11_, passthrough_entry_ptag__10_, passthrough_entry_ptag__9_, passthrough_entry_ptag__8_, passthrough_entry_ptag__7_, passthrough_entry_ptag__6_, passthrough_entry_ptag__5_, passthrough_entry_ptag__4_, passthrough_entry_ptag__3_, passthrough_entry_ptag__2_, passthrough_entry_ptag__1_, passthrough_entry_ptag__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N7 = trans_r;
  assign N8 = N26;
  assign tlb_v_lo = (N7)? tlb_r_v_r : 
                    (N8)? r_v_r : 1'b0;
  assign N9 = ~r_ptw_i;
  assign N10 = ~r_cbo_i;
  assign N12 = ~N11;
  assign N13 = ~r_size_i[0];
  assign N15 = ~N14;
  assign N16 = ~r_size_i[1];
  assign N18 = ~N17;
  assign N21 = r_eaddr_i[1] | r_eaddr_i[0];
  assign N22 = N38 | r_eaddr_i[0];
  assign N38 = r_eaddr_i[2] | r_eaddr_i[1];
  assign trans_li = trans_en_i & N39;
  assign N39 = ~r_ptw_i;
  assign tlb_r_v_li = r_v_i | flush_i;
  assign tlb_v_li = tlb_r_v_li | w_v_i;
  assign N24 = ~w_v_i;
  assign N25 = w_v_i;
  assign N26 = ~trans_r;
  assign eaddr_fault_v = N65 & N90;
  assign N65 = ~N64;
  assign N64 = N63 & passthrough_entry_ptag__26_;
  assign N63 = N62 & passthrough_entry_ptag__27_;
  assign N62 = N61 & r_etag_r[28];
  assign N61 = N60 & r_etag_r[29];
  assign N60 = N59 & r_etag_r[30];
  assign N59 = N58 & r_etag_r[31];
  assign N58 = N57 & r_etag_r[32];
  assign N57 = N56 & r_etag_r[33];
  assign N56 = N55 & r_etag_r[34];
  assign N55 = N54 & r_etag_r[35];
  assign N54 = N53 & r_etag_r[36];
  assign N53 = N52 & r_etag_r[37];
  assign N52 = N51 & r_etag_r[38];
  assign N51 = N50 & r_etag_r[39];
  assign N50 = N49 & r_etag_r[40];
  assign N49 = N48 & r_etag_r[41];
  assign N48 = N47 & r_etag_r[42];
  assign N47 = N46 & r_etag_r[43];
  assign N46 = N45 & r_etag_r[44];
  assign N45 = N44 & r_etag_r[45];
  assign N44 = N43 & r_etag_r[46];
  assign N43 = N42 & r_etag_r[47];
  assign N42 = N41 & r_etag_r[48];
  assign N41 = N40 & r_etag_r[49];
  assign N40 = r_etag_r[51] & r_etag_r[50];
  assign N90 = N89 | passthrough_entry_ptag__26_;
  assign N89 = N88 | passthrough_entry_ptag__27_;
  assign N88 = N87 | r_etag_r[28];
  assign N87 = N86 | r_etag_r[29];
  assign N86 = N85 | r_etag_r[30];
  assign N85 = N84 | r_etag_r[31];
  assign N84 = N83 | r_etag_r[32];
  assign N83 = N82 | r_etag_r[33];
  assign N82 = N81 | r_etag_r[34];
  assign N81 = N80 | r_etag_r[35];
  assign N80 = N79 | r_etag_r[36];
  assign N79 = N78 | r_etag_r[37];
  assign N78 = N77 | r_etag_r[38];
  assign N77 = N76 | r_etag_r[39];
  assign N76 = N75 | r_etag_r[40];
  assign N75 = N74 | r_etag_r[41];
  assign N74 = N73 | r_etag_r[42];
  assign N73 = N72 | r_etag_r[43];
  assign N72 = N71 | r_etag_r[44];
  assign N71 = N70 | r_etag_r[45];
  assign N70 = N69 | r_etag_r[46];
  assign N69 = N68 | r_etag_r[47];
  assign N68 = N67 | r_etag_r[48];
  assign N67 = N66 | r_etag_r[49];
  assign N66 = r_etag_r[51] | r_etag_r[50];
  assign cached_fault_v = N91 & r_uncached_o;
  assign N91 = r_cbo_r & tlb_v_lo;
  assign hio_fault_v = N93 | N96;
  assign N93 = N92 & N32;
  assign N92 = r_instr_r & tlb_v_lo;
  assign N96 = N94 & N95;
  assign N94 = tlb_v_lo & r_ptag_o[21];
  assign N95 = ~hio_mask_i[0];
  assign instr_access_fault_v = r_instr_r & hio_fault_v;
  assign load_access_fault_v = r_load_r & cached_fault_v;
  assign store_access_fault_v = r_store_r & cached_fault_v;
  assign any_access_fault_v = N97 | store_access_fault_v;
  assign N97 = instr_access_fault_v | load_access_fault_v;
  assign instr_exe_page_fault_v = tlb_v_lo & N98;
  assign N98 = ~tlb_entry_lo_x_;
  assign instr_priv_page_fault_v = tlb_v_lo & N102;
  assign N102 = N99 | N101;
  assign N99 = N35 & tlb_entry_lo_u_;
  assign N101 = N37 & N100;
  assign N100 = ~tlb_entry_lo_u_;
  assign data_priv_page_fault = tlb_v_lo & N107;
  assign N107 = N105 | N106;
  assign N105 = N104 & tlb_entry_lo_u_;
  assign N104 = N35 & N103;
  assign N103 = ~sum_i;
  assign N106 = N37 & N100;
  assign data_read_page_fault = tlb_v_lo & N110;
  assign N110 = ~N109;
  assign N109 = tlb_entry_lo_r_ | N108;
  assign N108 = tlb_entry_lo_x_ & mxr_i;
  assign data_write_page_fault = tlb_v_lo & N112;
  assign N112 = ~N111;
  assign N111 = tlb_entry_lo_w_ & tlb_entry_lo_d_;
  assign instr_page_fault_v = N113 & N115;
  assign N113 = trans_r & r_instr_r;
  assign N115 = N114 | eaddr_fault_v;
  assign N114 = instr_priv_page_fault_v | instr_exe_page_fault_v;
  assign load_page_fault_v = N116 & N118;
  assign N116 = trans_r & r_load_r;
  assign N118 = N117 | eaddr_fault_v;
  assign N117 = data_priv_page_fault | data_read_page_fault;
  assign store_page_fault_v = N119 & N121;
  assign N119 = trans_r & r_store_r;
  assign N121 = N120 | eaddr_fault_v;
  assign N120 = data_priv_page_fault | data_write_page_fault;
  assign any_page_fault_v = N122 | store_page_fault_v;
  assign N122 = instr_page_fault_v | load_page_fault_v;
  assign any_fault_v = any_access_fault_v | any_page_fault_v;
  assign r_v_o = N123 & N124;
  assign N123 = r_v_r & tlb_v_lo;
  assign N124 = ~any_fault_v;
  assign r_instr_miss_o = N127 & r_instr_r;
  assign N127 = N126 & N124;
  assign N126 = r_v_r & N125;
  assign N125 = ~tlb_v_lo;
  assign r_load_miss_o = N129 & r_load_r;
  assign N129 = N128 & N124;
  assign N128 = r_v_r & N125;
  assign r_store_miss_o = N131 & r_store_r;
  assign N131 = N130 & N124;
  assign N130 = r_v_r & N125;
  assign r_instr_misaligned_o = N132 & r_instr_r;
  assign N132 = r_v_r & r_misaligned_r;
  assign r_load_misaligned_o = N133 & r_load_r;
  assign N133 = r_v_r & r_misaligned_r;
  assign r_store_misaligned_o = N134 & r_store_r;
  assign N134 = r_v_r & r_misaligned_r;
  assign r_instr_access_fault_o = r_v_r & instr_access_fault_v;
  assign r_load_access_fault_o = r_v_r & load_access_fault_v;
  assign r_store_access_fault_o = r_v_r & store_access_fault_v;
  assign r_instr_page_fault_o = r_v_r & instr_page_fault_v;
  assign r_load_page_fault_o = r_v_r & load_page_fault_v;
  assign r_store_page_fault_o = r_v_r & store_page_fault_v;

endmodule



module bp_be_dcache_decoder_00_00000ffe
(
  pkt_i,
  decode_o
);

  input [22:0] pkt_i;
  output [32:0] decode_o;
  wire [32:0] decode_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,decode_o_4_,decode_o_3_,
  decode_o_2_,decode_o_1_,decode_o_0_,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,
  N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,
  N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
  N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,
  N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,
  N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,
  N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,
  N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,
  N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,
  N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,
  N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,
  N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,
  N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,
  N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,
  N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,
  N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,
  N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,
  N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,
  N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,
  N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,
  N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,
  N362,N363,N364,N365,N366,N367,N368,N369,N371,N372,N373,N374,N375,N376,N377,N378,
  N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,
  N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,
  N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,
  N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,
  N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458;
  assign decode_o[17] = 1'b0;
  assign decode_o_4_ = pkt_i[22];
  assign decode_o[4] = decode_o_4_;
  assign decode_o_3_ = pkt_i[21];
  assign decode_o[3] = decode_o_3_;
  assign decode_o_2_ = pkt_i[20];
  assign decode_o[2] = decode_o_2_;
  assign decode_o_1_ = pkt_i[19];
  assign decode_o[1] = decode_o_1_;
  assign decode_o_0_ = pkt_i[18];
  assign decode_o[0] = decode_o_0_;
  assign N14 = N26 | N342;
  assign N15 = N105 | N14;
  assign N16 = ~N15;
  assign N17 = N105 | N23;
  assign N18 = ~N17;
  assign decode_o[16] = N16 | N18;
  assign N19 = ~pkt_i[14];
  assign N20 = pkt_i[16] | pkt_i[17];
  assign N21 = N255 | N20;
  assign N22 = N19 | N21;
  assign N23 = pkt_i[13] | N22;
  assign N24 = pkt_i[12] | N23;
  assign N25 = ~N24;
  assign N26 = ~pkt_i[13];
  assign N27 = N26 | N22;
  assign N28 = pkt_i[12] | N27;
  assign N29 = ~N28;
  assign decode_o[15] = N25 | N29;
  assign N30 = pkt_i[17] | pkt_i[16];
  assign N31 = N26 | N105;
  assign N32 = N30 | N278;
  assign N33 = N32 | N31;
  assign N34 = N30 | N261;
  assign N35 = N34 | N262;
  assign N37 = N34 | N273;
  assign N38 = N34 | N265;
  assign N40 = pkt_i[17] | N99;
  assign N41 = N40 | N272;
  assign N42 = N41 | N273;
  assign N43 = N255 | pkt_i[14];
  assign N44 = N40 | N43;
  assign N45 = N44 | N262;
  assign N47 = N41 | N262;
  assign N48 = N44 | N265;
  assign N50 = N41 | N265;
  assign N51 = N44 | N31;
  assign N53 = N41 | N31;
  assign N54 = N40 | N261;
  assign N55 = N54 | N273;
  assign N57 = N40 | N278;
  assign N58 = N57 | N273;
  assign N59 = N54 | N262;
  assign N61 = N57 | N262;
  assign N62 = N54 | N265;
  assign N64 = N57 | N265;
  assign N65 = N54 | N31;
  assign N67 = N57 | N31;
  assign N68 = N98 | pkt_i[16];
  assign N69 = N68 | N272;
  assign N70 = N69 | N273;
  assign N72 = N44 | N273;
  assign N73 = N69 | N262;
  assign N75 = N305 & N268;
  assign N76 = N99 & N255;
  assign N77 = N76 & N314;
  assign N78 = pkt_i[17] & pkt_i[13];
  assign N79 = pkt_i[13] & N105;
  assign N80 = N76 & N79;
  assign N81 = N329 & pkt_i[13];
  assign N82 = pkt_i[17] & pkt_i[14];
  assign N83 = pkt_i[14] & N105;
  assign N84 = N76 & N83;
  assign N85 = N305 & N19;
  assign N86 = N98 & N99;
  assign N87 = N86 & N19;
  assign N89 = N26 | N102;
  assign N90 = pkt_i[12] | N89;
  assign N91 = ~N90;
  assign decode_o[10] = N91 | N97;
  assign N92 = N105 | N103;
  assign N93 = ~N92;
  assign N94 = N19 | N101;
  assign N95 = pkt_i[13] | N94;
  assign N96 = pkt_i[12] | N95;
  assign N97 = ~N96;
  assign decode_o[11] = N93 | N97;
  assign N98 = ~pkt_i[17];
  assign N99 = ~pkt_i[16];
  assign N100 = N99 | N98;
  assign N101 = pkt_i[15] | N100;
  assign N102 = pkt_i[14] | N101;
  assign N103 = pkt_i[13] | N102;
  assign N104 = pkt_i[12] | N103;
  assign decode_o[9] = ~N104;
  assign N105 = ~pkt_i[12];
  assign N106 = pkt_i[13] | N109;
  assign N107 = N105 | N106;
  assign N108 = ~N107;
  assign decode_o[12] = N108 | N117;
  assign N109 = N19 | N256;
  assign N110 = N26 | N109;
  assign N111 = pkt_i[12] | N110;
  assign N112 = ~N111;
  assign N113 = pkt_i[16] & pkt_i[17];
  assign N114 = pkt_i[15] & N113;
  assign N115 = pkt_i[14] & N114;
  assign N116 = pkt_i[13] & N115;
  assign N117 = pkt_i[12] & N116;
  assign decode_o[13] = N112 | N117;
  assign N118 = N105 | N121;
  assign N119 = ~N118;
  assign N120 = N253 | N119;
  assign N121 = N26 | N128;
  assign N122 = pkt_i[12] | N121;
  assign N123 = ~N122;
  assign N124 = N120 | N123;
  assign N125 = N105 | N129;
  assign N126 = ~N125;
  assign N127 = N124 | N126;
  assign N128 = pkt_i[14] | N341;
  assign N129 = pkt_i[13] | N128;
  assign N130 = pkt_i[12] | N129;
  assign N131 = ~N130;
  assign N132 = N127 | N131;
  assign N133 = N132 | N337;
  assign N134 = N133 | N339;
  assign N135 = N134 | N345;
  assign N136 = ~N259;
  assign N137 = N135 | N136;
  assign N138 = N26 | N147;
  assign N139 = N105 | N138;
  assign N140 = ~N139;
  assign N141 = pkt_i[12] | N138;
  assign N142 = ~N141;
  assign N143 = N140 | N142;
  assign N144 = N105 | N148;
  assign N145 = ~N144;
  assign N146 = N143 | N145;
  assign N147 = pkt_i[14] | N21;
  assign N148 = pkt_i[13] | N147;
  assign N149 = pkt_i[12] | N148;
  assign N150 = ~N149;
  assign N151 = N146 | N150;
  assign N152 = pkt_i[12] | N158;
  assign N153 = ~N152;
  assign N154 = N151 | N153;
  assign N155 = pkt_i[16] | N98;
  assign N156 = pkt_i[15] | N155;
  assign N157 = N19 | N156;
  assign N158 = pkt_i[13] | N157;
  assign N159 = N105 | N158;
  assign N160 = ~N159;
  assign N161 = N154 | N160;
  assign N162 = ~N104;
  assign N163 = N161 | N162;
  assign N164 = N131 | N126;
  assign N165 = N164 | N123;
  assign N166 = N165 | N119;
  assign N167 = N166 | N345;
  assign N168 = N167 | N339;
  assign N169 = N168 | N337;
  assign N170 = N169 | N150;
  assign N171 = N170 | N145;
  assign N172 = N171 | N142;
  assign N173 = N172 | N140;
  assign N174 = N173 | N16;
  assign N175 = N174 | N25;
  assign N176 = N175 | N18;
  assign N177 = N176 | N29;
  assign N178 = pkt_i[12] | N181;
  assign N179 = ~N178;
  assign N180 = N177 | N179;
  assign N181 = pkt_i[13] | N188;
  assign N182 = N105 | N181;
  assign N183 = ~N182;
  assign N184 = N180 | N183;
  assign N185 = pkt_i[12] | N189;
  assign N186 = ~N185;
  assign N187 = N184 | N186;
  assign N188 = pkt_i[14] | N203;
  assign N189 = N26 | N188;
  assign N190 = N105 | N189;
  assign N191 = ~N190;
  assign N192 = N187 | N191;
  assign N193 = pkt_i[12] | N196;
  assign N194 = ~N193;
  assign N195 = N192 | N194;
  assign N196 = pkt_i[13] | N204;
  assign N197 = N105 | N196;
  assign N198 = ~N197;
  assign N199 = N195 | N198;
  assign N200 = pkt_i[12] | N205;
  assign N201 = ~N200;
  assign N202 = N199 | N201;
  assign N203 = pkt_i[15] | N234;
  assign N204 = N19 | N203;
  assign N205 = N26 | N204;
  assign N206 = N105 | N205;
  assign N207 = ~N206;
  assign N208 = N202 | N207;
  assign N209 = pkt_i[12] | N212;
  assign N210 = ~N209;
  assign N211 = N208 | N210;
  assign N212 = pkt_i[13] | N219;
  assign N213 = N105 | N212;
  assign N214 = ~N213;
  assign N215 = N211 | N214;
  assign N216 = pkt_i[12] | N220;
  assign N217 = ~N216;
  assign N218 = N215 | N217;
  assign N219 = pkt_i[14] | N235;
  assign N220 = N26 | N219;
  assign N221 = N105 | N220;
  assign N222 = ~N221;
  assign N223 = N218 | N222;
  assign N224 = pkt_i[12] | N227;
  assign N225 = ~N224;
  assign N226 = N223 | N225;
  assign N227 = pkt_i[13] | N236;
  assign N228 = N105 | N227;
  assign N229 = ~N228;
  assign N230 = N226 | N229;
  assign N231 = pkt_i[12] | N237;
  assign N232 = ~N231;
  assign N233 = N230 | N232;
  assign N234 = N99 | pkt_i[17];
  assign N235 = N255 | N234;
  assign N236 = N19 | N235;
  assign N237 = N26 | N236;
  assign N238 = N105 | N237;
  assign N239 = ~N238;
  assign N240 = N233 | N239;
  assign N241 = pkt_i[12] | N244;
  assign N242 = ~N241;
  assign N243 = N240 | N242;
  assign N244 = pkt_i[13] | N247;
  assign N245 = N105 | N244;
  assign N246 = ~N245;
  assign decode_o[25] = N243 | N246;
  assign N247 = pkt_i[14] | N156;
  assign N248 = N26 | N247;
  assign N249 = pkt_i[12] | N248;
  assign N250 = ~N249;
  assign N251 = N105 | N248;
  assign N252 = ~N251;
  assign N253 = N250 | N252;
  assign N254 = N253 | N153;
  assign decode_o[26] = N254 | N160;
  assign N255 = ~pkt_i[15];
  assign N256 = N255 | N100;
  assign N257 = pkt_i[14] | N256;
  assign N258 = pkt_i[13] | N257;
  assign N259 = pkt_i[12] | N258;
  assign decode_o[24] = ~N259;
  assign N260 = N98 | N99;
  assign N261 = N255 | N19;
  assign N262 = pkt_i[13] | N105;
  assign N263 = N260 | N261;
  assign N264 = N263 | N262;
  assign N265 = N26 | pkt_i[12];
  assign N266 = N263 | N265;
  assign N267 = pkt_i[17] & pkt_i[16];
  assign N268 = pkt_i[13] & pkt_i[12];
  assign N269 = N267 & N310;
  assign N270 = N269 & N268;
  assign N272 = pkt_i[15] | pkt_i[14];
  assign N273 = pkt_i[13] | pkt_i[12];
  assign N274 = N260 | N272;
  assign N275 = N274 | N273;
  assign N276 = N274 | N265;
  assign N277 = N274 | N262;
  assign N278 = pkt_i[15] | N19;
  assign N279 = N260 | N278;
  assign N280 = N279 | N273;
  assign N282 = N255 & N19;
  assign N283 = N26 & N105;
  assign N284 = N86 & N282;
  assign N285 = N284 & N283;
  assign N286 = N32 | N273;
  assign N287 = N296 | N273;
  assign N289 = N293 | N262;
  assign N290 = N32 | N262;
  assign N291 = N296 | N262;
  assign N293 = N30 | N272;
  assign N294 = N293 | N265;
  assign N295 = N32 | N265;
  assign N296 = N30 | N43;
  assign N297 = N296 | N265;
  assign N298 = N69 | N265;
  assign N299 = N68 | N278;
  assign N300 = N299 | N273;
  assign N302 = N98 & pkt_i[15];
  assign N303 = pkt_i[14] & pkt_i[12];
  assign N304 = N302 & N303;
  assign N305 = N99 & pkt_i[15];
  assign N306 = N305 & N303;
  assign N307 = pkt_i[17] & N255;
  assign N308 = N307 & N303;
  assign N309 = N98 & pkt_i[16];
  assign N310 = pkt_i[15] & pkt_i[14];
  assign N311 = N309 & N310;
  assign N312 = pkt_i[14] & pkt_i[13];
  assign N313 = N307 & N312;
  assign N314 = pkt_i[14] & N26;
  assign N315 = N322 & N314;
  assign N316 = N315 & N105;
  assign N317 = N320 & N312;
  assign N318 = N317 & N105;
  assign N319 = N305 & N312;
  assign N320 = pkt_i[17] & N99;
  assign N321 = N320 & pkt_i[15];
  assign N322 = pkt_i[16] & pkt_i[15];
  assign N323 = N19 & pkt_i[12];
  assign N324 = N322 & N323;
  assign N325 = pkt_i[17] & N19;
  assign N326 = N325 & N268;
  assign N327 = N19 & pkt_i[13];
  assign N328 = N322 & N327;
  assign N329 = N99 & N19;
  assign N330 = N329 & N268;
  assign N331 = pkt_i[17] & pkt_i[15];
  assign N332 = N331 & N19;
  assign N333 = N19 & N26;
  assign N334 = N320 & N333;
  assign N336 = pkt_i[12] | N14;
  assign N337 = ~N336;
  assign N338 = N105 | N343;
  assign N339 = ~N338;
  assign N340 = N337 | N339;
  assign N341 = pkt_i[15] | N20;
  assign N342 = N19 | N341;
  assign N343 = pkt_i[13] | N342;
  assign N344 = pkt_i[12] | N343;
  assign N345 = ~N344;
  assign N346 = N340 | N345;
  assign N364 = decode_o_3_ | decode_o_4_;
  assign N365 = decode_o_2_ | N364;
  assign N366 = decode_o_1_ | N365;
  assign N367 = decode_o_0_ | N366;
  assign N368 = decode_o[7] | decode_o[8];
  assign N369 = decode_o[6] | N368;
  assign decode_o[14] = decode_o[5] | N369;
  assign decode_o[8:5] = (N0)? { 1'b0, 1'b0, 1'b0, 1'b1 } : 
                         (N1)? { 1'b0, 1'b0, 1'b1, 1'b0 } : 
                         (N2)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                         (N3)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                         (N4)? { 1'b0, 1'b1, 1'b0, 1'b1 } : 
                         (N5)? { 1'b0, 1'b1, 1'b1, 1'b0 } : 
                         (N6)? { 1'b0, 1'b1, 1'b1, 1'b1 } : 
                         (N7)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                         (N8)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                         (N9)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                         (N10)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                         (N11)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N36;
  assign N1 = N39;
  assign N2 = N46;
  assign N3 = N49;
  assign N4 = N52;
  assign N5 = N56;
  assign N6 = N60;
  assign N7 = N63;
  assign N8 = N66;
  assign N9 = N71;
  assign N10 = N74;
  assign N11 = N88;
  assign decode_o[31] = (N12)? 1'b1 : 
                        (N357)? 1'b0 : 
                        (N360)? 1'b1 : 
                        (N363)? 1'b1 : 
                        (N354)? 1'b0 : 1'b0;
  assign N12 = N347;
  assign decode_o[32] = (N12)? 1'b1 : 
                        (N357)? 1'b1 : 
                        (N355)? 1'b0 : 
                        (N13)? 1'b0 : 
                        (N13)? 1'b0 : 1'b0;
  assign N13 = 1'b0;
  assign N36 = N371 | N372;
  assign N371 = ~N33;
  assign N372 = ~N35;
  assign N39 = N373 | N374;
  assign N373 = ~N37;
  assign N374 = ~N38;
  assign N46 = N375 | N376;
  assign N375 = ~N42;
  assign N376 = ~N45;
  assign N49 = N377 | N378;
  assign N377 = ~N47;
  assign N378 = ~N48;
  assign N52 = N379 | N380;
  assign N379 = ~N50;
  assign N380 = ~N51;
  assign N56 = N381 | N382;
  assign N381 = ~N53;
  assign N382 = ~N55;
  assign N60 = N383 | N384;
  assign N383 = ~N58;
  assign N384 = ~N59;
  assign N63 = N385 | N386;
  assign N385 = ~N61;
  assign N386 = ~N62;
  assign N66 = N387 | N388;
  assign N387 = ~N64;
  assign N388 = ~N65;
  assign N71 = N389 | N390;
  assign N389 = ~N67;
  assign N390 = ~N70;
  assign N74 = N391 | N392;
  assign N391 = ~N72;
  assign N392 = ~N73;
  assign N88 = N75 | N401;
  assign N401 = N77 | N400;
  assign N400 = N78 | N399;
  assign N399 = N80 | N398;
  assign N398 = N81 | N397;
  assign N397 = N82 | N396;
  assign N396 = N84 | N395;
  assign N395 = N331 | N394;
  assign N394 = N85 | N393;
  assign N393 = N267 | N87;
  assign decode_o[30] = N402 | N137;
  assign N402 = decode_o[14] | decode_o[16];
  assign decode_o[28] = N404 | N163;
  assign N404 = decode_o[14] & N403;
  assign N403 = ~decode_o[16];
  assign N271 = N407 | N270;
  assign N407 = N405 | N406;
  assign N405 = ~N264;
  assign N406 = ~N266;
  assign N281 = N412 | N413;
  assign N412 = N410 | N411;
  assign N410 = N408 | N409;
  assign N408 = ~N275;
  assign N409 = ~N276;
  assign N411 = ~N277;
  assign N413 = ~N280;
  assign N288 = N415 | N416;
  assign N415 = N285 | N414;
  assign N414 = ~N286;
  assign N416 = ~N287;
  assign N292 = N419 | N420;
  assign N419 = N417 | N418;
  assign N417 = ~N289;
  assign N418 = ~N290;
  assign N420 = ~N291;
  assign N301 = N439 | N373;
  assign N439 = N438 | N371;
  assign N438 = N436 | N437;
  assign N436 = N434 | N435;
  assign N434 = N432 | N433;
  assign N432 = N430 | N431;
  assign N430 = N428 | N429;
  assign N428 = N427 | N391;
  assign N427 = N426 | N389;
  assign N426 = N425 | N387;
  assign N425 = N424 | N385;
  assign N424 = N423 | N383;
  assign N423 = N422 | N381;
  assign N422 = N421 | N379;
  assign N421 = N375 | N377;
  assign N429 = ~N294;
  assign N431 = ~N295;
  assign N433 = ~N297;
  assign N435 = ~N298;
  assign N437 = ~N300;
  assign N335 = N304 | N452;
  assign N452 = N306 | N451;
  assign N451 = N308 | N450;
  assign N450 = N311 | N449;
  assign N449 = N313 | N448;
  assign N448 = N316 | N447;
  assign N447 = N318 | N446;
  assign N446 = N319 | N445;
  assign N445 = N321 | N444;
  assign N444 = N324 | N443;
  assign N443 = N326 | N442;
  assign N442 = N328 | N441;
  assign N441 = N330 | N440;
  assign N440 = N332 | N334;
  assign decode_o[23] = N271;
  assign decode_o[22] = N281;
  assign decode_o[18] = N288;
  assign decode_o[19] = N292;
  assign decode_o[20] = N301;
  assign decode_o[21] = N335;
  assign decode_o[27] = N454 & N455;
  assign N454 = N453 | decode_o[20];
  assign N453 = decode_o[18] | decode_o[19];
  assign N455 = ~N346;
  assign N347 = decode_o[25] & decode_o[18];
  assign N348 = decode_o[25] & decode_o[19];
  assign N349 = decode_o[25] & decode_o[20];
  assign N350 = decode_o[26] & decode_o[20];
  assign N351 = N348 | N347;
  assign N352 = N349 | N351;
  assign N353 = N350 | N352;
  assign N354 = ~N353;
  assign N355 = ~N351;
  assign decode_o[29] = decode_o[30] & N458;
  assign N458 = N456 | N457;
  assign N456 = decode_o[24] | decode_o[26];
  assign N457 = decode_o[25] & N367;
  assign N356 = ~N347;
  assign N357 = N348 & N356;
  assign N358 = ~N348;
  assign N359 = N356 & N358;
  assign N360 = N349 & N359;
  assign N361 = ~N349;
  assign N362 = N359 & N361;
  assign N363 = N350 & N362;

endmodule



module bsg_mem_1rw_sync_mask_write_bit_000000b8_00000040_1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [183:0] data_i;
  input [5:0] addr_i;
  input [183:0] w_mask_i;
  output [183:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [183:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  addr_i,
  data_i,
  write_mask_i,
  data_o
);

  input [8:0] addr_i;
  input [63:0] data_i;
  input [7:0] write_mask_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [63:0] data_o;

  bsg_mem_1rw_sync_mask_write_byte_synth
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .w_i(w_i),
    .addr_i(addr_i),
    .data_i(data_i),
    .write_mask_i(write_mask_i),
    .data_o(data_o)
  );


endmodule



module bsg_dff_reset_width_p1
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  wire [0:0] data_o;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_width_p45
(
  clk_i,
  data_i,
  data_o
);

  input [44:0] data_i;
  output [44:0] data_o;
  input clk_i;
  wire [44:0] data_o;
  reg data_o_44_sv2v_reg,data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,
  data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,
  data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,
  data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,
  data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,
  data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,
  data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,
  data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mux_000002aa_2
(
  data_i,
  sel_i,
  data_o
);

  input [1363:0] data_i;
  input [0:0] sel_i;
  output [681:0] data_o;
  wire [681:0] data_o;
  wire N0,N1;
  assign data_o[681] = (N1)? data_i[681] : 
                       (N0)? data_i[1363] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[680] = (N1)? data_i[680] : 
                       (N0)? data_i[1362] : 1'b0;
  assign data_o[679] = (N1)? data_i[679] : 
                       (N0)? data_i[1361] : 1'b0;
  assign data_o[678] = (N1)? data_i[678] : 
                       (N0)? data_i[1360] : 1'b0;
  assign data_o[677] = (N1)? data_i[677] : 
                       (N0)? data_i[1359] : 1'b0;
  assign data_o[676] = (N1)? data_i[676] : 
                       (N0)? data_i[1358] : 1'b0;
  assign data_o[675] = (N1)? data_i[675] : 
                       (N0)? data_i[1357] : 1'b0;
  assign data_o[674] = (N1)? data_i[674] : 
                       (N0)? data_i[1356] : 1'b0;
  assign data_o[673] = (N1)? data_i[673] : 
                       (N0)? data_i[1355] : 1'b0;
  assign data_o[672] = (N1)? data_i[672] : 
                       (N0)? data_i[1354] : 1'b0;
  assign data_o[671] = (N1)? data_i[671] : 
                       (N0)? data_i[1353] : 1'b0;
  assign data_o[670] = (N1)? data_i[670] : 
                       (N0)? data_i[1352] : 1'b0;
  assign data_o[669] = (N1)? data_i[669] : 
                       (N0)? data_i[1351] : 1'b0;
  assign data_o[668] = (N1)? data_i[668] : 
                       (N0)? data_i[1350] : 1'b0;
  assign data_o[667] = (N1)? data_i[667] : 
                       (N0)? data_i[1349] : 1'b0;
  assign data_o[666] = (N1)? data_i[666] : 
                       (N0)? data_i[1348] : 1'b0;
  assign data_o[665] = (N1)? data_i[665] : 
                       (N0)? data_i[1347] : 1'b0;
  assign data_o[664] = (N1)? data_i[664] : 
                       (N0)? data_i[1346] : 1'b0;
  assign data_o[663] = (N1)? data_i[663] : 
                       (N0)? data_i[1345] : 1'b0;
  assign data_o[662] = (N1)? data_i[662] : 
                       (N0)? data_i[1344] : 1'b0;
  assign data_o[661] = (N1)? data_i[661] : 
                       (N0)? data_i[1343] : 1'b0;
  assign data_o[660] = (N1)? data_i[660] : 
                       (N0)? data_i[1342] : 1'b0;
  assign data_o[659] = (N1)? data_i[659] : 
                       (N0)? data_i[1341] : 1'b0;
  assign data_o[658] = (N1)? data_i[658] : 
                       (N0)? data_i[1340] : 1'b0;
  assign data_o[657] = (N1)? data_i[657] : 
                       (N0)? data_i[1339] : 1'b0;
  assign data_o[656] = (N1)? data_i[656] : 
                       (N0)? data_i[1338] : 1'b0;
  assign data_o[655] = (N1)? data_i[655] : 
                       (N0)? data_i[1337] : 1'b0;
  assign data_o[654] = (N1)? data_i[654] : 
                       (N0)? data_i[1336] : 1'b0;
  assign data_o[653] = (N1)? data_i[653] : 
                       (N0)? data_i[1335] : 1'b0;
  assign data_o[652] = (N1)? data_i[652] : 
                       (N0)? data_i[1334] : 1'b0;
  assign data_o[651] = (N1)? data_i[651] : 
                       (N0)? data_i[1333] : 1'b0;
  assign data_o[650] = (N1)? data_i[650] : 
                       (N0)? data_i[1332] : 1'b0;
  assign data_o[649] = (N1)? data_i[649] : 
                       (N0)? data_i[1331] : 1'b0;
  assign data_o[648] = (N1)? data_i[648] : 
                       (N0)? data_i[1330] : 1'b0;
  assign data_o[647] = (N1)? data_i[647] : 
                       (N0)? data_i[1329] : 1'b0;
  assign data_o[646] = (N1)? data_i[646] : 
                       (N0)? data_i[1328] : 1'b0;
  assign data_o[645] = (N1)? data_i[645] : 
                       (N0)? data_i[1327] : 1'b0;
  assign data_o[644] = (N1)? data_i[644] : 
                       (N0)? data_i[1326] : 1'b0;
  assign data_o[643] = (N1)? data_i[643] : 
                       (N0)? data_i[1325] : 1'b0;
  assign data_o[642] = (N1)? data_i[642] : 
                       (N0)? data_i[1324] : 1'b0;
  assign data_o[641] = (N1)? data_i[641] : 
                       (N0)? data_i[1323] : 1'b0;
  assign data_o[640] = (N1)? data_i[640] : 
                       (N0)? data_i[1322] : 1'b0;
  assign data_o[639] = (N1)? data_i[639] : 
                       (N0)? data_i[1321] : 1'b0;
  assign data_o[638] = (N1)? data_i[638] : 
                       (N0)? data_i[1320] : 1'b0;
  assign data_o[637] = (N1)? data_i[637] : 
                       (N0)? data_i[1319] : 1'b0;
  assign data_o[636] = (N1)? data_i[636] : 
                       (N0)? data_i[1318] : 1'b0;
  assign data_o[635] = (N1)? data_i[635] : 
                       (N0)? data_i[1317] : 1'b0;
  assign data_o[634] = (N1)? data_i[634] : 
                       (N0)? data_i[1316] : 1'b0;
  assign data_o[633] = (N1)? data_i[633] : 
                       (N0)? data_i[1315] : 1'b0;
  assign data_o[632] = (N1)? data_i[632] : 
                       (N0)? data_i[1314] : 1'b0;
  assign data_o[631] = (N1)? data_i[631] : 
                       (N0)? data_i[1313] : 1'b0;
  assign data_o[630] = (N1)? data_i[630] : 
                       (N0)? data_i[1312] : 1'b0;
  assign data_o[629] = (N1)? data_i[629] : 
                       (N0)? data_i[1311] : 1'b0;
  assign data_o[628] = (N1)? data_i[628] : 
                       (N0)? data_i[1310] : 1'b0;
  assign data_o[627] = (N1)? data_i[627] : 
                       (N0)? data_i[1309] : 1'b0;
  assign data_o[626] = (N1)? data_i[626] : 
                       (N0)? data_i[1308] : 1'b0;
  assign data_o[625] = (N1)? data_i[625] : 
                       (N0)? data_i[1307] : 1'b0;
  assign data_o[624] = (N1)? data_i[624] : 
                       (N0)? data_i[1306] : 1'b0;
  assign data_o[623] = (N1)? data_i[623] : 
                       (N0)? data_i[1305] : 1'b0;
  assign data_o[622] = (N1)? data_i[622] : 
                       (N0)? data_i[1304] : 1'b0;
  assign data_o[621] = (N1)? data_i[621] : 
                       (N0)? data_i[1303] : 1'b0;
  assign data_o[620] = (N1)? data_i[620] : 
                       (N0)? data_i[1302] : 1'b0;
  assign data_o[619] = (N1)? data_i[619] : 
                       (N0)? data_i[1301] : 1'b0;
  assign data_o[618] = (N1)? data_i[618] : 
                       (N0)? data_i[1300] : 1'b0;
  assign data_o[617] = (N1)? data_i[617] : 
                       (N0)? data_i[1299] : 1'b0;
  assign data_o[616] = (N1)? data_i[616] : 
                       (N0)? data_i[1298] : 1'b0;
  assign data_o[615] = (N1)? data_i[615] : 
                       (N0)? data_i[1297] : 1'b0;
  assign data_o[614] = (N1)? data_i[614] : 
                       (N0)? data_i[1296] : 1'b0;
  assign data_o[613] = (N1)? data_i[613] : 
                       (N0)? data_i[1295] : 1'b0;
  assign data_o[612] = (N1)? data_i[612] : 
                       (N0)? data_i[1294] : 1'b0;
  assign data_o[611] = (N1)? data_i[611] : 
                       (N0)? data_i[1293] : 1'b0;
  assign data_o[610] = (N1)? data_i[610] : 
                       (N0)? data_i[1292] : 1'b0;
  assign data_o[609] = (N1)? data_i[609] : 
                       (N0)? data_i[1291] : 1'b0;
  assign data_o[608] = (N1)? data_i[608] : 
                       (N0)? data_i[1290] : 1'b0;
  assign data_o[607] = (N1)? data_i[607] : 
                       (N0)? data_i[1289] : 1'b0;
  assign data_o[606] = (N1)? data_i[606] : 
                       (N0)? data_i[1288] : 1'b0;
  assign data_o[605] = (N1)? data_i[605] : 
                       (N0)? data_i[1287] : 1'b0;
  assign data_o[604] = (N1)? data_i[604] : 
                       (N0)? data_i[1286] : 1'b0;
  assign data_o[603] = (N1)? data_i[603] : 
                       (N0)? data_i[1285] : 1'b0;
  assign data_o[602] = (N1)? data_i[602] : 
                       (N0)? data_i[1284] : 1'b0;
  assign data_o[601] = (N1)? data_i[601] : 
                       (N0)? data_i[1283] : 1'b0;
  assign data_o[600] = (N1)? data_i[600] : 
                       (N0)? data_i[1282] : 1'b0;
  assign data_o[599] = (N1)? data_i[599] : 
                       (N0)? data_i[1281] : 1'b0;
  assign data_o[598] = (N1)? data_i[598] : 
                       (N0)? data_i[1280] : 1'b0;
  assign data_o[597] = (N1)? data_i[597] : 
                       (N0)? data_i[1279] : 1'b0;
  assign data_o[596] = (N1)? data_i[596] : 
                       (N0)? data_i[1278] : 1'b0;
  assign data_o[595] = (N1)? data_i[595] : 
                       (N0)? data_i[1277] : 1'b0;
  assign data_o[594] = (N1)? data_i[594] : 
                       (N0)? data_i[1276] : 1'b0;
  assign data_o[593] = (N1)? data_i[593] : 
                       (N0)? data_i[1275] : 1'b0;
  assign data_o[592] = (N1)? data_i[592] : 
                       (N0)? data_i[1274] : 1'b0;
  assign data_o[591] = (N1)? data_i[591] : 
                       (N0)? data_i[1273] : 1'b0;
  assign data_o[590] = (N1)? data_i[590] : 
                       (N0)? data_i[1272] : 1'b0;
  assign data_o[589] = (N1)? data_i[589] : 
                       (N0)? data_i[1271] : 1'b0;
  assign data_o[588] = (N1)? data_i[588] : 
                       (N0)? data_i[1270] : 1'b0;
  assign data_o[587] = (N1)? data_i[587] : 
                       (N0)? data_i[1269] : 1'b0;
  assign data_o[586] = (N1)? data_i[586] : 
                       (N0)? data_i[1268] : 1'b0;
  assign data_o[585] = (N1)? data_i[585] : 
                       (N0)? data_i[1267] : 1'b0;
  assign data_o[584] = (N1)? data_i[584] : 
                       (N0)? data_i[1266] : 1'b0;
  assign data_o[583] = (N1)? data_i[583] : 
                       (N0)? data_i[1265] : 1'b0;
  assign data_o[582] = (N1)? data_i[582] : 
                       (N0)? data_i[1264] : 1'b0;
  assign data_o[581] = (N1)? data_i[581] : 
                       (N0)? data_i[1263] : 1'b0;
  assign data_o[580] = (N1)? data_i[580] : 
                       (N0)? data_i[1262] : 1'b0;
  assign data_o[579] = (N1)? data_i[579] : 
                       (N0)? data_i[1261] : 1'b0;
  assign data_o[578] = (N1)? data_i[578] : 
                       (N0)? data_i[1260] : 1'b0;
  assign data_o[577] = (N1)? data_i[577] : 
                       (N0)? data_i[1259] : 1'b0;
  assign data_o[576] = (N1)? data_i[576] : 
                       (N0)? data_i[1258] : 1'b0;
  assign data_o[575] = (N1)? data_i[575] : 
                       (N0)? data_i[1257] : 1'b0;
  assign data_o[574] = (N1)? data_i[574] : 
                       (N0)? data_i[1256] : 1'b0;
  assign data_o[573] = (N1)? data_i[573] : 
                       (N0)? data_i[1255] : 1'b0;
  assign data_o[572] = (N1)? data_i[572] : 
                       (N0)? data_i[1254] : 1'b0;
  assign data_o[571] = (N1)? data_i[571] : 
                       (N0)? data_i[1253] : 1'b0;
  assign data_o[570] = (N1)? data_i[570] : 
                       (N0)? data_i[1252] : 1'b0;
  assign data_o[569] = (N1)? data_i[569] : 
                       (N0)? data_i[1251] : 1'b0;
  assign data_o[568] = (N1)? data_i[568] : 
                       (N0)? data_i[1250] : 1'b0;
  assign data_o[567] = (N1)? data_i[567] : 
                       (N0)? data_i[1249] : 1'b0;
  assign data_o[566] = (N1)? data_i[566] : 
                       (N0)? data_i[1248] : 1'b0;
  assign data_o[565] = (N1)? data_i[565] : 
                       (N0)? data_i[1247] : 1'b0;
  assign data_o[564] = (N1)? data_i[564] : 
                       (N0)? data_i[1246] : 1'b0;
  assign data_o[563] = (N1)? data_i[563] : 
                       (N0)? data_i[1245] : 1'b0;
  assign data_o[562] = (N1)? data_i[562] : 
                       (N0)? data_i[1244] : 1'b0;
  assign data_o[561] = (N1)? data_i[561] : 
                       (N0)? data_i[1243] : 1'b0;
  assign data_o[560] = (N1)? data_i[560] : 
                       (N0)? data_i[1242] : 1'b0;
  assign data_o[559] = (N1)? data_i[559] : 
                       (N0)? data_i[1241] : 1'b0;
  assign data_o[558] = (N1)? data_i[558] : 
                       (N0)? data_i[1240] : 1'b0;
  assign data_o[557] = (N1)? data_i[557] : 
                       (N0)? data_i[1239] : 1'b0;
  assign data_o[556] = (N1)? data_i[556] : 
                       (N0)? data_i[1238] : 1'b0;
  assign data_o[555] = (N1)? data_i[555] : 
                       (N0)? data_i[1237] : 1'b0;
  assign data_o[554] = (N1)? data_i[554] : 
                       (N0)? data_i[1236] : 1'b0;
  assign data_o[553] = (N1)? data_i[553] : 
                       (N0)? data_i[1235] : 1'b0;
  assign data_o[552] = (N1)? data_i[552] : 
                       (N0)? data_i[1234] : 1'b0;
  assign data_o[551] = (N1)? data_i[551] : 
                       (N0)? data_i[1233] : 1'b0;
  assign data_o[550] = (N1)? data_i[550] : 
                       (N0)? data_i[1232] : 1'b0;
  assign data_o[549] = (N1)? data_i[549] : 
                       (N0)? data_i[1231] : 1'b0;
  assign data_o[548] = (N1)? data_i[548] : 
                       (N0)? data_i[1230] : 1'b0;
  assign data_o[547] = (N1)? data_i[547] : 
                       (N0)? data_i[1229] : 1'b0;
  assign data_o[546] = (N1)? data_i[546] : 
                       (N0)? data_i[1228] : 1'b0;
  assign data_o[545] = (N1)? data_i[545] : 
                       (N0)? data_i[1227] : 1'b0;
  assign data_o[544] = (N1)? data_i[544] : 
                       (N0)? data_i[1226] : 1'b0;
  assign data_o[543] = (N1)? data_i[543] : 
                       (N0)? data_i[1225] : 1'b0;
  assign data_o[542] = (N1)? data_i[542] : 
                       (N0)? data_i[1224] : 1'b0;
  assign data_o[541] = (N1)? data_i[541] : 
                       (N0)? data_i[1223] : 1'b0;
  assign data_o[540] = (N1)? data_i[540] : 
                       (N0)? data_i[1222] : 1'b0;
  assign data_o[539] = (N1)? data_i[539] : 
                       (N0)? data_i[1221] : 1'b0;
  assign data_o[538] = (N1)? data_i[538] : 
                       (N0)? data_i[1220] : 1'b0;
  assign data_o[537] = (N1)? data_i[537] : 
                       (N0)? data_i[1219] : 1'b0;
  assign data_o[536] = (N1)? data_i[536] : 
                       (N0)? data_i[1218] : 1'b0;
  assign data_o[535] = (N1)? data_i[535] : 
                       (N0)? data_i[1217] : 1'b0;
  assign data_o[534] = (N1)? data_i[534] : 
                       (N0)? data_i[1216] : 1'b0;
  assign data_o[533] = (N1)? data_i[533] : 
                       (N0)? data_i[1215] : 1'b0;
  assign data_o[532] = (N1)? data_i[532] : 
                       (N0)? data_i[1214] : 1'b0;
  assign data_o[531] = (N1)? data_i[531] : 
                       (N0)? data_i[1213] : 1'b0;
  assign data_o[530] = (N1)? data_i[530] : 
                       (N0)? data_i[1212] : 1'b0;
  assign data_o[529] = (N1)? data_i[529] : 
                       (N0)? data_i[1211] : 1'b0;
  assign data_o[528] = (N1)? data_i[528] : 
                       (N0)? data_i[1210] : 1'b0;
  assign data_o[527] = (N1)? data_i[527] : 
                       (N0)? data_i[1209] : 1'b0;
  assign data_o[526] = (N1)? data_i[526] : 
                       (N0)? data_i[1208] : 1'b0;
  assign data_o[525] = (N1)? data_i[525] : 
                       (N0)? data_i[1207] : 1'b0;
  assign data_o[524] = (N1)? data_i[524] : 
                       (N0)? data_i[1206] : 1'b0;
  assign data_o[523] = (N1)? data_i[523] : 
                       (N0)? data_i[1205] : 1'b0;
  assign data_o[522] = (N1)? data_i[522] : 
                       (N0)? data_i[1204] : 1'b0;
  assign data_o[521] = (N1)? data_i[521] : 
                       (N0)? data_i[1203] : 1'b0;
  assign data_o[520] = (N1)? data_i[520] : 
                       (N0)? data_i[1202] : 1'b0;
  assign data_o[519] = (N1)? data_i[519] : 
                       (N0)? data_i[1201] : 1'b0;
  assign data_o[518] = (N1)? data_i[518] : 
                       (N0)? data_i[1200] : 1'b0;
  assign data_o[517] = (N1)? data_i[517] : 
                       (N0)? data_i[1199] : 1'b0;
  assign data_o[516] = (N1)? data_i[516] : 
                       (N0)? data_i[1198] : 1'b0;
  assign data_o[515] = (N1)? data_i[515] : 
                       (N0)? data_i[1197] : 1'b0;
  assign data_o[514] = (N1)? data_i[514] : 
                       (N0)? data_i[1196] : 1'b0;
  assign data_o[513] = (N1)? data_i[513] : 
                       (N0)? data_i[1195] : 1'b0;
  assign data_o[512] = (N1)? data_i[512] : 
                       (N0)? data_i[1194] : 1'b0;
  assign data_o[511] = (N1)? data_i[511] : 
                       (N0)? data_i[1193] : 1'b0;
  assign data_o[510] = (N1)? data_i[510] : 
                       (N0)? data_i[1192] : 1'b0;
  assign data_o[509] = (N1)? data_i[509] : 
                       (N0)? data_i[1191] : 1'b0;
  assign data_o[508] = (N1)? data_i[508] : 
                       (N0)? data_i[1190] : 1'b0;
  assign data_o[507] = (N1)? data_i[507] : 
                       (N0)? data_i[1189] : 1'b0;
  assign data_o[506] = (N1)? data_i[506] : 
                       (N0)? data_i[1188] : 1'b0;
  assign data_o[505] = (N1)? data_i[505] : 
                       (N0)? data_i[1187] : 1'b0;
  assign data_o[504] = (N1)? data_i[504] : 
                       (N0)? data_i[1186] : 1'b0;
  assign data_o[503] = (N1)? data_i[503] : 
                       (N0)? data_i[1185] : 1'b0;
  assign data_o[502] = (N1)? data_i[502] : 
                       (N0)? data_i[1184] : 1'b0;
  assign data_o[501] = (N1)? data_i[501] : 
                       (N0)? data_i[1183] : 1'b0;
  assign data_o[500] = (N1)? data_i[500] : 
                       (N0)? data_i[1182] : 1'b0;
  assign data_o[499] = (N1)? data_i[499] : 
                       (N0)? data_i[1181] : 1'b0;
  assign data_o[498] = (N1)? data_i[498] : 
                       (N0)? data_i[1180] : 1'b0;
  assign data_o[497] = (N1)? data_i[497] : 
                       (N0)? data_i[1179] : 1'b0;
  assign data_o[496] = (N1)? data_i[496] : 
                       (N0)? data_i[1178] : 1'b0;
  assign data_o[495] = (N1)? data_i[495] : 
                       (N0)? data_i[1177] : 1'b0;
  assign data_o[494] = (N1)? data_i[494] : 
                       (N0)? data_i[1176] : 1'b0;
  assign data_o[493] = (N1)? data_i[493] : 
                       (N0)? data_i[1175] : 1'b0;
  assign data_o[492] = (N1)? data_i[492] : 
                       (N0)? data_i[1174] : 1'b0;
  assign data_o[491] = (N1)? data_i[491] : 
                       (N0)? data_i[1173] : 1'b0;
  assign data_o[490] = (N1)? data_i[490] : 
                       (N0)? data_i[1172] : 1'b0;
  assign data_o[489] = (N1)? data_i[489] : 
                       (N0)? data_i[1171] : 1'b0;
  assign data_o[488] = (N1)? data_i[488] : 
                       (N0)? data_i[1170] : 1'b0;
  assign data_o[487] = (N1)? data_i[487] : 
                       (N0)? data_i[1169] : 1'b0;
  assign data_o[486] = (N1)? data_i[486] : 
                       (N0)? data_i[1168] : 1'b0;
  assign data_o[485] = (N1)? data_i[485] : 
                       (N0)? data_i[1167] : 1'b0;
  assign data_o[484] = (N1)? data_i[484] : 
                       (N0)? data_i[1166] : 1'b0;
  assign data_o[483] = (N1)? data_i[483] : 
                       (N0)? data_i[1165] : 1'b0;
  assign data_o[482] = (N1)? data_i[482] : 
                       (N0)? data_i[1164] : 1'b0;
  assign data_o[481] = (N1)? data_i[481] : 
                       (N0)? data_i[1163] : 1'b0;
  assign data_o[480] = (N1)? data_i[480] : 
                       (N0)? data_i[1162] : 1'b0;
  assign data_o[479] = (N1)? data_i[479] : 
                       (N0)? data_i[1161] : 1'b0;
  assign data_o[478] = (N1)? data_i[478] : 
                       (N0)? data_i[1160] : 1'b0;
  assign data_o[477] = (N1)? data_i[477] : 
                       (N0)? data_i[1159] : 1'b0;
  assign data_o[476] = (N1)? data_i[476] : 
                       (N0)? data_i[1158] : 1'b0;
  assign data_o[475] = (N1)? data_i[475] : 
                       (N0)? data_i[1157] : 1'b0;
  assign data_o[474] = (N1)? data_i[474] : 
                       (N0)? data_i[1156] : 1'b0;
  assign data_o[473] = (N1)? data_i[473] : 
                       (N0)? data_i[1155] : 1'b0;
  assign data_o[472] = (N1)? data_i[472] : 
                       (N0)? data_i[1154] : 1'b0;
  assign data_o[471] = (N1)? data_i[471] : 
                       (N0)? data_i[1153] : 1'b0;
  assign data_o[470] = (N1)? data_i[470] : 
                       (N0)? data_i[1152] : 1'b0;
  assign data_o[469] = (N1)? data_i[469] : 
                       (N0)? data_i[1151] : 1'b0;
  assign data_o[468] = (N1)? data_i[468] : 
                       (N0)? data_i[1150] : 1'b0;
  assign data_o[467] = (N1)? data_i[467] : 
                       (N0)? data_i[1149] : 1'b0;
  assign data_o[466] = (N1)? data_i[466] : 
                       (N0)? data_i[1148] : 1'b0;
  assign data_o[465] = (N1)? data_i[465] : 
                       (N0)? data_i[1147] : 1'b0;
  assign data_o[464] = (N1)? data_i[464] : 
                       (N0)? data_i[1146] : 1'b0;
  assign data_o[463] = (N1)? data_i[463] : 
                       (N0)? data_i[1145] : 1'b0;
  assign data_o[462] = (N1)? data_i[462] : 
                       (N0)? data_i[1144] : 1'b0;
  assign data_o[461] = (N1)? data_i[461] : 
                       (N0)? data_i[1143] : 1'b0;
  assign data_o[460] = (N1)? data_i[460] : 
                       (N0)? data_i[1142] : 1'b0;
  assign data_o[459] = (N1)? data_i[459] : 
                       (N0)? data_i[1141] : 1'b0;
  assign data_o[458] = (N1)? data_i[458] : 
                       (N0)? data_i[1140] : 1'b0;
  assign data_o[457] = (N1)? data_i[457] : 
                       (N0)? data_i[1139] : 1'b0;
  assign data_o[456] = (N1)? data_i[456] : 
                       (N0)? data_i[1138] : 1'b0;
  assign data_o[455] = (N1)? data_i[455] : 
                       (N0)? data_i[1137] : 1'b0;
  assign data_o[454] = (N1)? data_i[454] : 
                       (N0)? data_i[1136] : 1'b0;
  assign data_o[453] = (N1)? data_i[453] : 
                       (N0)? data_i[1135] : 1'b0;
  assign data_o[452] = (N1)? data_i[452] : 
                       (N0)? data_i[1134] : 1'b0;
  assign data_o[451] = (N1)? data_i[451] : 
                       (N0)? data_i[1133] : 1'b0;
  assign data_o[450] = (N1)? data_i[450] : 
                       (N0)? data_i[1132] : 1'b0;
  assign data_o[449] = (N1)? data_i[449] : 
                       (N0)? data_i[1131] : 1'b0;
  assign data_o[448] = (N1)? data_i[448] : 
                       (N0)? data_i[1130] : 1'b0;
  assign data_o[447] = (N1)? data_i[447] : 
                       (N0)? data_i[1129] : 1'b0;
  assign data_o[446] = (N1)? data_i[446] : 
                       (N0)? data_i[1128] : 1'b0;
  assign data_o[445] = (N1)? data_i[445] : 
                       (N0)? data_i[1127] : 1'b0;
  assign data_o[444] = (N1)? data_i[444] : 
                       (N0)? data_i[1126] : 1'b0;
  assign data_o[443] = (N1)? data_i[443] : 
                       (N0)? data_i[1125] : 1'b0;
  assign data_o[442] = (N1)? data_i[442] : 
                       (N0)? data_i[1124] : 1'b0;
  assign data_o[441] = (N1)? data_i[441] : 
                       (N0)? data_i[1123] : 1'b0;
  assign data_o[440] = (N1)? data_i[440] : 
                       (N0)? data_i[1122] : 1'b0;
  assign data_o[439] = (N1)? data_i[439] : 
                       (N0)? data_i[1121] : 1'b0;
  assign data_o[438] = (N1)? data_i[438] : 
                       (N0)? data_i[1120] : 1'b0;
  assign data_o[437] = (N1)? data_i[437] : 
                       (N0)? data_i[1119] : 1'b0;
  assign data_o[436] = (N1)? data_i[436] : 
                       (N0)? data_i[1118] : 1'b0;
  assign data_o[435] = (N1)? data_i[435] : 
                       (N0)? data_i[1117] : 1'b0;
  assign data_o[434] = (N1)? data_i[434] : 
                       (N0)? data_i[1116] : 1'b0;
  assign data_o[433] = (N1)? data_i[433] : 
                       (N0)? data_i[1115] : 1'b0;
  assign data_o[432] = (N1)? data_i[432] : 
                       (N0)? data_i[1114] : 1'b0;
  assign data_o[431] = (N1)? data_i[431] : 
                       (N0)? data_i[1113] : 1'b0;
  assign data_o[430] = (N1)? data_i[430] : 
                       (N0)? data_i[1112] : 1'b0;
  assign data_o[429] = (N1)? data_i[429] : 
                       (N0)? data_i[1111] : 1'b0;
  assign data_o[428] = (N1)? data_i[428] : 
                       (N0)? data_i[1110] : 1'b0;
  assign data_o[427] = (N1)? data_i[427] : 
                       (N0)? data_i[1109] : 1'b0;
  assign data_o[426] = (N1)? data_i[426] : 
                       (N0)? data_i[1108] : 1'b0;
  assign data_o[425] = (N1)? data_i[425] : 
                       (N0)? data_i[1107] : 1'b0;
  assign data_o[424] = (N1)? data_i[424] : 
                       (N0)? data_i[1106] : 1'b0;
  assign data_o[423] = (N1)? data_i[423] : 
                       (N0)? data_i[1105] : 1'b0;
  assign data_o[422] = (N1)? data_i[422] : 
                       (N0)? data_i[1104] : 1'b0;
  assign data_o[421] = (N1)? data_i[421] : 
                       (N0)? data_i[1103] : 1'b0;
  assign data_o[420] = (N1)? data_i[420] : 
                       (N0)? data_i[1102] : 1'b0;
  assign data_o[419] = (N1)? data_i[419] : 
                       (N0)? data_i[1101] : 1'b0;
  assign data_o[418] = (N1)? data_i[418] : 
                       (N0)? data_i[1100] : 1'b0;
  assign data_o[417] = (N1)? data_i[417] : 
                       (N0)? data_i[1099] : 1'b0;
  assign data_o[416] = (N1)? data_i[416] : 
                       (N0)? data_i[1098] : 1'b0;
  assign data_o[415] = (N1)? data_i[415] : 
                       (N0)? data_i[1097] : 1'b0;
  assign data_o[414] = (N1)? data_i[414] : 
                       (N0)? data_i[1096] : 1'b0;
  assign data_o[413] = (N1)? data_i[413] : 
                       (N0)? data_i[1095] : 1'b0;
  assign data_o[412] = (N1)? data_i[412] : 
                       (N0)? data_i[1094] : 1'b0;
  assign data_o[411] = (N1)? data_i[411] : 
                       (N0)? data_i[1093] : 1'b0;
  assign data_o[410] = (N1)? data_i[410] : 
                       (N0)? data_i[1092] : 1'b0;
  assign data_o[409] = (N1)? data_i[409] : 
                       (N0)? data_i[1091] : 1'b0;
  assign data_o[408] = (N1)? data_i[408] : 
                       (N0)? data_i[1090] : 1'b0;
  assign data_o[407] = (N1)? data_i[407] : 
                       (N0)? data_i[1089] : 1'b0;
  assign data_o[406] = (N1)? data_i[406] : 
                       (N0)? data_i[1088] : 1'b0;
  assign data_o[405] = (N1)? data_i[405] : 
                       (N0)? data_i[1087] : 1'b0;
  assign data_o[404] = (N1)? data_i[404] : 
                       (N0)? data_i[1086] : 1'b0;
  assign data_o[403] = (N1)? data_i[403] : 
                       (N0)? data_i[1085] : 1'b0;
  assign data_o[402] = (N1)? data_i[402] : 
                       (N0)? data_i[1084] : 1'b0;
  assign data_o[401] = (N1)? data_i[401] : 
                       (N0)? data_i[1083] : 1'b0;
  assign data_o[400] = (N1)? data_i[400] : 
                       (N0)? data_i[1082] : 1'b0;
  assign data_o[399] = (N1)? data_i[399] : 
                       (N0)? data_i[1081] : 1'b0;
  assign data_o[398] = (N1)? data_i[398] : 
                       (N0)? data_i[1080] : 1'b0;
  assign data_o[397] = (N1)? data_i[397] : 
                       (N0)? data_i[1079] : 1'b0;
  assign data_o[396] = (N1)? data_i[396] : 
                       (N0)? data_i[1078] : 1'b0;
  assign data_o[395] = (N1)? data_i[395] : 
                       (N0)? data_i[1077] : 1'b0;
  assign data_o[394] = (N1)? data_i[394] : 
                       (N0)? data_i[1076] : 1'b0;
  assign data_o[393] = (N1)? data_i[393] : 
                       (N0)? data_i[1075] : 1'b0;
  assign data_o[392] = (N1)? data_i[392] : 
                       (N0)? data_i[1074] : 1'b0;
  assign data_o[391] = (N1)? data_i[391] : 
                       (N0)? data_i[1073] : 1'b0;
  assign data_o[390] = (N1)? data_i[390] : 
                       (N0)? data_i[1072] : 1'b0;
  assign data_o[389] = (N1)? data_i[389] : 
                       (N0)? data_i[1071] : 1'b0;
  assign data_o[388] = (N1)? data_i[388] : 
                       (N0)? data_i[1070] : 1'b0;
  assign data_o[387] = (N1)? data_i[387] : 
                       (N0)? data_i[1069] : 1'b0;
  assign data_o[386] = (N1)? data_i[386] : 
                       (N0)? data_i[1068] : 1'b0;
  assign data_o[385] = (N1)? data_i[385] : 
                       (N0)? data_i[1067] : 1'b0;
  assign data_o[384] = (N1)? data_i[384] : 
                       (N0)? data_i[1066] : 1'b0;
  assign data_o[383] = (N1)? data_i[383] : 
                       (N0)? data_i[1065] : 1'b0;
  assign data_o[382] = (N1)? data_i[382] : 
                       (N0)? data_i[1064] : 1'b0;
  assign data_o[381] = (N1)? data_i[381] : 
                       (N0)? data_i[1063] : 1'b0;
  assign data_o[380] = (N1)? data_i[380] : 
                       (N0)? data_i[1062] : 1'b0;
  assign data_o[379] = (N1)? data_i[379] : 
                       (N0)? data_i[1061] : 1'b0;
  assign data_o[378] = (N1)? data_i[378] : 
                       (N0)? data_i[1060] : 1'b0;
  assign data_o[377] = (N1)? data_i[377] : 
                       (N0)? data_i[1059] : 1'b0;
  assign data_o[376] = (N1)? data_i[376] : 
                       (N0)? data_i[1058] : 1'b0;
  assign data_o[375] = (N1)? data_i[375] : 
                       (N0)? data_i[1057] : 1'b0;
  assign data_o[374] = (N1)? data_i[374] : 
                       (N0)? data_i[1056] : 1'b0;
  assign data_o[373] = (N1)? data_i[373] : 
                       (N0)? data_i[1055] : 1'b0;
  assign data_o[372] = (N1)? data_i[372] : 
                       (N0)? data_i[1054] : 1'b0;
  assign data_o[371] = (N1)? data_i[371] : 
                       (N0)? data_i[1053] : 1'b0;
  assign data_o[370] = (N1)? data_i[370] : 
                       (N0)? data_i[1052] : 1'b0;
  assign data_o[369] = (N1)? data_i[369] : 
                       (N0)? data_i[1051] : 1'b0;
  assign data_o[368] = (N1)? data_i[368] : 
                       (N0)? data_i[1050] : 1'b0;
  assign data_o[367] = (N1)? data_i[367] : 
                       (N0)? data_i[1049] : 1'b0;
  assign data_o[366] = (N1)? data_i[366] : 
                       (N0)? data_i[1048] : 1'b0;
  assign data_o[365] = (N1)? data_i[365] : 
                       (N0)? data_i[1047] : 1'b0;
  assign data_o[364] = (N1)? data_i[364] : 
                       (N0)? data_i[1046] : 1'b0;
  assign data_o[363] = (N1)? data_i[363] : 
                       (N0)? data_i[1045] : 1'b0;
  assign data_o[362] = (N1)? data_i[362] : 
                       (N0)? data_i[1044] : 1'b0;
  assign data_o[361] = (N1)? data_i[361] : 
                       (N0)? data_i[1043] : 1'b0;
  assign data_o[360] = (N1)? data_i[360] : 
                       (N0)? data_i[1042] : 1'b0;
  assign data_o[359] = (N1)? data_i[359] : 
                       (N0)? data_i[1041] : 1'b0;
  assign data_o[358] = (N1)? data_i[358] : 
                       (N0)? data_i[1040] : 1'b0;
  assign data_o[357] = (N1)? data_i[357] : 
                       (N0)? data_i[1039] : 1'b0;
  assign data_o[356] = (N1)? data_i[356] : 
                       (N0)? data_i[1038] : 1'b0;
  assign data_o[355] = (N1)? data_i[355] : 
                       (N0)? data_i[1037] : 1'b0;
  assign data_o[354] = (N1)? data_i[354] : 
                       (N0)? data_i[1036] : 1'b0;
  assign data_o[353] = (N1)? data_i[353] : 
                       (N0)? data_i[1035] : 1'b0;
  assign data_o[352] = (N1)? data_i[352] : 
                       (N0)? data_i[1034] : 1'b0;
  assign data_o[351] = (N1)? data_i[351] : 
                       (N0)? data_i[1033] : 1'b0;
  assign data_o[350] = (N1)? data_i[350] : 
                       (N0)? data_i[1032] : 1'b0;
  assign data_o[349] = (N1)? data_i[349] : 
                       (N0)? data_i[1031] : 1'b0;
  assign data_o[348] = (N1)? data_i[348] : 
                       (N0)? data_i[1030] : 1'b0;
  assign data_o[347] = (N1)? data_i[347] : 
                       (N0)? data_i[1029] : 1'b0;
  assign data_o[346] = (N1)? data_i[346] : 
                       (N0)? data_i[1028] : 1'b0;
  assign data_o[345] = (N1)? data_i[345] : 
                       (N0)? data_i[1027] : 1'b0;
  assign data_o[344] = (N1)? data_i[344] : 
                       (N0)? data_i[1026] : 1'b0;
  assign data_o[343] = (N1)? data_i[343] : 
                       (N0)? data_i[1025] : 1'b0;
  assign data_o[342] = (N1)? data_i[342] : 
                       (N0)? data_i[1024] : 1'b0;
  assign data_o[341] = (N1)? data_i[341] : 
                       (N0)? data_i[1023] : 1'b0;
  assign data_o[340] = (N1)? data_i[340] : 
                       (N0)? data_i[1022] : 1'b0;
  assign data_o[339] = (N1)? data_i[339] : 
                       (N0)? data_i[1021] : 1'b0;
  assign data_o[338] = (N1)? data_i[338] : 
                       (N0)? data_i[1020] : 1'b0;
  assign data_o[337] = (N1)? data_i[337] : 
                       (N0)? data_i[1019] : 1'b0;
  assign data_o[336] = (N1)? data_i[336] : 
                       (N0)? data_i[1018] : 1'b0;
  assign data_o[335] = (N1)? data_i[335] : 
                       (N0)? data_i[1017] : 1'b0;
  assign data_o[334] = (N1)? data_i[334] : 
                       (N0)? data_i[1016] : 1'b0;
  assign data_o[333] = (N1)? data_i[333] : 
                       (N0)? data_i[1015] : 1'b0;
  assign data_o[332] = (N1)? data_i[332] : 
                       (N0)? data_i[1014] : 1'b0;
  assign data_o[331] = (N1)? data_i[331] : 
                       (N0)? data_i[1013] : 1'b0;
  assign data_o[330] = (N1)? data_i[330] : 
                       (N0)? data_i[1012] : 1'b0;
  assign data_o[329] = (N1)? data_i[329] : 
                       (N0)? data_i[1011] : 1'b0;
  assign data_o[328] = (N1)? data_i[328] : 
                       (N0)? data_i[1010] : 1'b0;
  assign data_o[327] = (N1)? data_i[327] : 
                       (N0)? data_i[1009] : 1'b0;
  assign data_o[326] = (N1)? data_i[326] : 
                       (N0)? data_i[1008] : 1'b0;
  assign data_o[325] = (N1)? data_i[325] : 
                       (N0)? data_i[1007] : 1'b0;
  assign data_o[324] = (N1)? data_i[324] : 
                       (N0)? data_i[1006] : 1'b0;
  assign data_o[323] = (N1)? data_i[323] : 
                       (N0)? data_i[1005] : 1'b0;
  assign data_o[322] = (N1)? data_i[322] : 
                       (N0)? data_i[1004] : 1'b0;
  assign data_o[321] = (N1)? data_i[321] : 
                       (N0)? data_i[1003] : 1'b0;
  assign data_o[320] = (N1)? data_i[320] : 
                       (N0)? data_i[1002] : 1'b0;
  assign data_o[319] = (N1)? data_i[319] : 
                       (N0)? data_i[1001] : 1'b0;
  assign data_o[318] = (N1)? data_i[318] : 
                       (N0)? data_i[1000] : 1'b0;
  assign data_o[317] = (N1)? data_i[317] : 
                       (N0)? data_i[999] : 1'b0;
  assign data_o[316] = (N1)? data_i[316] : 
                       (N0)? data_i[998] : 1'b0;
  assign data_o[315] = (N1)? data_i[315] : 
                       (N0)? data_i[997] : 1'b0;
  assign data_o[314] = (N1)? data_i[314] : 
                       (N0)? data_i[996] : 1'b0;
  assign data_o[313] = (N1)? data_i[313] : 
                       (N0)? data_i[995] : 1'b0;
  assign data_o[312] = (N1)? data_i[312] : 
                       (N0)? data_i[994] : 1'b0;
  assign data_o[311] = (N1)? data_i[311] : 
                       (N0)? data_i[993] : 1'b0;
  assign data_o[310] = (N1)? data_i[310] : 
                       (N0)? data_i[992] : 1'b0;
  assign data_o[309] = (N1)? data_i[309] : 
                       (N0)? data_i[991] : 1'b0;
  assign data_o[308] = (N1)? data_i[308] : 
                       (N0)? data_i[990] : 1'b0;
  assign data_o[307] = (N1)? data_i[307] : 
                       (N0)? data_i[989] : 1'b0;
  assign data_o[306] = (N1)? data_i[306] : 
                       (N0)? data_i[988] : 1'b0;
  assign data_o[305] = (N1)? data_i[305] : 
                       (N0)? data_i[987] : 1'b0;
  assign data_o[304] = (N1)? data_i[304] : 
                       (N0)? data_i[986] : 1'b0;
  assign data_o[303] = (N1)? data_i[303] : 
                       (N0)? data_i[985] : 1'b0;
  assign data_o[302] = (N1)? data_i[302] : 
                       (N0)? data_i[984] : 1'b0;
  assign data_o[301] = (N1)? data_i[301] : 
                       (N0)? data_i[983] : 1'b0;
  assign data_o[300] = (N1)? data_i[300] : 
                       (N0)? data_i[982] : 1'b0;
  assign data_o[299] = (N1)? data_i[299] : 
                       (N0)? data_i[981] : 1'b0;
  assign data_o[298] = (N1)? data_i[298] : 
                       (N0)? data_i[980] : 1'b0;
  assign data_o[297] = (N1)? data_i[297] : 
                       (N0)? data_i[979] : 1'b0;
  assign data_o[296] = (N1)? data_i[296] : 
                       (N0)? data_i[978] : 1'b0;
  assign data_o[295] = (N1)? data_i[295] : 
                       (N0)? data_i[977] : 1'b0;
  assign data_o[294] = (N1)? data_i[294] : 
                       (N0)? data_i[976] : 1'b0;
  assign data_o[293] = (N1)? data_i[293] : 
                       (N0)? data_i[975] : 1'b0;
  assign data_o[292] = (N1)? data_i[292] : 
                       (N0)? data_i[974] : 1'b0;
  assign data_o[291] = (N1)? data_i[291] : 
                       (N0)? data_i[973] : 1'b0;
  assign data_o[290] = (N1)? data_i[290] : 
                       (N0)? data_i[972] : 1'b0;
  assign data_o[289] = (N1)? data_i[289] : 
                       (N0)? data_i[971] : 1'b0;
  assign data_o[288] = (N1)? data_i[288] : 
                       (N0)? data_i[970] : 1'b0;
  assign data_o[287] = (N1)? data_i[287] : 
                       (N0)? data_i[969] : 1'b0;
  assign data_o[286] = (N1)? data_i[286] : 
                       (N0)? data_i[968] : 1'b0;
  assign data_o[285] = (N1)? data_i[285] : 
                       (N0)? data_i[967] : 1'b0;
  assign data_o[284] = (N1)? data_i[284] : 
                       (N0)? data_i[966] : 1'b0;
  assign data_o[283] = (N1)? data_i[283] : 
                       (N0)? data_i[965] : 1'b0;
  assign data_o[282] = (N1)? data_i[282] : 
                       (N0)? data_i[964] : 1'b0;
  assign data_o[281] = (N1)? data_i[281] : 
                       (N0)? data_i[963] : 1'b0;
  assign data_o[280] = (N1)? data_i[280] : 
                       (N0)? data_i[962] : 1'b0;
  assign data_o[279] = (N1)? data_i[279] : 
                       (N0)? data_i[961] : 1'b0;
  assign data_o[278] = (N1)? data_i[278] : 
                       (N0)? data_i[960] : 1'b0;
  assign data_o[277] = (N1)? data_i[277] : 
                       (N0)? data_i[959] : 1'b0;
  assign data_o[276] = (N1)? data_i[276] : 
                       (N0)? data_i[958] : 1'b0;
  assign data_o[275] = (N1)? data_i[275] : 
                       (N0)? data_i[957] : 1'b0;
  assign data_o[274] = (N1)? data_i[274] : 
                       (N0)? data_i[956] : 1'b0;
  assign data_o[273] = (N1)? data_i[273] : 
                       (N0)? data_i[955] : 1'b0;
  assign data_o[272] = (N1)? data_i[272] : 
                       (N0)? data_i[954] : 1'b0;
  assign data_o[271] = (N1)? data_i[271] : 
                       (N0)? data_i[953] : 1'b0;
  assign data_o[270] = (N1)? data_i[270] : 
                       (N0)? data_i[952] : 1'b0;
  assign data_o[269] = (N1)? data_i[269] : 
                       (N0)? data_i[951] : 1'b0;
  assign data_o[268] = (N1)? data_i[268] : 
                       (N0)? data_i[950] : 1'b0;
  assign data_o[267] = (N1)? data_i[267] : 
                       (N0)? data_i[949] : 1'b0;
  assign data_o[266] = (N1)? data_i[266] : 
                       (N0)? data_i[948] : 1'b0;
  assign data_o[265] = (N1)? data_i[265] : 
                       (N0)? data_i[947] : 1'b0;
  assign data_o[264] = (N1)? data_i[264] : 
                       (N0)? data_i[946] : 1'b0;
  assign data_o[263] = (N1)? data_i[263] : 
                       (N0)? data_i[945] : 1'b0;
  assign data_o[262] = (N1)? data_i[262] : 
                       (N0)? data_i[944] : 1'b0;
  assign data_o[261] = (N1)? data_i[261] : 
                       (N0)? data_i[943] : 1'b0;
  assign data_o[260] = (N1)? data_i[260] : 
                       (N0)? data_i[942] : 1'b0;
  assign data_o[259] = (N1)? data_i[259] : 
                       (N0)? data_i[941] : 1'b0;
  assign data_o[258] = (N1)? data_i[258] : 
                       (N0)? data_i[940] : 1'b0;
  assign data_o[257] = (N1)? data_i[257] : 
                       (N0)? data_i[939] : 1'b0;
  assign data_o[256] = (N1)? data_i[256] : 
                       (N0)? data_i[938] : 1'b0;
  assign data_o[255] = (N1)? data_i[255] : 
                       (N0)? data_i[937] : 1'b0;
  assign data_o[254] = (N1)? data_i[254] : 
                       (N0)? data_i[936] : 1'b0;
  assign data_o[253] = (N1)? data_i[253] : 
                       (N0)? data_i[935] : 1'b0;
  assign data_o[252] = (N1)? data_i[252] : 
                       (N0)? data_i[934] : 1'b0;
  assign data_o[251] = (N1)? data_i[251] : 
                       (N0)? data_i[933] : 1'b0;
  assign data_o[250] = (N1)? data_i[250] : 
                       (N0)? data_i[932] : 1'b0;
  assign data_o[249] = (N1)? data_i[249] : 
                       (N0)? data_i[931] : 1'b0;
  assign data_o[248] = (N1)? data_i[248] : 
                       (N0)? data_i[930] : 1'b0;
  assign data_o[247] = (N1)? data_i[247] : 
                       (N0)? data_i[929] : 1'b0;
  assign data_o[246] = (N1)? data_i[246] : 
                       (N0)? data_i[928] : 1'b0;
  assign data_o[245] = (N1)? data_i[245] : 
                       (N0)? data_i[927] : 1'b0;
  assign data_o[244] = (N1)? data_i[244] : 
                       (N0)? data_i[926] : 1'b0;
  assign data_o[243] = (N1)? data_i[243] : 
                       (N0)? data_i[925] : 1'b0;
  assign data_o[242] = (N1)? data_i[242] : 
                       (N0)? data_i[924] : 1'b0;
  assign data_o[241] = (N1)? data_i[241] : 
                       (N0)? data_i[923] : 1'b0;
  assign data_o[240] = (N1)? data_i[240] : 
                       (N0)? data_i[922] : 1'b0;
  assign data_o[239] = (N1)? data_i[239] : 
                       (N0)? data_i[921] : 1'b0;
  assign data_o[238] = (N1)? data_i[238] : 
                       (N0)? data_i[920] : 1'b0;
  assign data_o[237] = (N1)? data_i[237] : 
                       (N0)? data_i[919] : 1'b0;
  assign data_o[236] = (N1)? data_i[236] : 
                       (N0)? data_i[918] : 1'b0;
  assign data_o[235] = (N1)? data_i[235] : 
                       (N0)? data_i[917] : 1'b0;
  assign data_o[234] = (N1)? data_i[234] : 
                       (N0)? data_i[916] : 1'b0;
  assign data_o[233] = (N1)? data_i[233] : 
                       (N0)? data_i[915] : 1'b0;
  assign data_o[232] = (N1)? data_i[232] : 
                       (N0)? data_i[914] : 1'b0;
  assign data_o[231] = (N1)? data_i[231] : 
                       (N0)? data_i[913] : 1'b0;
  assign data_o[230] = (N1)? data_i[230] : 
                       (N0)? data_i[912] : 1'b0;
  assign data_o[229] = (N1)? data_i[229] : 
                       (N0)? data_i[911] : 1'b0;
  assign data_o[228] = (N1)? data_i[228] : 
                       (N0)? data_i[910] : 1'b0;
  assign data_o[227] = (N1)? data_i[227] : 
                       (N0)? data_i[909] : 1'b0;
  assign data_o[226] = (N1)? data_i[226] : 
                       (N0)? data_i[908] : 1'b0;
  assign data_o[225] = (N1)? data_i[225] : 
                       (N0)? data_i[907] : 1'b0;
  assign data_o[224] = (N1)? data_i[224] : 
                       (N0)? data_i[906] : 1'b0;
  assign data_o[223] = (N1)? data_i[223] : 
                       (N0)? data_i[905] : 1'b0;
  assign data_o[222] = (N1)? data_i[222] : 
                       (N0)? data_i[904] : 1'b0;
  assign data_o[221] = (N1)? data_i[221] : 
                       (N0)? data_i[903] : 1'b0;
  assign data_o[220] = (N1)? data_i[220] : 
                       (N0)? data_i[902] : 1'b0;
  assign data_o[219] = (N1)? data_i[219] : 
                       (N0)? data_i[901] : 1'b0;
  assign data_o[218] = (N1)? data_i[218] : 
                       (N0)? data_i[900] : 1'b0;
  assign data_o[217] = (N1)? data_i[217] : 
                       (N0)? data_i[899] : 1'b0;
  assign data_o[216] = (N1)? data_i[216] : 
                       (N0)? data_i[898] : 1'b0;
  assign data_o[215] = (N1)? data_i[215] : 
                       (N0)? data_i[897] : 1'b0;
  assign data_o[214] = (N1)? data_i[214] : 
                       (N0)? data_i[896] : 1'b0;
  assign data_o[213] = (N1)? data_i[213] : 
                       (N0)? data_i[895] : 1'b0;
  assign data_o[212] = (N1)? data_i[212] : 
                       (N0)? data_i[894] : 1'b0;
  assign data_o[211] = (N1)? data_i[211] : 
                       (N0)? data_i[893] : 1'b0;
  assign data_o[210] = (N1)? data_i[210] : 
                       (N0)? data_i[892] : 1'b0;
  assign data_o[209] = (N1)? data_i[209] : 
                       (N0)? data_i[891] : 1'b0;
  assign data_o[208] = (N1)? data_i[208] : 
                       (N0)? data_i[890] : 1'b0;
  assign data_o[207] = (N1)? data_i[207] : 
                       (N0)? data_i[889] : 1'b0;
  assign data_o[206] = (N1)? data_i[206] : 
                       (N0)? data_i[888] : 1'b0;
  assign data_o[205] = (N1)? data_i[205] : 
                       (N0)? data_i[887] : 1'b0;
  assign data_o[204] = (N1)? data_i[204] : 
                       (N0)? data_i[886] : 1'b0;
  assign data_o[203] = (N1)? data_i[203] : 
                       (N0)? data_i[885] : 1'b0;
  assign data_o[202] = (N1)? data_i[202] : 
                       (N0)? data_i[884] : 1'b0;
  assign data_o[201] = (N1)? data_i[201] : 
                       (N0)? data_i[883] : 1'b0;
  assign data_o[200] = (N1)? data_i[200] : 
                       (N0)? data_i[882] : 1'b0;
  assign data_o[199] = (N1)? data_i[199] : 
                       (N0)? data_i[881] : 1'b0;
  assign data_o[198] = (N1)? data_i[198] : 
                       (N0)? data_i[880] : 1'b0;
  assign data_o[197] = (N1)? data_i[197] : 
                       (N0)? data_i[879] : 1'b0;
  assign data_o[196] = (N1)? data_i[196] : 
                       (N0)? data_i[878] : 1'b0;
  assign data_o[195] = (N1)? data_i[195] : 
                       (N0)? data_i[877] : 1'b0;
  assign data_o[194] = (N1)? data_i[194] : 
                       (N0)? data_i[876] : 1'b0;
  assign data_o[193] = (N1)? data_i[193] : 
                       (N0)? data_i[875] : 1'b0;
  assign data_o[192] = (N1)? data_i[192] : 
                       (N0)? data_i[874] : 1'b0;
  assign data_o[191] = (N1)? data_i[191] : 
                       (N0)? data_i[873] : 1'b0;
  assign data_o[190] = (N1)? data_i[190] : 
                       (N0)? data_i[872] : 1'b0;
  assign data_o[189] = (N1)? data_i[189] : 
                       (N0)? data_i[871] : 1'b0;
  assign data_o[188] = (N1)? data_i[188] : 
                       (N0)? data_i[870] : 1'b0;
  assign data_o[187] = (N1)? data_i[187] : 
                       (N0)? data_i[869] : 1'b0;
  assign data_o[186] = (N1)? data_i[186] : 
                       (N0)? data_i[868] : 1'b0;
  assign data_o[185] = (N1)? data_i[185] : 
                       (N0)? data_i[867] : 1'b0;
  assign data_o[184] = (N1)? data_i[184] : 
                       (N0)? data_i[866] : 1'b0;
  assign data_o[183] = (N1)? data_i[183] : 
                       (N0)? data_i[865] : 1'b0;
  assign data_o[182] = (N1)? data_i[182] : 
                       (N0)? data_i[864] : 1'b0;
  assign data_o[181] = (N1)? data_i[181] : 
                       (N0)? data_i[863] : 1'b0;
  assign data_o[180] = (N1)? data_i[180] : 
                       (N0)? data_i[862] : 1'b0;
  assign data_o[179] = (N1)? data_i[179] : 
                       (N0)? data_i[861] : 1'b0;
  assign data_o[178] = (N1)? data_i[178] : 
                       (N0)? data_i[860] : 1'b0;
  assign data_o[177] = (N1)? data_i[177] : 
                       (N0)? data_i[859] : 1'b0;
  assign data_o[176] = (N1)? data_i[176] : 
                       (N0)? data_i[858] : 1'b0;
  assign data_o[175] = (N1)? data_i[175] : 
                       (N0)? data_i[857] : 1'b0;
  assign data_o[174] = (N1)? data_i[174] : 
                       (N0)? data_i[856] : 1'b0;
  assign data_o[173] = (N1)? data_i[173] : 
                       (N0)? data_i[855] : 1'b0;
  assign data_o[172] = (N1)? data_i[172] : 
                       (N0)? data_i[854] : 1'b0;
  assign data_o[171] = (N1)? data_i[171] : 
                       (N0)? data_i[853] : 1'b0;
  assign data_o[170] = (N1)? data_i[170] : 
                       (N0)? data_i[852] : 1'b0;
  assign data_o[169] = (N1)? data_i[169] : 
                       (N0)? data_i[851] : 1'b0;
  assign data_o[168] = (N1)? data_i[168] : 
                       (N0)? data_i[850] : 1'b0;
  assign data_o[167] = (N1)? data_i[167] : 
                       (N0)? data_i[849] : 1'b0;
  assign data_o[166] = (N1)? data_i[166] : 
                       (N0)? data_i[848] : 1'b0;
  assign data_o[165] = (N1)? data_i[165] : 
                       (N0)? data_i[847] : 1'b0;
  assign data_o[164] = (N1)? data_i[164] : 
                       (N0)? data_i[846] : 1'b0;
  assign data_o[163] = (N1)? data_i[163] : 
                       (N0)? data_i[845] : 1'b0;
  assign data_o[162] = (N1)? data_i[162] : 
                       (N0)? data_i[844] : 1'b0;
  assign data_o[161] = (N1)? data_i[161] : 
                       (N0)? data_i[843] : 1'b0;
  assign data_o[160] = (N1)? data_i[160] : 
                       (N0)? data_i[842] : 1'b0;
  assign data_o[159] = (N1)? data_i[159] : 
                       (N0)? data_i[841] : 1'b0;
  assign data_o[158] = (N1)? data_i[158] : 
                       (N0)? data_i[840] : 1'b0;
  assign data_o[157] = (N1)? data_i[157] : 
                       (N0)? data_i[839] : 1'b0;
  assign data_o[156] = (N1)? data_i[156] : 
                       (N0)? data_i[838] : 1'b0;
  assign data_o[155] = (N1)? data_i[155] : 
                       (N0)? data_i[837] : 1'b0;
  assign data_o[154] = (N1)? data_i[154] : 
                       (N0)? data_i[836] : 1'b0;
  assign data_o[153] = (N1)? data_i[153] : 
                       (N0)? data_i[835] : 1'b0;
  assign data_o[152] = (N1)? data_i[152] : 
                       (N0)? data_i[834] : 1'b0;
  assign data_o[151] = (N1)? data_i[151] : 
                       (N0)? data_i[833] : 1'b0;
  assign data_o[150] = (N1)? data_i[150] : 
                       (N0)? data_i[832] : 1'b0;
  assign data_o[149] = (N1)? data_i[149] : 
                       (N0)? data_i[831] : 1'b0;
  assign data_o[148] = (N1)? data_i[148] : 
                       (N0)? data_i[830] : 1'b0;
  assign data_o[147] = (N1)? data_i[147] : 
                       (N0)? data_i[829] : 1'b0;
  assign data_o[146] = (N1)? data_i[146] : 
                       (N0)? data_i[828] : 1'b0;
  assign data_o[145] = (N1)? data_i[145] : 
                       (N0)? data_i[827] : 1'b0;
  assign data_o[144] = (N1)? data_i[144] : 
                       (N0)? data_i[826] : 1'b0;
  assign data_o[143] = (N1)? data_i[143] : 
                       (N0)? data_i[825] : 1'b0;
  assign data_o[142] = (N1)? data_i[142] : 
                       (N0)? data_i[824] : 1'b0;
  assign data_o[141] = (N1)? data_i[141] : 
                       (N0)? data_i[823] : 1'b0;
  assign data_o[140] = (N1)? data_i[140] : 
                       (N0)? data_i[822] : 1'b0;
  assign data_o[139] = (N1)? data_i[139] : 
                       (N0)? data_i[821] : 1'b0;
  assign data_o[138] = (N1)? data_i[138] : 
                       (N0)? data_i[820] : 1'b0;
  assign data_o[137] = (N1)? data_i[137] : 
                       (N0)? data_i[819] : 1'b0;
  assign data_o[136] = (N1)? data_i[136] : 
                       (N0)? data_i[818] : 1'b0;
  assign data_o[135] = (N1)? data_i[135] : 
                       (N0)? data_i[817] : 1'b0;
  assign data_o[134] = (N1)? data_i[134] : 
                       (N0)? data_i[816] : 1'b0;
  assign data_o[133] = (N1)? data_i[133] : 
                       (N0)? data_i[815] : 1'b0;
  assign data_o[132] = (N1)? data_i[132] : 
                       (N0)? data_i[814] : 1'b0;
  assign data_o[131] = (N1)? data_i[131] : 
                       (N0)? data_i[813] : 1'b0;
  assign data_o[130] = (N1)? data_i[130] : 
                       (N0)? data_i[812] : 1'b0;
  assign data_o[129] = (N1)? data_i[129] : 
                       (N0)? data_i[811] : 1'b0;
  assign data_o[128] = (N1)? data_i[128] : 
                       (N0)? data_i[810] : 1'b0;
  assign data_o[127] = (N1)? data_i[127] : 
                       (N0)? data_i[809] : 1'b0;
  assign data_o[126] = (N1)? data_i[126] : 
                       (N0)? data_i[808] : 1'b0;
  assign data_o[125] = (N1)? data_i[125] : 
                       (N0)? data_i[807] : 1'b0;
  assign data_o[124] = (N1)? data_i[124] : 
                       (N0)? data_i[806] : 1'b0;
  assign data_o[123] = (N1)? data_i[123] : 
                       (N0)? data_i[805] : 1'b0;
  assign data_o[122] = (N1)? data_i[122] : 
                       (N0)? data_i[804] : 1'b0;
  assign data_o[121] = (N1)? data_i[121] : 
                       (N0)? data_i[803] : 1'b0;
  assign data_o[120] = (N1)? data_i[120] : 
                       (N0)? data_i[802] : 1'b0;
  assign data_o[119] = (N1)? data_i[119] : 
                       (N0)? data_i[801] : 1'b0;
  assign data_o[118] = (N1)? data_i[118] : 
                       (N0)? data_i[800] : 1'b0;
  assign data_o[117] = (N1)? data_i[117] : 
                       (N0)? data_i[799] : 1'b0;
  assign data_o[116] = (N1)? data_i[116] : 
                       (N0)? data_i[798] : 1'b0;
  assign data_o[115] = (N1)? data_i[115] : 
                       (N0)? data_i[797] : 1'b0;
  assign data_o[114] = (N1)? data_i[114] : 
                       (N0)? data_i[796] : 1'b0;
  assign data_o[113] = (N1)? data_i[113] : 
                       (N0)? data_i[795] : 1'b0;
  assign data_o[112] = (N1)? data_i[112] : 
                       (N0)? data_i[794] : 1'b0;
  assign data_o[111] = (N1)? data_i[111] : 
                       (N0)? data_i[793] : 1'b0;
  assign data_o[110] = (N1)? data_i[110] : 
                       (N0)? data_i[792] : 1'b0;
  assign data_o[109] = (N1)? data_i[109] : 
                       (N0)? data_i[791] : 1'b0;
  assign data_o[108] = (N1)? data_i[108] : 
                       (N0)? data_i[790] : 1'b0;
  assign data_o[107] = (N1)? data_i[107] : 
                       (N0)? data_i[789] : 1'b0;
  assign data_o[106] = (N1)? data_i[106] : 
                       (N0)? data_i[788] : 1'b0;
  assign data_o[105] = (N1)? data_i[105] : 
                       (N0)? data_i[787] : 1'b0;
  assign data_o[104] = (N1)? data_i[104] : 
                       (N0)? data_i[786] : 1'b0;
  assign data_o[103] = (N1)? data_i[103] : 
                       (N0)? data_i[785] : 1'b0;
  assign data_o[102] = (N1)? data_i[102] : 
                       (N0)? data_i[784] : 1'b0;
  assign data_o[101] = (N1)? data_i[101] : 
                       (N0)? data_i[783] : 1'b0;
  assign data_o[100] = (N1)? data_i[100] : 
                       (N0)? data_i[782] : 1'b0;
  assign data_o[99] = (N1)? data_i[99] : 
                      (N0)? data_i[781] : 1'b0;
  assign data_o[98] = (N1)? data_i[98] : 
                      (N0)? data_i[780] : 1'b0;
  assign data_o[97] = (N1)? data_i[97] : 
                      (N0)? data_i[779] : 1'b0;
  assign data_o[96] = (N1)? data_i[96] : 
                      (N0)? data_i[778] : 1'b0;
  assign data_o[95] = (N1)? data_i[95] : 
                      (N0)? data_i[777] : 1'b0;
  assign data_o[94] = (N1)? data_i[94] : 
                      (N0)? data_i[776] : 1'b0;
  assign data_o[93] = (N1)? data_i[93] : 
                      (N0)? data_i[775] : 1'b0;
  assign data_o[92] = (N1)? data_i[92] : 
                      (N0)? data_i[774] : 1'b0;
  assign data_o[91] = (N1)? data_i[91] : 
                      (N0)? data_i[773] : 1'b0;
  assign data_o[90] = (N1)? data_i[90] : 
                      (N0)? data_i[772] : 1'b0;
  assign data_o[89] = (N1)? data_i[89] : 
                      (N0)? data_i[771] : 1'b0;
  assign data_o[88] = (N1)? data_i[88] : 
                      (N0)? data_i[770] : 1'b0;
  assign data_o[87] = (N1)? data_i[87] : 
                      (N0)? data_i[769] : 1'b0;
  assign data_o[86] = (N1)? data_i[86] : 
                      (N0)? data_i[768] : 1'b0;
  assign data_o[85] = (N1)? data_i[85] : 
                      (N0)? data_i[767] : 1'b0;
  assign data_o[84] = (N1)? data_i[84] : 
                      (N0)? data_i[766] : 1'b0;
  assign data_o[83] = (N1)? data_i[83] : 
                      (N0)? data_i[765] : 1'b0;
  assign data_o[82] = (N1)? data_i[82] : 
                      (N0)? data_i[764] : 1'b0;
  assign data_o[81] = (N1)? data_i[81] : 
                      (N0)? data_i[763] : 1'b0;
  assign data_o[80] = (N1)? data_i[80] : 
                      (N0)? data_i[762] : 1'b0;
  assign data_o[79] = (N1)? data_i[79] : 
                      (N0)? data_i[761] : 1'b0;
  assign data_o[78] = (N1)? data_i[78] : 
                      (N0)? data_i[760] : 1'b0;
  assign data_o[77] = (N1)? data_i[77] : 
                      (N0)? data_i[759] : 1'b0;
  assign data_o[76] = (N1)? data_i[76] : 
                      (N0)? data_i[758] : 1'b0;
  assign data_o[75] = (N1)? data_i[75] : 
                      (N0)? data_i[757] : 1'b0;
  assign data_o[74] = (N1)? data_i[74] : 
                      (N0)? data_i[756] : 1'b0;
  assign data_o[73] = (N1)? data_i[73] : 
                      (N0)? data_i[755] : 1'b0;
  assign data_o[72] = (N1)? data_i[72] : 
                      (N0)? data_i[754] : 1'b0;
  assign data_o[71] = (N1)? data_i[71] : 
                      (N0)? data_i[753] : 1'b0;
  assign data_o[70] = (N1)? data_i[70] : 
                      (N0)? data_i[752] : 1'b0;
  assign data_o[69] = (N1)? data_i[69] : 
                      (N0)? data_i[751] : 1'b0;
  assign data_o[68] = (N1)? data_i[68] : 
                      (N0)? data_i[750] : 1'b0;
  assign data_o[67] = (N1)? data_i[67] : 
                      (N0)? data_i[749] : 1'b0;
  assign data_o[66] = (N1)? data_i[66] : 
                      (N0)? data_i[748] : 1'b0;
  assign data_o[65] = (N1)? data_i[65] : 
                      (N0)? data_i[747] : 1'b0;
  assign data_o[64] = (N1)? data_i[64] : 
                      (N0)? data_i[746] : 1'b0;
  assign data_o[63] = (N1)? data_i[63] : 
                      (N0)? data_i[745] : 1'b0;
  assign data_o[62] = (N1)? data_i[62] : 
                      (N0)? data_i[744] : 1'b0;
  assign data_o[61] = (N1)? data_i[61] : 
                      (N0)? data_i[743] : 1'b0;
  assign data_o[60] = (N1)? data_i[60] : 
                      (N0)? data_i[742] : 1'b0;
  assign data_o[59] = (N1)? data_i[59] : 
                      (N0)? data_i[741] : 1'b0;
  assign data_o[58] = (N1)? data_i[58] : 
                      (N0)? data_i[740] : 1'b0;
  assign data_o[57] = (N1)? data_i[57] : 
                      (N0)? data_i[739] : 1'b0;
  assign data_o[56] = (N1)? data_i[56] : 
                      (N0)? data_i[738] : 1'b0;
  assign data_o[55] = (N1)? data_i[55] : 
                      (N0)? data_i[737] : 1'b0;
  assign data_o[54] = (N1)? data_i[54] : 
                      (N0)? data_i[736] : 1'b0;
  assign data_o[53] = (N1)? data_i[53] : 
                      (N0)? data_i[735] : 1'b0;
  assign data_o[52] = (N1)? data_i[52] : 
                      (N0)? data_i[734] : 1'b0;
  assign data_o[51] = (N1)? data_i[51] : 
                      (N0)? data_i[733] : 1'b0;
  assign data_o[50] = (N1)? data_i[50] : 
                      (N0)? data_i[732] : 1'b0;
  assign data_o[49] = (N1)? data_i[49] : 
                      (N0)? data_i[731] : 1'b0;
  assign data_o[48] = (N1)? data_i[48] : 
                      (N0)? data_i[730] : 1'b0;
  assign data_o[47] = (N1)? data_i[47] : 
                      (N0)? data_i[729] : 1'b0;
  assign data_o[46] = (N1)? data_i[46] : 
                      (N0)? data_i[728] : 1'b0;
  assign data_o[45] = (N1)? data_i[45] : 
                      (N0)? data_i[727] : 1'b0;
  assign data_o[44] = (N1)? data_i[44] : 
                      (N0)? data_i[726] : 1'b0;
  assign data_o[43] = (N1)? data_i[43] : 
                      (N0)? data_i[725] : 1'b0;
  assign data_o[42] = (N1)? data_i[42] : 
                      (N0)? data_i[724] : 1'b0;
  assign data_o[41] = (N1)? data_i[41] : 
                      (N0)? data_i[723] : 1'b0;
  assign data_o[40] = (N1)? data_i[40] : 
                      (N0)? data_i[722] : 1'b0;
  assign data_o[39] = (N1)? data_i[39] : 
                      (N0)? data_i[721] : 1'b0;
  assign data_o[38] = (N1)? data_i[38] : 
                      (N0)? data_i[720] : 1'b0;
  assign data_o[37] = (N1)? data_i[37] : 
                      (N0)? data_i[719] : 1'b0;
  assign data_o[36] = (N1)? data_i[36] : 
                      (N0)? data_i[718] : 1'b0;
  assign data_o[35] = (N1)? data_i[35] : 
                      (N0)? data_i[717] : 1'b0;
  assign data_o[34] = (N1)? data_i[34] : 
                      (N0)? data_i[716] : 1'b0;
  assign data_o[33] = (N1)? data_i[33] : 
                      (N0)? data_i[715] : 1'b0;
  assign data_o[32] = (N1)? data_i[32] : 
                      (N0)? data_i[714] : 1'b0;
  assign data_o[31] = (N1)? data_i[31] : 
                      (N0)? data_i[713] : 1'b0;
  assign data_o[30] = (N1)? data_i[30] : 
                      (N0)? data_i[712] : 1'b0;
  assign data_o[29] = (N1)? data_i[29] : 
                      (N0)? data_i[711] : 1'b0;
  assign data_o[28] = (N1)? data_i[28] : 
                      (N0)? data_i[710] : 1'b0;
  assign data_o[27] = (N1)? data_i[27] : 
                      (N0)? data_i[709] : 1'b0;
  assign data_o[26] = (N1)? data_i[26] : 
                      (N0)? data_i[708] : 1'b0;
  assign data_o[25] = (N1)? data_i[25] : 
                      (N0)? data_i[707] : 1'b0;
  assign data_o[24] = (N1)? data_i[24] : 
                      (N0)? data_i[706] : 1'b0;
  assign data_o[23] = (N1)? data_i[23] : 
                      (N0)? data_i[705] : 1'b0;
  assign data_o[22] = (N1)? data_i[22] : 
                      (N0)? data_i[704] : 1'b0;
  assign data_o[21] = (N1)? data_i[21] : 
                      (N0)? data_i[703] : 1'b0;
  assign data_o[20] = (N1)? data_i[20] : 
                      (N0)? data_i[702] : 1'b0;
  assign data_o[19] = (N1)? data_i[19] : 
                      (N0)? data_i[701] : 1'b0;
  assign data_o[18] = (N1)? data_i[18] : 
                      (N0)? data_i[700] : 1'b0;
  assign data_o[17] = (N1)? data_i[17] : 
                      (N0)? data_i[699] : 1'b0;
  assign data_o[16] = (N1)? data_i[16] : 
                      (N0)? data_i[698] : 1'b0;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[697] : 1'b0;
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[696] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[695] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[694] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[693] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[692] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[691] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[690] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[689] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[688] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[687] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[686] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[685] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[684] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[683] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[682] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_dff_000002ab
(
  clk_i,
  data_i,
  data_o
);

  input [682:0] data_i;
  output [682:0] data_o;
  input clk_i;
  wire [682:0] data_o;
  reg data_o_682_sv2v_reg,data_o_681_sv2v_reg,data_o_680_sv2v_reg,data_o_679_sv2v_reg,
  data_o_678_sv2v_reg,data_o_677_sv2v_reg,data_o_676_sv2v_reg,data_o_675_sv2v_reg,
  data_o_674_sv2v_reg,data_o_673_sv2v_reg,data_o_672_sv2v_reg,data_o_671_sv2v_reg,
  data_o_670_sv2v_reg,data_o_669_sv2v_reg,data_o_668_sv2v_reg,data_o_667_sv2v_reg,
  data_o_666_sv2v_reg,data_o_665_sv2v_reg,data_o_664_sv2v_reg,data_o_663_sv2v_reg,
  data_o_662_sv2v_reg,data_o_661_sv2v_reg,data_o_660_sv2v_reg,data_o_659_sv2v_reg,
  data_o_658_sv2v_reg,data_o_657_sv2v_reg,data_o_656_sv2v_reg,data_o_655_sv2v_reg,
  data_o_654_sv2v_reg,data_o_653_sv2v_reg,data_o_652_sv2v_reg,data_o_651_sv2v_reg,
  data_o_650_sv2v_reg,data_o_649_sv2v_reg,data_o_648_sv2v_reg,data_o_647_sv2v_reg,
  data_o_646_sv2v_reg,data_o_645_sv2v_reg,data_o_644_sv2v_reg,data_o_643_sv2v_reg,
  data_o_642_sv2v_reg,data_o_641_sv2v_reg,data_o_640_sv2v_reg,data_o_639_sv2v_reg,
  data_o_638_sv2v_reg,data_o_637_sv2v_reg,data_o_636_sv2v_reg,data_o_635_sv2v_reg,
  data_o_634_sv2v_reg,data_o_633_sv2v_reg,data_o_632_sv2v_reg,data_o_631_sv2v_reg,
  data_o_630_sv2v_reg,data_o_629_sv2v_reg,data_o_628_sv2v_reg,data_o_627_sv2v_reg,
  data_o_626_sv2v_reg,data_o_625_sv2v_reg,data_o_624_sv2v_reg,data_o_623_sv2v_reg,
  data_o_622_sv2v_reg,data_o_621_sv2v_reg,data_o_620_sv2v_reg,data_o_619_sv2v_reg,
  data_o_618_sv2v_reg,data_o_617_sv2v_reg,data_o_616_sv2v_reg,data_o_615_sv2v_reg,
  data_o_614_sv2v_reg,data_o_613_sv2v_reg,data_o_612_sv2v_reg,data_o_611_sv2v_reg,
  data_o_610_sv2v_reg,data_o_609_sv2v_reg,data_o_608_sv2v_reg,data_o_607_sv2v_reg,
  data_o_606_sv2v_reg,data_o_605_sv2v_reg,data_o_604_sv2v_reg,data_o_603_sv2v_reg,
  data_o_602_sv2v_reg,data_o_601_sv2v_reg,data_o_600_sv2v_reg,data_o_599_sv2v_reg,
  data_o_598_sv2v_reg,data_o_597_sv2v_reg,data_o_596_sv2v_reg,data_o_595_sv2v_reg,
  data_o_594_sv2v_reg,data_o_593_sv2v_reg,data_o_592_sv2v_reg,data_o_591_sv2v_reg,
  data_o_590_sv2v_reg,data_o_589_sv2v_reg,data_o_588_sv2v_reg,data_o_587_sv2v_reg,
  data_o_586_sv2v_reg,data_o_585_sv2v_reg,data_o_584_sv2v_reg,data_o_583_sv2v_reg,
  data_o_582_sv2v_reg,data_o_581_sv2v_reg,data_o_580_sv2v_reg,data_o_579_sv2v_reg,
  data_o_578_sv2v_reg,data_o_577_sv2v_reg,data_o_576_sv2v_reg,data_o_575_sv2v_reg,
  data_o_574_sv2v_reg,data_o_573_sv2v_reg,data_o_572_sv2v_reg,data_o_571_sv2v_reg,
  data_o_570_sv2v_reg,data_o_569_sv2v_reg,data_o_568_sv2v_reg,data_o_567_sv2v_reg,
  data_o_566_sv2v_reg,data_o_565_sv2v_reg,data_o_564_sv2v_reg,data_o_563_sv2v_reg,
  data_o_562_sv2v_reg,data_o_561_sv2v_reg,data_o_560_sv2v_reg,data_o_559_sv2v_reg,
  data_o_558_sv2v_reg,data_o_557_sv2v_reg,data_o_556_sv2v_reg,data_o_555_sv2v_reg,
  data_o_554_sv2v_reg,data_o_553_sv2v_reg,data_o_552_sv2v_reg,data_o_551_sv2v_reg,
  data_o_550_sv2v_reg,data_o_549_sv2v_reg,data_o_548_sv2v_reg,data_o_547_sv2v_reg,
  data_o_546_sv2v_reg,data_o_545_sv2v_reg,data_o_544_sv2v_reg,data_o_543_sv2v_reg,
  data_o_542_sv2v_reg,data_o_541_sv2v_reg,data_o_540_sv2v_reg,data_o_539_sv2v_reg,
  data_o_538_sv2v_reg,data_o_537_sv2v_reg,data_o_536_sv2v_reg,data_o_535_sv2v_reg,
  data_o_534_sv2v_reg,data_o_533_sv2v_reg,data_o_532_sv2v_reg,data_o_531_sv2v_reg,
  data_o_530_sv2v_reg,data_o_529_sv2v_reg,data_o_528_sv2v_reg,data_o_527_sv2v_reg,
  data_o_526_sv2v_reg,data_o_525_sv2v_reg,data_o_524_sv2v_reg,data_o_523_sv2v_reg,
  data_o_522_sv2v_reg,data_o_521_sv2v_reg,data_o_520_sv2v_reg,data_o_519_sv2v_reg,
  data_o_518_sv2v_reg,data_o_517_sv2v_reg,data_o_516_sv2v_reg,data_o_515_sv2v_reg,
  data_o_514_sv2v_reg,data_o_513_sv2v_reg,data_o_512_sv2v_reg,data_o_511_sv2v_reg,
  data_o_510_sv2v_reg,data_o_509_sv2v_reg,data_o_508_sv2v_reg,data_o_507_sv2v_reg,
  data_o_506_sv2v_reg,data_o_505_sv2v_reg,data_o_504_sv2v_reg,data_o_503_sv2v_reg,
  data_o_502_sv2v_reg,data_o_501_sv2v_reg,data_o_500_sv2v_reg,data_o_499_sv2v_reg,
  data_o_498_sv2v_reg,data_o_497_sv2v_reg,data_o_496_sv2v_reg,data_o_495_sv2v_reg,
  data_o_494_sv2v_reg,data_o_493_sv2v_reg,data_o_492_sv2v_reg,data_o_491_sv2v_reg,
  data_o_490_sv2v_reg,data_o_489_sv2v_reg,data_o_488_sv2v_reg,data_o_487_sv2v_reg,
  data_o_486_sv2v_reg,data_o_485_sv2v_reg,data_o_484_sv2v_reg,data_o_483_sv2v_reg,
  data_o_482_sv2v_reg,data_o_481_sv2v_reg,data_o_480_sv2v_reg,data_o_479_sv2v_reg,
  data_o_478_sv2v_reg,data_o_477_sv2v_reg,data_o_476_sv2v_reg,data_o_475_sv2v_reg,
  data_o_474_sv2v_reg,data_o_473_sv2v_reg,data_o_472_sv2v_reg,data_o_471_sv2v_reg,
  data_o_470_sv2v_reg,data_o_469_sv2v_reg,data_o_468_sv2v_reg,data_o_467_sv2v_reg,
  data_o_466_sv2v_reg,data_o_465_sv2v_reg,data_o_464_sv2v_reg,data_o_463_sv2v_reg,
  data_o_462_sv2v_reg,data_o_461_sv2v_reg,data_o_460_sv2v_reg,data_o_459_sv2v_reg,
  data_o_458_sv2v_reg,data_o_457_sv2v_reg,data_o_456_sv2v_reg,data_o_455_sv2v_reg,
  data_o_454_sv2v_reg,data_o_453_sv2v_reg,data_o_452_sv2v_reg,data_o_451_sv2v_reg,
  data_o_450_sv2v_reg,data_o_449_sv2v_reg,data_o_448_sv2v_reg,data_o_447_sv2v_reg,
  data_o_446_sv2v_reg,data_o_445_sv2v_reg,data_o_444_sv2v_reg,data_o_443_sv2v_reg,
  data_o_442_sv2v_reg,data_o_441_sv2v_reg,data_o_440_sv2v_reg,data_o_439_sv2v_reg,
  data_o_438_sv2v_reg,data_o_437_sv2v_reg,data_o_436_sv2v_reg,data_o_435_sv2v_reg,
  data_o_434_sv2v_reg,data_o_433_sv2v_reg,data_o_432_sv2v_reg,data_o_431_sv2v_reg,
  data_o_430_sv2v_reg,data_o_429_sv2v_reg,data_o_428_sv2v_reg,data_o_427_sv2v_reg,
  data_o_426_sv2v_reg,data_o_425_sv2v_reg,data_o_424_sv2v_reg,data_o_423_sv2v_reg,
  data_o_422_sv2v_reg,data_o_421_sv2v_reg,data_o_420_sv2v_reg,data_o_419_sv2v_reg,
  data_o_418_sv2v_reg,data_o_417_sv2v_reg,data_o_416_sv2v_reg,data_o_415_sv2v_reg,
  data_o_414_sv2v_reg,data_o_413_sv2v_reg,data_o_412_sv2v_reg,data_o_411_sv2v_reg,
  data_o_410_sv2v_reg,data_o_409_sv2v_reg,data_o_408_sv2v_reg,data_o_407_sv2v_reg,
  data_o_406_sv2v_reg,data_o_405_sv2v_reg,data_o_404_sv2v_reg,data_o_403_sv2v_reg,
  data_o_402_sv2v_reg,data_o_401_sv2v_reg,data_o_400_sv2v_reg,data_o_399_sv2v_reg,
  data_o_398_sv2v_reg,data_o_397_sv2v_reg,data_o_396_sv2v_reg,data_o_395_sv2v_reg,
  data_o_394_sv2v_reg,data_o_393_sv2v_reg,data_o_392_sv2v_reg,data_o_391_sv2v_reg,
  data_o_390_sv2v_reg,data_o_389_sv2v_reg,data_o_388_sv2v_reg,data_o_387_sv2v_reg,
  data_o_386_sv2v_reg,data_o_385_sv2v_reg,data_o_384_sv2v_reg,data_o_383_sv2v_reg,
  data_o_382_sv2v_reg,data_o_381_sv2v_reg,data_o_380_sv2v_reg,data_o_379_sv2v_reg,
  data_o_378_sv2v_reg,data_o_377_sv2v_reg,data_o_376_sv2v_reg,data_o_375_sv2v_reg,
  data_o_374_sv2v_reg,data_o_373_sv2v_reg,data_o_372_sv2v_reg,data_o_371_sv2v_reg,
  data_o_370_sv2v_reg,data_o_369_sv2v_reg,data_o_368_sv2v_reg,data_o_367_sv2v_reg,
  data_o_366_sv2v_reg,data_o_365_sv2v_reg,data_o_364_sv2v_reg,data_o_363_sv2v_reg,
  data_o_362_sv2v_reg,data_o_361_sv2v_reg,data_o_360_sv2v_reg,data_o_359_sv2v_reg,
  data_o_358_sv2v_reg,data_o_357_sv2v_reg,data_o_356_sv2v_reg,data_o_355_sv2v_reg,
  data_o_354_sv2v_reg,data_o_353_sv2v_reg,data_o_352_sv2v_reg,data_o_351_sv2v_reg,
  data_o_350_sv2v_reg,data_o_349_sv2v_reg,data_o_348_sv2v_reg,data_o_347_sv2v_reg,
  data_o_346_sv2v_reg,data_o_345_sv2v_reg,data_o_344_sv2v_reg,data_o_343_sv2v_reg,
  data_o_342_sv2v_reg,data_o_341_sv2v_reg,data_o_340_sv2v_reg,data_o_339_sv2v_reg,
  data_o_338_sv2v_reg,data_o_337_sv2v_reg,data_o_336_sv2v_reg,data_o_335_sv2v_reg,
  data_o_334_sv2v_reg,data_o_333_sv2v_reg,data_o_332_sv2v_reg,data_o_331_sv2v_reg,
  data_o_330_sv2v_reg,data_o_329_sv2v_reg,data_o_328_sv2v_reg,data_o_327_sv2v_reg,
  data_o_326_sv2v_reg,data_o_325_sv2v_reg,data_o_324_sv2v_reg,data_o_323_sv2v_reg,
  data_o_322_sv2v_reg,data_o_321_sv2v_reg,data_o_320_sv2v_reg,data_o_319_sv2v_reg,
  data_o_318_sv2v_reg,data_o_317_sv2v_reg,data_o_316_sv2v_reg,data_o_315_sv2v_reg,
  data_o_314_sv2v_reg,data_o_313_sv2v_reg,data_o_312_sv2v_reg,data_o_311_sv2v_reg,
  data_o_310_sv2v_reg,data_o_309_sv2v_reg,data_o_308_sv2v_reg,data_o_307_sv2v_reg,
  data_o_306_sv2v_reg,data_o_305_sv2v_reg,data_o_304_sv2v_reg,data_o_303_sv2v_reg,
  data_o_302_sv2v_reg,data_o_301_sv2v_reg,data_o_300_sv2v_reg,data_o_299_sv2v_reg,
  data_o_298_sv2v_reg,data_o_297_sv2v_reg,data_o_296_sv2v_reg,data_o_295_sv2v_reg,
  data_o_294_sv2v_reg,data_o_293_sv2v_reg,data_o_292_sv2v_reg,data_o_291_sv2v_reg,
  data_o_290_sv2v_reg,data_o_289_sv2v_reg,data_o_288_sv2v_reg,data_o_287_sv2v_reg,
  data_o_286_sv2v_reg,data_o_285_sv2v_reg,data_o_284_sv2v_reg,data_o_283_sv2v_reg,
  data_o_282_sv2v_reg,data_o_281_sv2v_reg,data_o_280_sv2v_reg,data_o_279_sv2v_reg,
  data_o_278_sv2v_reg,data_o_277_sv2v_reg,data_o_276_sv2v_reg,data_o_275_sv2v_reg,
  data_o_274_sv2v_reg,data_o_273_sv2v_reg,data_o_272_sv2v_reg,data_o_271_sv2v_reg,
  data_o_270_sv2v_reg,data_o_269_sv2v_reg,data_o_268_sv2v_reg,data_o_267_sv2v_reg,
  data_o_266_sv2v_reg,data_o_265_sv2v_reg,data_o_264_sv2v_reg,data_o_263_sv2v_reg,
  data_o_262_sv2v_reg,data_o_261_sv2v_reg,data_o_260_sv2v_reg,data_o_259_sv2v_reg,
  data_o_258_sv2v_reg,data_o_257_sv2v_reg,data_o_256_sv2v_reg,data_o_255_sv2v_reg,
  data_o_254_sv2v_reg,data_o_253_sv2v_reg,data_o_252_sv2v_reg,data_o_251_sv2v_reg,
  data_o_250_sv2v_reg,data_o_249_sv2v_reg,data_o_248_sv2v_reg,data_o_247_sv2v_reg,
  data_o_246_sv2v_reg,data_o_245_sv2v_reg,data_o_244_sv2v_reg,data_o_243_sv2v_reg,
  data_o_242_sv2v_reg,data_o_241_sv2v_reg,data_o_240_sv2v_reg,data_o_239_sv2v_reg,
  data_o_238_sv2v_reg,data_o_237_sv2v_reg,data_o_236_sv2v_reg,data_o_235_sv2v_reg,
  data_o_234_sv2v_reg,data_o_233_sv2v_reg,data_o_232_sv2v_reg,data_o_231_sv2v_reg,
  data_o_230_sv2v_reg,data_o_229_sv2v_reg,data_o_228_sv2v_reg,data_o_227_sv2v_reg,
  data_o_226_sv2v_reg,data_o_225_sv2v_reg,data_o_224_sv2v_reg,data_o_223_sv2v_reg,
  data_o_222_sv2v_reg,data_o_221_sv2v_reg,data_o_220_sv2v_reg,data_o_219_sv2v_reg,
  data_o_218_sv2v_reg,data_o_217_sv2v_reg,data_o_216_sv2v_reg,data_o_215_sv2v_reg,
  data_o_214_sv2v_reg,data_o_213_sv2v_reg,data_o_212_sv2v_reg,data_o_211_sv2v_reg,
  data_o_210_sv2v_reg,data_o_209_sv2v_reg,data_o_208_sv2v_reg,data_o_207_sv2v_reg,
  data_o_206_sv2v_reg,data_o_205_sv2v_reg,data_o_204_sv2v_reg,data_o_203_sv2v_reg,
  data_o_202_sv2v_reg,data_o_201_sv2v_reg,data_o_200_sv2v_reg,data_o_199_sv2v_reg,
  data_o_198_sv2v_reg,data_o_197_sv2v_reg,data_o_196_sv2v_reg,data_o_195_sv2v_reg,
  data_o_194_sv2v_reg,data_o_193_sv2v_reg,data_o_192_sv2v_reg,data_o_191_sv2v_reg,
  data_o_190_sv2v_reg,data_o_189_sv2v_reg,data_o_188_sv2v_reg,data_o_187_sv2v_reg,
  data_o_186_sv2v_reg,data_o_185_sv2v_reg,data_o_184_sv2v_reg,data_o_183_sv2v_reg,
  data_o_182_sv2v_reg,data_o_181_sv2v_reg,data_o_180_sv2v_reg,data_o_179_sv2v_reg,
  data_o_178_sv2v_reg,data_o_177_sv2v_reg,data_o_176_sv2v_reg,data_o_175_sv2v_reg,
  data_o_174_sv2v_reg,data_o_173_sv2v_reg,data_o_172_sv2v_reg,data_o_171_sv2v_reg,
  data_o_170_sv2v_reg,data_o_169_sv2v_reg,data_o_168_sv2v_reg,data_o_167_sv2v_reg,
  data_o_166_sv2v_reg,data_o_165_sv2v_reg,data_o_164_sv2v_reg,data_o_163_sv2v_reg,
  data_o_162_sv2v_reg,data_o_161_sv2v_reg,data_o_160_sv2v_reg,data_o_159_sv2v_reg,
  data_o_158_sv2v_reg,data_o_157_sv2v_reg,data_o_156_sv2v_reg,data_o_155_sv2v_reg,
  data_o_154_sv2v_reg,data_o_153_sv2v_reg,data_o_152_sv2v_reg,data_o_151_sv2v_reg,
  data_o_150_sv2v_reg,data_o_149_sv2v_reg,data_o_148_sv2v_reg,data_o_147_sv2v_reg,
  data_o_146_sv2v_reg,data_o_145_sv2v_reg,data_o_144_sv2v_reg,data_o_143_sv2v_reg,
  data_o_142_sv2v_reg,data_o_141_sv2v_reg,data_o_140_sv2v_reg,data_o_139_sv2v_reg,
  data_o_138_sv2v_reg,data_o_137_sv2v_reg,data_o_136_sv2v_reg,data_o_135_sv2v_reg,
  data_o_134_sv2v_reg,data_o_133_sv2v_reg,data_o_132_sv2v_reg,data_o_131_sv2v_reg,
  data_o_130_sv2v_reg,data_o_129_sv2v_reg,data_o_128_sv2v_reg,data_o_127_sv2v_reg,
  data_o_126_sv2v_reg,data_o_125_sv2v_reg,data_o_124_sv2v_reg,data_o_123_sv2v_reg,
  data_o_122_sv2v_reg,data_o_121_sv2v_reg,data_o_120_sv2v_reg,data_o_119_sv2v_reg,
  data_o_118_sv2v_reg,data_o_117_sv2v_reg,data_o_116_sv2v_reg,data_o_115_sv2v_reg,
  data_o_114_sv2v_reg,data_o_113_sv2v_reg,data_o_112_sv2v_reg,data_o_111_sv2v_reg,
  data_o_110_sv2v_reg,data_o_109_sv2v_reg,data_o_108_sv2v_reg,data_o_107_sv2v_reg,
  data_o_106_sv2v_reg,data_o_105_sv2v_reg,data_o_104_sv2v_reg,data_o_103_sv2v_reg,
  data_o_102_sv2v_reg,data_o_101_sv2v_reg,data_o_100_sv2v_reg,data_o_99_sv2v_reg,
  data_o_98_sv2v_reg,data_o_97_sv2v_reg,data_o_96_sv2v_reg,data_o_95_sv2v_reg,
  data_o_94_sv2v_reg,data_o_93_sv2v_reg,data_o_92_sv2v_reg,data_o_91_sv2v_reg,
  data_o_90_sv2v_reg,data_o_89_sv2v_reg,data_o_88_sv2v_reg,data_o_87_sv2v_reg,
  data_o_86_sv2v_reg,data_o_85_sv2v_reg,data_o_84_sv2v_reg,data_o_83_sv2v_reg,
  data_o_82_sv2v_reg,data_o_81_sv2v_reg,data_o_80_sv2v_reg,data_o_79_sv2v_reg,data_o_78_sv2v_reg,
  data_o_77_sv2v_reg,data_o_76_sv2v_reg,data_o_75_sv2v_reg,data_o_74_sv2v_reg,
  data_o_73_sv2v_reg,data_o_72_sv2v_reg,data_o_71_sv2v_reg,data_o_70_sv2v_reg,
  data_o_69_sv2v_reg,data_o_68_sv2v_reg,data_o_67_sv2v_reg,data_o_66_sv2v_reg,
  data_o_65_sv2v_reg,data_o_64_sv2v_reg,data_o_63_sv2v_reg,data_o_62_sv2v_reg,
  data_o_61_sv2v_reg,data_o_60_sv2v_reg,data_o_59_sv2v_reg,data_o_58_sv2v_reg,data_o_57_sv2v_reg,
  data_o_56_sv2v_reg,data_o_55_sv2v_reg,data_o_54_sv2v_reg,data_o_53_sv2v_reg,
  data_o_52_sv2v_reg,data_o_51_sv2v_reg,data_o_50_sv2v_reg,data_o_49_sv2v_reg,
  data_o_48_sv2v_reg,data_o_47_sv2v_reg,data_o_46_sv2v_reg,data_o_45_sv2v_reg,
  data_o_44_sv2v_reg,data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,
  data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,
  data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,
  data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,
  data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,
  data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[682] = data_o_682_sv2v_reg;
  assign data_o[681] = data_o_681_sv2v_reg;
  assign data_o[680] = data_o_680_sv2v_reg;
  assign data_o[679] = data_o_679_sv2v_reg;
  assign data_o[678] = data_o_678_sv2v_reg;
  assign data_o[677] = data_o_677_sv2v_reg;
  assign data_o[676] = data_o_676_sv2v_reg;
  assign data_o[675] = data_o_675_sv2v_reg;
  assign data_o[674] = data_o_674_sv2v_reg;
  assign data_o[673] = data_o_673_sv2v_reg;
  assign data_o[672] = data_o_672_sv2v_reg;
  assign data_o[671] = data_o_671_sv2v_reg;
  assign data_o[670] = data_o_670_sv2v_reg;
  assign data_o[669] = data_o_669_sv2v_reg;
  assign data_o[668] = data_o_668_sv2v_reg;
  assign data_o[667] = data_o_667_sv2v_reg;
  assign data_o[666] = data_o_666_sv2v_reg;
  assign data_o[665] = data_o_665_sv2v_reg;
  assign data_o[664] = data_o_664_sv2v_reg;
  assign data_o[663] = data_o_663_sv2v_reg;
  assign data_o[662] = data_o_662_sv2v_reg;
  assign data_o[661] = data_o_661_sv2v_reg;
  assign data_o[660] = data_o_660_sv2v_reg;
  assign data_o[659] = data_o_659_sv2v_reg;
  assign data_o[658] = data_o_658_sv2v_reg;
  assign data_o[657] = data_o_657_sv2v_reg;
  assign data_o[656] = data_o_656_sv2v_reg;
  assign data_o[655] = data_o_655_sv2v_reg;
  assign data_o[654] = data_o_654_sv2v_reg;
  assign data_o[653] = data_o_653_sv2v_reg;
  assign data_o[652] = data_o_652_sv2v_reg;
  assign data_o[651] = data_o_651_sv2v_reg;
  assign data_o[650] = data_o_650_sv2v_reg;
  assign data_o[649] = data_o_649_sv2v_reg;
  assign data_o[648] = data_o_648_sv2v_reg;
  assign data_o[647] = data_o_647_sv2v_reg;
  assign data_o[646] = data_o_646_sv2v_reg;
  assign data_o[645] = data_o_645_sv2v_reg;
  assign data_o[644] = data_o_644_sv2v_reg;
  assign data_o[643] = data_o_643_sv2v_reg;
  assign data_o[642] = data_o_642_sv2v_reg;
  assign data_o[641] = data_o_641_sv2v_reg;
  assign data_o[640] = data_o_640_sv2v_reg;
  assign data_o[639] = data_o_639_sv2v_reg;
  assign data_o[638] = data_o_638_sv2v_reg;
  assign data_o[637] = data_o_637_sv2v_reg;
  assign data_o[636] = data_o_636_sv2v_reg;
  assign data_o[635] = data_o_635_sv2v_reg;
  assign data_o[634] = data_o_634_sv2v_reg;
  assign data_o[633] = data_o_633_sv2v_reg;
  assign data_o[632] = data_o_632_sv2v_reg;
  assign data_o[631] = data_o_631_sv2v_reg;
  assign data_o[630] = data_o_630_sv2v_reg;
  assign data_o[629] = data_o_629_sv2v_reg;
  assign data_o[628] = data_o_628_sv2v_reg;
  assign data_o[627] = data_o_627_sv2v_reg;
  assign data_o[626] = data_o_626_sv2v_reg;
  assign data_o[625] = data_o_625_sv2v_reg;
  assign data_o[624] = data_o_624_sv2v_reg;
  assign data_o[623] = data_o_623_sv2v_reg;
  assign data_o[622] = data_o_622_sv2v_reg;
  assign data_o[621] = data_o_621_sv2v_reg;
  assign data_o[620] = data_o_620_sv2v_reg;
  assign data_o[619] = data_o_619_sv2v_reg;
  assign data_o[618] = data_o_618_sv2v_reg;
  assign data_o[617] = data_o_617_sv2v_reg;
  assign data_o[616] = data_o_616_sv2v_reg;
  assign data_o[615] = data_o_615_sv2v_reg;
  assign data_o[614] = data_o_614_sv2v_reg;
  assign data_o[613] = data_o_613_sv2v_reg;
  assign data_o[612] = data_o_612_sv2v_reg;
  assign data_o[611] = data_o_611_sv2v_reg;
  assign data_o[610] = data_o_610_sv2v_reg;
  assign data_o[609] = data_o_609_sv2v_reg;
  assign data_o[608] = data_o_608_sv2v_reg;
  assign data_o[607] = data_o_607_sv2v_reg;
  assign data_o[606] = data_o_606_sv2v_reg;
  assign data_o[605] = data_o_605_sv2v_reg;
  assign data_o[604] = data_o_604_sv2v_reg;
  assign data_o[603] = data_o_603_sv2v_reg;
  assign data_o[602] = data_o_602_sv2v_reg;
  assign data_o[601] = data_o_601_sv2v_reg;
  assign data_o[600] = data_o_600_sv2v_reg;
  assign data_o[599] = data_o_599_sv2v_reg;
  assign data_o[598] = data_o_598_sv2v_reg;
  assign data_o[597] = data_o_597_sv2v_reg;
  assign data_o[596] = data_o_596_sv2v_reg;
  assign data_o[595] = data_o_595_sv2v_reg;
  assign data_o[594] = data_o_594_sv2v_reg;
  assign data_o[593] = data_o_593_sv2v_reg;
  assign data_o[592] = data_o_592_sv2v_reg;
  assign data_o[591] = data_o_591_sv2v_reg;
  assign data_o[590] = data_o_590_sv2v_reg;
  assign data_o[589] = data_o_589_sv2v_reg;
  assign data_o[588] = data_o_588_sv2v_reg;
  assign data_o[587] = data_o_587_sv2v_reg;
  assign data_o[586] = data_o_586_sv2v_reg;
  assign data_o[585] = data_o_585_sv2v_reg;
  assign data_o[584] = data_o_584_sv2v_reg;
  assign data_o[583] = data_o_583_sv2v_reg;
  assign data_o[582] = data_o_582_sv2v_reg;
  assign data_o[581] = data_o_581_sv2v_reg;
  assign data_o[580] = data_o_580_sv2v_reg;
  assign data_o[579] = data_o_579_sv2v_reg;
  assign data_o[578] = data_o_578_sv2v_reg;
  assign data_o[577] = data_o_577_sv2v_reg;
  assign data_o[576] = data_o_576_sv2v_reg;
  assign data_o[575] = data_o_575_sv2v_reg;
  assign data_o[574] = data_o_574_sv2v_reg;
  assign data_o[573] = data_o_573_sv2v_reg;
  assign data_o[572] = data_o_572_sv2v_reg;
  assign data_o[571] = data_o_571_sv2v_reg;
  assign data_o[570] = data_o_570_sv2v_reg;
  assign data_o[569] = data_o_569_sv2v_reg;
  assign data_o[568] = data_o_568_sv2v_reg;
  assign data_o[567] = data_o_567_sv2v_reg;
  assign data_o[566] = data_o_566_sv2v_reg;
  assign data_o[565] = data_o_565_sv2v_reg;
  assign data_o[564] = data_o_564_sv2v_reg;
  assign data_o[563] = data_o_563_sv2v_reg;
  assign data_o[562] = data_o_562_sv2v_reg;
  assign data_o[561] = data_o_561_sv2v_reg;
  assign data_o[560] = data_o_560_sv2v_reg;
  assign data_o[559] = data_o_559_sv2v_reg;
  assign data_o[558] = data_o_558_sv2v_reg;
  assign data_o[557] = data_o_557_sv2v_reg;
  assign data_o[556] = data_o_556_sv2v_reg;
  assign data_o[555] = data_o_555_sv2v_reg;
  assign data_o[554] = data_o_554_sv2v_reg;
  assign data_o[553] = data_o_553_sv2v_reg;
  assign data_o[552] = data_o_552_sv2v_reg;
  assign data_o[551] = data_o_551_sv2v_reg;
  assign data_o[550] = data_o_550_sv2v_reg;
  assign data_o[549] = data_o_549_sv2v_reg;
  assign data_o[548] = data_o_548_sv2v_reg;
  assign data_o[547] = data_o_547_sv2v_reg;
  assign data_o[546] = data_o_546_sv2v_reg;
  assign data_o[545] = data_o_545_sv2v_reg;
  assign data_o[544] = data_o_544_sv2v_reg;
  assign data_o[543] = data_o_543_sv2v_reg;
  assign data_o[542] = data_o_542_sv2v_reg;
  assign data_o[541] = data_o_541_sv2v_reg;
  assign data_o[540] = data_o_540_sv2v_reg;
  assign data_o[539] = data_o_539_sv2v_reg;
  assign data_o[538] = data_o_538_sv2v_reg;
  assign data_o[537] = data_o_537_sv2v_reg;
  assign data_o[536] = data_o_536_sv2v_reg;
  assign data_o[535] = data_o_535_sv2v_reg;
  assign data_o[534] = data_o_534_sv2v_reg;
  assign data_o[533] = data_o_533_sv2v_reg;
  assign data_o[532] = data_o_532_sv2v_reg;
  assign data_o[531] = data_o_531_sv2v_reg;
  assign data_o[530] = data_o_530_sv2v_reg;
  assign data_o[529] = data_o_529_sv2v_reg;
  assign data_o[528] = data_o_528_sv2v_reg;
  assign data_o[527] = data_o_527_sv2v_reg;
  assign data_o[526] = data_o_526_sv2v_reg;
  assign data_o[525] = data_o_525_sv2v_reg;
  assign data_o[524] = data_o_524_sv2v_reg;
  assign data_o[523] = data_o_523_sv2v_reg;
  assign data_o[522] = data_o_522_sv2v_reg;
  assign data_o[521] = data_o_521_sv2v_reg;
  assign data_o[520] = data_o_520_sv2v_reg;
  assign data_o[519] = data_o_519_sv2v_reg;
  assign data_o[518] = data_o_518_sv2v_reg;
  assign data_o[517] = data_o_517_sv2v_reg;
  assign data_o[516] = data_o_516_sv2v_reg;
  assign data_o[515] = data_o_515_sv2v_reg;
  assign data_o[514] = data_o_514_sv2v_reg;
  assign data_o[513] = data_o_513_sv2v_reg;
  assign data_o[512] = data_o_512_sv2v_reg;
  assign data_o[511] = data_o_511_sv2v_reg;
  assign data_o[510] = data_o_510_sv2v_reg;
  assign data_o[509] = data_o_509_sv2v_reg;
  assign data_o[508] = data_o_508_sv2v_reg;
  assign data_o[507] = data_o_507_sv2v_reg;
  assign data_o[506] = data_o_506_sv2v_reg;
  assign data_o[505] = data_o_505_sv2v_reg;
  assign data_o[504] = data_o_504_sv2v_reg;
  assign data_o[503] = data_o_503_sv2v_reg;
  assign data_o[502] = data_o_502_sv2v_reg;
  assign data_o[501] = data_o_501_sv2v_reg;
  assign data_o[500] = data_o_500_sv2v_reg;
  assign data_o[499] = data_o_499_sv2v_reg;
  assign data_o[498] = data_o_498_sv2v_reg;
  assign data_o[497] = data_o_497_sv2v_reg;
  assign data_o[496] = data_o_496_sv2v_reg;
  assign data_o[495] = data_o_495_sv2v_reg;
  assign data_o[494] = data_o_494_sv2v_reg;
  assign data_o[493] = data_o_493_sv2v_reg;
  assign data_o[492] = data_o_492_sv2v_reg;
  assign data_o[491] = data_o_491_sv2v_reg;
  assign data_o[490] = data_o_490_sv2v_reg;
  assign data_o[489] = data_o_489_sv2v_reg;
  assign data_o[488] = data_o_488_sv2v_reg;
  assign data_o[487] = data_o_487_sv2v_reg;
  assign data_o[486] = data_o_486_sv2v_reg;
  assign data_o[485] = data_o_485_sv2v_reg;
  assign data_o[484] = data_o_484_sv2v_reg;
  assign data_o[483] = data_o_483_sv2v_reg;
  assign data_o[482] = data_o_482_sv2v_reg;
  assign data_o[481] = data_o_481_sv2v_reg;
  assign data_o[480] = data_o_480_sv2v_reg;
  assign data_o[479] = data_o_479_sv2v_reg;
  assign data_o[478] = data_o_478_sv2v_reg;
  assign data_o[477] = data_o_477_sv2v_reg;
  assign data_o[476] = data_o_476_sv2v_reg;
  assign data_o[475] = data_o_475_sv2v_reg;
  assign data_o[474] = data_o_474_sv2v_reg;
  assign data_o[473] = data_o_473_sv2v_reg;
  assign data_o[472] = data_o_472_sv2v_reg;
  assign data_o[471] = data_o_471_sv2v_reg;
  assign data_o[470] = data_o_470_sv2v_reg;
  assign data_o[469] = data_o_469_sv2v_reg;
  assign data_o[468] = data_o_468_sv2v_reg;
  assign data_o[467] = data_o_467_sv2v_reg;
  assign data_o[466] = data_o_466_sv2v_reg;
  assign data_o[465] = data_o_465_sv2v_reg;
  assign data_o[464] = data_o_464_sv2v_reg;
  assign data_o[463] = data_o_463_sv2v_reg;
  assign data_o[462] = data_o_462_sv2v_reg;
  assign data_o[461] = data_o_461_sv2v_reg;
  assign data_o[460] = data_o_460_sv2v_reg;
  assign data_o[459] = data_o_459_sv2v_reg;
  assign data_o[458] = data_o_458_sv2v_reg;
  assign data_o[457] = data_o_457_sv2v_reg;
  assign data_o[456] = data_o_456_sv2v_reg;
  assign data_o[455] = data_o_455_sv2v_reg;
  assign data_o[454] = data_o_454_sv2v_reg;
  assign data_o[453] = data_o_453_sv2v_reg;
  assign data_o[452] = data_o_452_sv2v_reg;
  assign data_o[451] = data_o_451_sv2v_reg;
  assign data_o[450] = data_o_450_sv2v_reg;
  assign data_o[449] = data_o_449_sv2v_reg;
  assign data_o[448] = data_o_448_sv2v_reg;
  assign data_o[447] = data_o_447_sv2v_reg;
  assign data_o[446] = data_o_446_sv2v_reg;
  assign data_o[445] = data_o_445_sv2v_reg;
  assign data_o[444] = data_o_444_sv2v_reg;
  assign data_o[443] = data_o_443_sv2v_reg;
  assign data_o[442] = data_o_442_sv2v_reg;
  assign data_o[441] = data_o_441_sv2v_reg;
  assign data_o[440] = data_o_440_sv2v_reg;
  assign data_o[439] = data_o_439_sv2v_reg;
  assign data_o[438] = data_o_438_sv2v_reg;
  assign data_o[437] = data_o_437_sv2v_reg;
  assign data_o[436] = data_o_436_sv2v_reg;
  assign data_o[435] = data_o_435_sv2v_reg;
  assign data_o[434] = data_o_434_sv2v_reg;
  assign data_o[433] = data_o_433_sv2v_reg;
  assign data_o[432] = data_o_432_sv2v_reg;
  assign data_o[431] = data_o_431_sv2v_reg;
  assign data_o[430] = data_o_430_sv2v_reg;
  assign data_o[429] = data_o_429_sv2v_reg;
  assign data_o[428] = data_o_428_sv2v_reg;
  assign data_o[427] = data_o_427_sv2v_reg;
  assign data_o[426] = data_o_426_sv2v_reg;
  assign data_o[425] = data_o_425_sv2v_reg;
  assign data_o[424] = data_o_424_sv2v_reg;
  assign data_o[423] = data_o_423_sv2v_reg;
  assign data_o[422] = data_o_422_sv2v_reg;
  assign data_o[421] = data_o_421_sv2v_reg;
  assign data_o[420] = data_o_420_sv2v_reg;
  assign data_o[419] = data_o_419_sv2v_reg;
  assign data_o[418] = data_o_418_sv2v_reg;
  assign data_o[417] = data_o_417_sv2v_reg;
  assign data_o[416] = data_o_416_sv2v_reg;
  assign data_o[415] = data_o_415_sv2v_reg;
  assign data_o[414] = data_o_414_sv2v_reg;
  assign data_o[413] = data_o_413_sv2v_reg;
  assign data_o[412] = data_o_412_sv2v_reg;
  assign data_o[411] = data_o_411_sv2v_reg;
  assign data_o[410] = data_o_410_sv2v_reg;
  assign data_o[409] = data_o_409_sv2v_reg;
  assign data_o[408] = data_o_408_sv2v_reg;
  assign data_o[407] = data_o_407_sv2v_reg;
  assign data_o[406] = data_o_406_sv2v_reg;
  assign data_o[405] = data_o_405_sv2v_reg;
  assign data_o[404] = data_o_404_sv2v_reg;
  assign data_o[403] = data_o_403_sv2v_reg;
  assign data_o[402] = data_o_402_sv2v_reg;
  assign data_o[401] = data_o_401_sv2v_reg;
  assign data_o[400] = data_o_400_sv2v_reg;
  assign data_o[399] = data_o_399_sv2v_reg;
  assign data_o[398] = data_o_398_sv2v_reg;
  assign data_o[397] = data_o_397_sv2v_reg;
  assign data_o[396] = data_o_396_sv2v_reg;
  assign data_o[395] = data_o_395_sv2v_reg;
  assign data_o[394] = data_o_394_sv2v_reg;
  assign data_o[393] = data_o_393_sv2v_reg;
  assign data_o[392] = data_o_392_sv2v_reg;
  assign data_o[391] = data_o_391_sv2v_reg;
  assign data_o[390] = data_o_390_sv2v_reg;
  assign data_o[389] = data_o_389_sv2v_reg;
  assign data_o[388] = data_o_388_sv2v_reg;
  assign data_o[387] = data_o_387_sv2v_reg;
  assign data_o[386] = data_o_386_sv2v_reg;
  assign data_o[385] = data_o_385_sv2v_reg;
  assign data_o[384] = data_o_384_sv2v_reg;
  assign data_o[383] = data_o_383_sv2v_reg;
  assign data_o[382] = data_o_382_sv2v_reg;
  assign data_o[381] = data_o_381_sv2v_reg;
  assign data_o[380] = data_o_380_sv2v_reg;
  assign data_o[379] = data_o_379_sv2v_reg;
  assign data_o[378] = data_o_378_sv2v_reg;
  assign data_o[377] = data_o_377_sv2v_reg;
  assign data_o[376] = data_o_376_sv2v_reg;
  assign data_o[375] = data_o_375_sv2v_reg;
  assign data_o[374] = data_o_374_sv2v_reg;
  assign data_o[373] = data_o_373_sv2v_reg;
  assign data_o[372] = data_o_372_sv2v_reg;
  assign data_o[371] = data_o_371_sv2v_reg;
  assign data_o[370] = data_o_370_sv2v_reg;
  assign data_o[369] = data_o_369_sv2v_reg;
  assign data_o[368] = data_o_368_sv2v_reg;
  assign data_o[367] = data_o_367_sv2v_reg;
  assign data_o[366] = data_o_366_sv2v_reg;
  assign data_o[365] = data_o_365_sv2v_reg;
  assign data_o[364] = data_o_364_sv2v_reg;
  assign data_o[363] = data_o_363_sv2v_reg;
  assign data_o[362] = data_o_362_sv2v_reg;
  assign data_o[361] = data_o_361_sv2v_reg;
  assign data_o[360] = data_o_360_sv2v_reg;
  assign data_o[359] = data_o_359_sv2v_reg;
  assign data_o[358] = data_o_358_sv2v_reg;
  assign data_o[357] = data_o_357_sv2v_reg;
  assign data_o[356] = data_o_356_sv2v_reg;
  assign data_o[355] = data_o_355_sv2v_reg;
  assign data_o[354] = data_o_354_sv2v_reg;
  assign data_o[353] = data_o_353_sv2v_reg;
  assign data_o[352] = data_o_352_sv2v_reg;
  assign data_o[351] = data_o_351_sv2v_reg;
  assign data_o[350] = data_o_350_sv2v_reg;
  assign data_o[349] = data_o_349_sv2v_reg;
  assign data_o[348] = data_o_348_sv2v_reg;
  assign data_o[347] = data_o_347_sv2v_reg;
  assign data_o[346] = data_o_346_sv2v_reg;
  assign data_o[345] = data_o_345_sv2v_reg;
  assign data_o[344] = data_o_344_sv2v_reg;
  assign data_o[343] = data_o_343_sv2v_reg;
  assign data_o[342] = data_o_342_sv2v_reg;
  assign data_o[341] = data_o_341_sv2v_reg;
  assign data_o[340] = data_o_340_sv2v_reg;
  assign data_o[339] = data_o_339_sv2v_reg;
  assign data_o[338] = data_o_338_sv2v_reg;
  assign data_o[337] = data_o_337_sv2v_reg;
  assign data_o[336] = data_o_336_sv2v_reg;
  assign data_o[335] = data_o_335_sv2v_reg;
  assign data_o[334] = data_o_334_sv2v_reg;
  assign data_o[333] = data_o_333_sv2v_reg;
  assign data_o[332] = data_o_332_sv2v_reg;
  assign data_o[331] = data_o_331_sv2v_reg;
  assign data_o[330] = data_o_330_sv2v_reg;
  assign data_o[329] = data_o_329_sv2v_reg;
  assign data_o[328] = data_o_328_sv2v_reg;
  assign data_o[327] = data_o_327_sv2v_reg;
  assign data_o[326] = data_o_326_sv2v_reg;
  assign data_o[325] = data_o_325_sv2v_reg;
  assign data_o[324] = data_o_324_sv2v_reg;
  assign data_o[323] = data_o_323_sv2v_reg;
  assign data_o[322] = data_o_322_sv2v_reg;
  assign data_o[321] = data_o_321_sv2v_reg;
  assign data_o[320] = data_o_320_sv2v_reg;
  assign data_o[319] = data_o_319_sv2v_reg;
  assign data_o[318] = data_o_318_sv2v_reg;
  assign data_o[317] = data_o_317_sv2v_reg;
  assign data_o[316] = data_o_316_sv2v_reg;
  assign data_o[315] = data_o_315_sv2v_reg;
  assign data_o[314] = data_o_314_sv2v_reg;
  assign data_o[313] = data_o_313_sv2v_reg;
  assign data_o[312] = data_o_312_sv2v_reg;
  assign data_o[311] = data_o_311_sv2v_reg;
  assign data_o[310] = data_o_310_sv2v_reg;
  assign data_o[309] = data_o_309_sv2v_reg;
  assign data_o[308] = data_o_308_sv2v_reg;
  assign data_o[307] = data_o_307_sv2v_reg;
  assign data_o[306] = data_o_306_sv2v_reg;
  assign data_o[305] = data_o_305_sv2v_reg;
  assign data_o[304] = data_o_304_sv2v_reg;
  assign data_o[303] = data_o_303_sv2v_reg;
  assign data_o[302] = data_o_302_sv2v_reg;
  assign data_o[301] = data_o_301_sv2v_reg;
  assign data_o[300] = data_o_300_sv2v_reg;
  assign data_o[299] = data_o_299_sv2v_reg;
  assign data_o[298] = data_o_298_sv2v_reg;
  assign data_o[297] = data_o_297_sv2v_reg;
  assign data_o[296] = data_o_296_sv2v_reg;
  assign data_o[295] = data_o_295_sv2v_reg;
  assign data_o[294] = data_o_294_sv2v_reg;
  assign data_o[293] = data_o_293_sv2v_reg;
  assign data_o[292] = data_o_292_sv2v_reg;
  assign data_o[291] = data_o_291_sv2v_reg;
  assign data_o[290] = data_o_290_sv2v_reg;
  assign data_o[289] = data_o_289_sv2v_reg;
  assign data_o[288] = data_o_288_sv2v_reg;
  assign data_o[287] = data_o_287_sv2v_reg;
  assign data_o[286] = data_o_286_sv2v_reg;
  assign data_o[285] = data_o_285_sv2v_reg;
  assign data_o[284] = data_o_284_sv2v_reg;
  assign data_o[283] = data_o_283_sv2v_reg;
  assign data_o[282] = data_o_282_sv2v_reg;
  assign data_o[281] = data_o_281_sv2v_reg;
  assign data_o[280] = data_o_280_sv2v_reg;
  assign data_o[279] = data_o_279_sv2v_reg;
  assign data_o[278] = data_o_278_sv2v_reg;
  assign data_o[277] = data_o_277_sv2v_reg;
  assign data_o[276] = data_o_276_sv2v_reg;
  assign data_o[275] = data_o_275_sv2v_reg;
  assign data_o[274] = data_o_274_sv2v_reg;
  assign data_o[273] = data_o_273_sv2v_reg;
  assign data_o[272] = data_o_272_sv2v_reg;
  assign data_o[271] = data_o_271_sv2v_reg;
  assign data_o[270] = data_o_270_sv2v_reg;
  assign data_o[269] = data_o_269_sv2v_reg;
  assign data_o[268] = data_o_268_sv2v_reg;
  assign data_o[267] = data_o_267_sv2v_reg;
  assign data_o[266] = data_o_266_sv2v_reg;
  assign data_o[265] = data_o_265_sv2v_reg;
  assign data_o[264] = data_o_264_sv2v_reg;
  assign data_o[263] = data_o_263_sv2v_reg;
  assign data_o[262] = data_o_262_sv2v_reg;
  assign data_o[261] = data_o_261_sv2v_reg;
  assign data_o[260] = data_o_260_sv2v_reg;
  assign data_o[259] = data_o_259_sv2v_reg;
  assign data_o[258] = data_o_258_sv2v_reg;
  assign data_o[257] = data_o_257_sv2v_reg;
  assign data_o[256] = data_o_256_sv2v_reg;
  assign data_o[255] = data_o_255_sv2v_reg;
  assign data_o[254] = data_o_254_sv2v_reg;
  assign data_o[253] = data_o_253_sv2v_reg;
  assign data_o[252] = data_o_252_sv2v_reg;
  assign data_o[251] = data_o_251_sv2v_reg;
  assign data_o[250] = data_o_250_sv2v_reg;
  assign data_o[249] = data_o_249_sv2v_reg;
  assign data_o[248] = data_o_248_sv2v_reg;
  assign data_o[247] = data_o_247_sv2v_reg;
  assign data_o[246] = data_o_246_sv2v_reg;
  assign data_o[245] = data_o_245_sv2v_reg;
  assign data_o[244] = data_o_244_sv2v_reg;
  assign data_o[243] = data_o_243_sv2v_reg;
  assign data_o[242] = data_o_242_sv2v_reg;
  assign data_o[241] = data_o_241_sv2v_reg;
  assign data_o[240] = data_o_240_sv2v_reg;
  assign data_o[239] = data_o_239_sv2v_reg;
  assign data_o[238] = data_o_238_sv2v_reg;
  assign data_o[237] = data_o_237_sv2v_reg;
  assign data_o[236] = data_o_236_sv2v_reg;
  assign data_o[235] = data_o_235_sv2v_reg;
  assign data_o[234] = data_o_234_sv2v_reg;
  assign data_o[233] = data_o_233_sv2v_reg;
  assign data_o[232] = data_o_232_sv2v_reg;
  assign data_o[231] = data_o_231_sv2v_reg;
  assign data_o[230] = data_o_230_sv2v_reg;
  assign data_o[229] = data_o_229_sv2v_reg;
  assign data_o[228] = data_o_228_sv2v_reg;
  assign data_o[227] = data_o_227_sv2v_reg;
  assign data_o[226] = data_o_226_sv2v_reg;
  assign data_o[225] = data_o_225_sv2v_reg;
  assign data_o[224] = data_o_224_sv2v_reg;
  assign data_o[223] = data_o_223_sv2v_reg;
  assign data_o[222] = data_o_222_sv2v_reg;
  assign data_o[221] = data_o_221_sv2v_reg;
  assign data_o[220] = data_o_220_sv2v_reg;
  assign data_o[219] = data_o_219_sv2v_reg;
  assign data_o[218] = data_o_218_sv2v_reg;
  assign data_o[217] = data_o_217_sv2v_reg;
  assign data_o[216] = data_o_216_sv2v_reg;
  assign data_o[215] = data_o_215_sv2v_reg;
  assign data_o[214] = data_o_214_sv2v_reg;
  assign data_o[213] = data_o_213_sv2v_reg;
  assign data_o[212] = data_o_212_sv2v_reg;
  assign data_o[211] = data_o_211_sv2v_reg;
  assign data_o[210] = data_o_210_sv2v_reg;
  assign data_o[209] = data_o_209_sv2v_reg;
  assign data_o[208] = data_o_208_sv2v_reg;
  assign data_o[207] = data_o_207_sv2v_reg;
  assign data_o[206] = data_o_206_sv2v_reg;
  assign data_o[205] = data_o_205_sv2v_reg;
  assign data_o[204] = data_o_204_sv2v_reg;
  assign data_o[203] = data_o_203_sv2v_reg;
  assign data_o[202] = data_o_202_sv2v_reg;
  assign data_o[201] = data_o_201_sv2v_reg;
  assign data_o[200] = data_o_200_sv2v_reg;
  assign data_o[199] = data_o_199_sv2v_reg;
  assign data_o[198] = data_o_198_sv2v_reg;
  assign data_o[197] = data_o_197_sv2v_reg;
  assign data_o[196] = data_o_196_sv2v_reg;
  assign data_o[195] = data_o_195_sv2v_reg;
  assign data_o[194] = data_o_194_sv2v_reg;
  assign data_o[193] = data_o_193_sv2v_reg;
  assign data_o[192] = data_o_192_sv2v_reg;
  assign data_o[191] = data_o_191_sv2v_reg;
  assign data_o[190] = data_o_190_sv2v_reg;
  assign data_o[189] = data_o_189_sv2v_reg;
  assign data_o[188] = data_o_188_sv2v_reg;
  assign data_o[187] = data_o_187_sv2v_reg;
  assign data_o[186] = data_o_186_sv2v_reg;
  assign data_o[185] = data_o_185_sv2v_reg;
  assign data_o[184] = data_o_184_sv2v_reg;
  assign data_o[183] = data_o_183_sv2v_reg;
  assign data_o[182] = data_o_182_sv2v_reg;
  assign data_o[181] = data_o_181_sv2v_reg;
  assign data_o[180] = data_o_180_sv2v_reg;
  assign data_o[179] = data_o_179_sv2v_reg;
  assign data_o[178] = data_o_178_sv2v_reg;
  assign data_o[177] = data_o_177_sv2v_reg;
  assign data_o[176] = data_o_176_sv2v_reg;
  assign data_o[175] = data_o_175_sv2v_reg;
  assign data_o[174] = data_o_174_sv2v_reg;
  assign data_o[173] = data_o_173_sv2v_reg;
  assign data_o[172] = data_o_172_sv2v_reg;
  assign data_o[171] = data_o_171_sv2v_reg;
  assign data_o[170] = data_o_170_sv2v_reg;
  assign data_o[169] = data_o_169_sv2v_reg;
  assign data_o[168] = data_o_168_sv2v_reg;
  assign data_o[167] = data_o_167_sv2v_reg;
  assign data_o[166] = data_o_166_sv2v_reg;
  assign data_o[165] = data_o_165_sv2v_reg;
  assign data_o[164] = data_o_164_sv2v_reg;
  assign data_o[163] = data_o_163_sv2v_reg;
  assign data_o[162] = data_o_162_sv2v_reg;
  assign data_o[161] = data_o_161_sv2v_reg;
  assign data_o[160] = data_o_160_sv2v_reg;
  assign data_o[159] = data_o_159_sv2v_reg;
  assign data_o[158] = data_o_158_sv2v_reg;
  assign data_o[157] = data_o_157_sv2v_reg;
  assign data_o[156] = data_o_156_sv2v_reg;
  assign data_o[155] = data_o_155_sv2v_reg;
  assign data_o[154] = data_o_154_sv2v_reg;
  assign data_o[153] = data_o_153_sv2v_reg;
  assign data_o[152] = data_o_152_sv2v_reg;
  assign data_o[151] = data_o_151_sv2v_reg;
  assign data_o[150] = data_o_150_sv2v_reg;
  assign data_o[149] = data_o_149_sv2v_reg;
  assign data_o[148] = data_o_148_sv2v_reg;
  assign data_o[147] = data_o_147_sv2v_reg;
  assign data_o[146] = data_o_146_sv2v_reg;
  assign data_o[145] = data_o_145_sv2v_reg;
  assign data_o[144] = data_o_144_sv2v_reg;
  assign data_o[143] = data_o_143_sv2v_reg;
  assign data_o[142] = data_o_142_sv2v_reg;
  assign data_o[141] = data_o_141_sv2v_reg;
  assign data_o[140] = data_o_140_sv2v_reg;
  assign data_o[139] = data_o_139_sv2v_reg;
  assign data_o[138] = data_o_138_sv2v_reg;
  assign data_o[137] = data_o_137_sv2v_reg;
  assign data_o[136] = data_o_136_sv2v_reg;
  assign data_o[135] = data_o_135_sv2v_reg;
  assign data_o[134] = data_o_134_sv2v_reg;
  assign data_o[133] = data_o_133_sv2v_reg;
  assign data_o[132] = data_o_132_sv2v_reg;
  assign data_o[131] = data_o_131_sv2v_reg;
  assign data_o[130] = data_o_130_sv2v_reg;
  assign data_o[129] = data_o_129_sv2v_reg;
  assign data_o[128] = data_o_128_sv2v_reg;
  assign data_o[127] = data_o_127_sv2v_reg;
  assign data_o[126] = data_o_126_sv2v_reg;
  assign data_o[125] = data_o_125_sv2v_reg;
  assign data_o[124] = data_o_124_sv2v_reg;
  assign data_o[123] = data_o_123_sv2v_reg;
  assign data_o[122] = data_o_122_sv2v_reg;
  assign data_o[121] = data_o_121_sv2v_reg;
  assign data_o[120] = data_o_120_sv2v_reg;
  assign data_o[119] = data_o_119_sv2v_reg;
  assign data_o[118] = data_o_118_sv2v_reg;
  assign data_o[117] = data_o_117_sv2v_reg;
  assign data_o[116] = data_o_116_sv2v_reg;
  assign data_o[115] = data_o_115_sv2v_reg;
  assign data_o[114] = data_o_114_sv2v_reg;
  assign data_o[113] = data_o_113_sv2v_reg;
  assign data_o[112] = data_o_112_sv2v_reg;
  assign data_o[111] = data_o_111_sv2v_reg;
  assign data_o[110] = data_o_110_sv2v_reg;
  assign data_o[109] = data_o_109_sv2v_reg;
  assign data_o[108] = data_o_108_sv2v_reg;
  assign data_o[107] = data_o_107_sv2v_reg;
  assign data_o[106] = data_o_106_sv2v_reg;
  assign data_o[105] = data_o_105_sv2v_reg;
  assign data_o[104] = data_o_104_sv2v_reg;
  assign data_o[103] = data_o_103_sv2v_reg;
  assign data_o[102] = data_o_102_sv2v_reg;
  assign data_o[101] = data_o_101_sv2v_reg;
  assign data_o[100] = data_o_100_sv2v_reg;
  assign data_o[99] = data_o_99_sv2v_reg;
  assign data_o[98] = data_o_98_sv2v_reg;
  assign data_o[97] = data_o_97_sv2v_reg;
  assign data_o[96] = data_o_96_sv2v_reg;
  assign data_o[95] = data_o_95_sv2v_reg;
  assign data_o[94] = data_o_94_sv2v_reg;
  assign data_o[93] = data_o_93_sv2v_reg;
  assign data_o[92] = data_o_92_sv2v_reg;
  assign data_o[91] = data_o_91_sv2v_reg;
  assign data_o[90] = data_o_90_sv2v_reg;
  assign data_o[89] = data_o_89_sv2v_reg;
  assign data_o[88] = data_o_88_sv2v_reg;
  assign data_o[87] = data_o_87_sv2v_reg;
  assign data_o[86] = data_o_86_sv2v_reg;
  assign data_o[85] = data_o_85_sv2v_reg;
  assign data_o[84] = data_o_84_sv2v_reg;
  assign data_o[83] = data_o_83_sv2v_reg;
  assign data_o[82] = data_o_82_sv2v_reg;
  assign data_o[81] = data_o_81_sv2v_reg;
  assign data_o[80] = data_o_80_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_682_sv2v_reg <= data_i[682];
      data_o_681_sv2v_reg <= data_i[681];
      data_o_680_sv2v_reg <= data_i[680];
      data_o_679_sv2v_reg <= data_i[679];
      data_o_678_sv2v_reg <= data_i[678];
      data_o_677_sv2v_reg <= data_i[677];
      data_o_676_sv2v_reg <= data_i[676];
      data_o_675_sv2v_reg <= data_i[675];
      data_o_674_sv2v_reg <= data_i[674];
      data_o_673_sv2v_reg <= data_i[673];
      data_o_672_sv2v_reg <= data_i[672];
      data_o_671_sv2v_reg <= data_i[671];
      data_o_670_sv2v_reg <= data_i[670];
      data_o_669_sv2v_reg <= data_i[669];
      data_o_668_sv2v_reg <= data_i[668];
      data_o_667_sv2v_reg <= data_i[667];
      data_o_666_sv2v_reg <= data_i[666];
      data_o_665_sv2v_reg <= data_i[665];
      data_o_664_sv2v_reg <= data_i[664];
      data_o_663_sv2v_reg <= data_i[663];
      data_o_662_sv2v_reg <= data_i[662];
      data_o_661_sv2v_reg <= data_i[661];
      data_o_660_sv2v_reg <= data_i[660];
      data_o_659_sv2v_reg <= data_i[659];
      data_o_658_sv2v_reg <= data_i[658];
      data_o_657_sv2v_reg <= data_i[657];
      data_o_656_sv2v_reg <= data_i[656];
      data_o_655_sv2v_reg <= data_i[655];
      data_o_654_sv2v_reg <= data_i[654];
      data_o_653_sv2v_reg <= data_i[653];
      data_o_652_sv2v_reg <= data_i[652];
      data_o_651_sv2v_reg <= data_i[651];
      data_o_650_sv2v_reg <= data_i[650];
      data_o_649_sv2v_reg <= data_i[649];
      data_o_648_sv2v_reg <= data_i[648];
      data_o_647_sv2v_reg <= data_i[647];
      data_o_646_sv2v_reg <= data_i[646];
      data_o_645_sv2v_reg <= data_i[645];
      data_o_644_sv2v_reg <= data_i[644];
      data_o_643_sv2v_reg <= data_i[643];
      data_o_642_sv2v_reg <= data_i[642];
      data_o_641_sv2v_reg <= data_i[641];
      data_o_640_sv2v_reg <= data_i[640];
      data_o_639_sv2v_reg <= data_i[639];
      data_o_638_sv2v_reg <= data_i[638];
      data_o_637_sv2v_reg <= data_i[637];
      data_o_636_sv2v_reg <= data_i[636];
      data_o_635_sv2v_reg <= data_i[635];
      data_o_634_sv2v_reg <= data_i[634];
      data_o_633_sv2v_reg <= data_i[633];
      data_o_632_sv2v_reg <= data_i[632];
      data_o_631_sv2v_reg <= data_i[631];
      data_o_630_sv2v_reg <= data_i[630];
      data_o_629_sv2v_reg <= data_i[629];
      data_o_628_sv2v_reg <= data_i[628];
      data_o_627_sv2v_reg <= data_i[627];
      data_o_626_sv2v_reg <= data_i[626];
      data_o_625_sv2v_reg <= data_i[625];
      data_o_624_sv2v_reg <= data_i[624];
      data_o_623_sv2v_reg <= data_i[623];
      data_o_622_sv2v_reg <= data_i[622];
      data_o_621_sv2v_reg <= data_i[621];
      data_o_620_sv2v_reg <= data_i[620];
      data_o_619_sv2v_reg <= data_i[619];
      data_o_618_sv2v_reg <= data_i[618];
      data_o_617_sv2v_reg <= data_i[617];
      data_o_616_sv2v_reg <= data_i[616];
      data_o_615_sv2v_reg <= data_i[615];
      data_o_614_sv2v_reg <= data_i[614];
      data_o_613_sv2v_reg <= data_i[613];
      data_o_612_sv2v_reg <= data_i[612];
      data_o_611_sv2v_reg <= data_i[611];
      data_o_610_sv2v_reg <= data_i[610];
      data_o_609_sv2v_reg <= data_i[609];
      data_o_608_sv2v_reg <= data_i[608];
      data_o_607_sv2v_reg <= data_i[607];
      data_o_606_sv2v_reg <= data_i[606];
      data_o_605_sv2v_reg <= data_i[605];
      data_o_604_sv2v_reg <= data_i[604];
      data_o_603_sv2v_reg <= data_i[603];
      data_o_602_sv2v_reg <= data_i[602];
      data_o_601_sv2v_reg <= data_i[601];
      data_o_600_sv2v_reg <= data_i[600];
      data_o_599_sv2v_reg <= data_i[599];
      data_o_598_sv2v_reg <= data_i[598];
      data_o_597_sv2v_reg <= data_i[597];
      data_o_596_sv2v_reg <= data_i[596];
      data_o_595_sv2v_reg <= data_i[595];
      data_o_594_sv2v_reg <= data_i[594];
      data_o_593_sv2v_reg <= data_i[593];
      data_o_592_sv2v_reg <= data_i[592];
      data_o_591_sv2v_reg <= data_i[591];
      data_o_590_sv2v_reg <= data_i[590];
      data_o_589_sv2v_reg <= data_i[589];
      data_o_588_sv2v_reg <= data_i[588];
      data_o_587_sv2v_reg <= data_i[587];
      data_o_586_sv2v_reg <= data_i[586];
      data_o_585_sv2v_reg <= data_i[585];
      data_o_584_sv2v_reg <= data_i[584];
      data_o_583_sv2v_reg <= data_i[583];
      data_o_582_sv2v_reg <= data_i[582];
      data_o_581_sv2v_reg <= data_i[581];
      data_o_580_sv2v_reg <= data_i[580];
      data_o_579_sv2v_reg <= data_i[579];
      data_o_578_sv2v_reg <= data_i[578];
      data_o_577_sv2v_reg <= data_i[577];
      data_o_576_sv2v_reg <= data_i[576];
      data_o_575_sv2v_reg <= data_i[575];
      data_o_574_sv2v_reg <= data_i[574];
      data_o_573_sv2v_reg <= data_i[573];
      data_o_572_sv2v_reg <= data_i[572];
      data_o_571_sv2v_reg <= data_i[571];
      data_o_570_sv2v_reg <= data_i[570];
      data_o_569_sv2v_reg <= data_i[569];
      data_o_568_sv2v_reg <= data_i[568];
      data_o_567_sv2v_reg <= data_i[567];
      data_o_566_sv2v_reg <= data_i[566];
      data_o_565_sv2v_reg <= data_i[565];
      data_o_564_sv2v_reg <= data_i[564];
      data_o_563_sv2v_reg <= data_i[563];
      data_o_562_sv2v_reg <= data_i[562];
      data_o_561_sv2v_reg <= data_i[561];
      data_o_560_sv2v_reg <= data_i[560];
      data_o_559_sv2v_reg <= data_i[559];
      data_o_558_sv2v_reg <= data_i[558];
      data_o_557_sv2v_reg <= data_i[557];
      data_o_556_sv2v_reg <= data_i[556];
      data_o_555_sv2v_reg <= data_i[555];
      data_o_554_sv2v_reg <= data_i[554];
      data_o_553_sv2v_reg <= data_i[553];
      data_o_552_sv2v_reg <= data_i[552];
      data_o_551_sv2v_reg <= data_i[551];
      data_o_550_sv2v_reg <= data_i[550];
      data_o_549_sv2v_reg <= data_i[549];
      data_o_548_sv2v_reg <= data_i[548];
      data_o_547_sv2v_reg <= data_i[547];
      data_o_546_sv2v_reg <= data_i[546];
      data_o_545_sv2v_reg <= data_i[545];
      data_o_544_sv2v_reg <= data_i[544];
      data_o_543_sv2v_reg <= data_i[543];
      data_o_542_sv2v_reg <= data_i[542];
      data_o_541_sv2v_reg <= data_i[541];
      data_o_540_sv2v_reg <= data_i[540];
      data_o_539_sv2v_reg <= data_i[539];
      data_o_538_sv2v_reg <= data_i[538];
      data_o_537_sv2v_reg <= data_i[537];
      data_o_536_sv2v_reg <= data_i[536];
      data_o_535_sv2v_reg <= data_i[535];
      data_o_534_sv2v_reg <= data_i[534];
      data_o_533_sv2v_reg <= data_i[533];
      data_o_532_sv2v_reg <= data_i[532];
      data_o_531_sv2v_reg <= data_i[531];
      data_o_530_sv2v_reg <= data_i[530];
      data_o_529_sv2v_reg <= data_i[529];
      data_o_528_sv2v_reg <= data_i[528];
      data_o_527_sv2v_reg <= data_i[527];
      data_o_526_sv2v_reg <= data_i[526];
      data_o_525_sv2v_reg <= data_i[525];
      data_o_524_sv2v_reg <= data_i[524];
      data_o_523_sv2v_reg <= data_i[523];
      data_o_522_sv2v_reg <= data_i[522];
      data_o_521_sv2v_reg <= data_i[521];
      data_o_520_sv2v_reg <= data_i[520];
      data_o_519_sv2v_reg <= data_i[519];
      data_o_518_sv2v_reg <= data_i[518];
      data_o_517_sv2v_reg <= data_i[517];
      data_o_516_sv2v_reg <= data_i[516];
      data_o_515_sv2v_reg <= data_i[515];
      data_o_514_sv2v_reg <= data_i[514];
      data_o_513_sv2v_reg <= data_i[513];
      data_o_512_sv2v_reg <= data_i[512];
      data_o_511_sv2v_reg <= data_i[511];
      data_o_510_sv2v_reg <= data_i[510];
      data_o_509_sv2v_reg <= data_i[509];
      data_o_508_sv2v_reg <= data_i[508];
      data_o_507_sv2v_reg <= data_i[507];
      data_o_506_sv2v_reg <= data_i[506];
      data_o_505_sv2v_reg <= data_i[505];
      data_o_504_sv2v_reg <= data_i[504];
      data_o_503_sv2v_reg <= data_i[503];
      data_o_502_sv2v_reg <= data_i[502];
      data_o_501_sv2v_reg <= data_i[501];
      data_o_500_sv2v_reg <= data_i[500];
      data_o_499_sv2v_reg <= data_i[499];
      data_o_498_sv2v_reg <= data_i[498];
      data_o_497_sv2v_reg <= data_i[497];
      data_o_496_sv2v_reg <= data_i[496];
      data_o_495_sv2v_reg <= data_i[495];
      data_o_494_sv2v_reg <= data_i[494];
      data_o_493_sv2v_reg <= data_i[493];
      data_o_492_sv2v_reg <= data_i[492];
      data_o_491_sv2v_reg <= data_i[491];
      data_o_490_sv2v_reg <= data_i[490];
      data_o_489_sv2v_reg <= data_i[489];
      data_o_488_sv2v_reg <= data_i[488];
      data_o_487_sv2v_reg <= data_i[487];
      data_o_486_sv2v_reg <= data_i[486];
      data_o_485_sv2v_reg <= data_i[485];
      data_o_484_sv2v_reg <= data_i[484];
      data_o_483_sv2v_reg <= data_i[483];
      data_o_482_sv2v_reg <= data_i[482];
      data_o_481_sv2v_reg <= data_i[481];
      data_o_480_sv2v_reg <= data_i[480];
      data_o_479_sv2v_reg <= data_i[479];
      data_o_478_sv2v_reg <= data_i[478];
      data_o_477_sv2v_reg <= data_i[477];
      data_o_476_sv2v_reg <= data_i[476];
      data_o_475_sv2v_reg <= data_i[475];
      data_o_474_sv2v_reg <= data_i[474];
      data_o_473_sv2v_reg <= data_i[473];
      data_o_472_sv2v_reg <= data_i[472];
      data_o_471_sv2v_reg <= data_i[471];
      data_o_470_sv2v_reg <= data_i[470];
      data_o_469_sv2v_reg <= data_i[469];
      data_o_468_sv2v_reg <= data_i[468];
      data_o_467_sv2v_reg <= data_i[467];
      data_o_466_sv2v_reg <= data_i[466];
      data_o_465_sv2v_reg <= data_i[465];
      data_o_464_sv2v_reg <= data_i[464];
      data_o_463_sv2v_reg <= data_i[463];
      data_o_462_sv2v_reg <= data_i[462];
      data_o_461_sv2v_reg <= data_i[461];
      data_o_460_sv2v_reg <= data_i[460];
      data_o_459_sv2v_reg <= data_i[459];
      data_o_458_sv2v_reg <= data_i[458];
      data_o_457_sv2v_reg <= data_i[457];
      data_o_456_sv2v_reg <= data_i[456];
      data_o_455_sv2v_reg <= data_i[455];
      data_o_454_sv2v_reg <= data_i[454];
      data_o_453_sv2v_reg <= data_i[453];
      data_o_452_sv2v_reg <= data_i[452];
      data_o_451_sv2v_reg <= data_i[451];
      data_o_450_sv2v_reg <= data_i[450];
      data_o_449_sv2v_reg <= data_i[449];
      data_o_448_sv2v_reg <= data_i[448];
      data_o_447_sv2v_reg <= data_i[447];
      data_o_446_sv2v_reg <= data_i[446];
      data_o_445_sv2v_reg <= data_i[445];
      data_o_444_sv2v_reg <= data_i[444];
      data_o_443_sv2v_reg <= data_i[443];
      data_o_442_sv2v_reg <= data_i[442];
      data_o_441_sv2v_reg <= data_i[441];
      data_o_440_sv2v_reg <= data_i[440];
      data_o_439_sv2v_reg <= data_i[439];
      data_o_438_sv2v_reg <= data_i[438];
      data_o_437_sv2v_reg <= data_i[437];
      data_o_436_sv2v_reg <= data_i[436];
      data_o_435_sv2v_reg <= data_i[435];
      data_o_434_sv2v_reg <= data_i[434];
      data_o_433_sv2v_reg <= data_i[433];
      data_o_432_sv2v_reg <= data_i[432];
      data_o_431_sv2v_reg <= data_i[431];
      data_o_430_sv2v_reg <= data_i[430];
      data_o_429_sv2v_reg <= data_i[429];
      data_o_428_sv2v_reg <= data_i[428];
      data_o_427_sv2v_reg <= data_i[427];
      data_o_426_sv2v_reg <= data_i[426];
      data_o_425_sv2v_reg <= data_i[425];
      data_o_424_sv2v_reg <= data_i[424];
      data_o_423_sv2v_reg <= data_i[423];
      data_o_422_sv2v_reg <= data_i[422];
      data_o_421_sv2v_reg <= data_i[421];
      data_o_420_sv2v_reg <= data_i[420];
      data_o_419_sv2v_reg <= data_i[419];
      data_o_418_sv2v_reg <= data_i[418];
      data_o_417_sv2v_reg <= data_i[417];
      data_o_416_sv2v_reg <= data_i[416];
      data_o_415_sv2v_reg <= data_i[415];
      data_o_414_sv2v_reg <= data_i[414];
      data_o_413_sv2v_reg <= data_i[413];
      data_o_412_sv2v_reg <= data_i[412];
      data_o_411_sv2v_reg <= data_i[411];
      data_o_410_sv2v_reg <= data_i[410];
      data_o_409_sv2v_reg <= data_i[409];
      data_o_408_sv2v_reg <= data_i[408];
      data_o_407_sv2v_reg <= data_i[407];
      data_o_406_sv2v_reg <= data_i[406];
      data_o_405_sv2v_reg <= data_i[405];
      data_o_404_sv2v_reg <= data_i[404];
      data_o_403_sv2v_reg <= data_i[403];
      data_o_402_sv2v_reg <= data_i[402];
      data_o_401_sv2v_reg <= data_i[401];
      data_o_400_sv2v_reg <= data_i[400];
      data_o_399_sv2v_reg <= data_i[399];
      data_o_398_sv2v_reg <= data_i[398];
      data_o_397_sv2v_reg <= data_i[397];
      data_o_396_sv2v_reg <= data_i[396];
      data_o_395_sv2v_reg <= data_i[395];
      data_o_394_sv2v_reg <= data_i[394];
      data_o_393_sv2v_reg <= data_i[393];
      data_o_392_sv2v_reg <= data_i[392];
      data_o_391_sv2v_reg <= data_i[391];
      data_o_390_sv2v_reg <= data_i[390];
      data_o_389_sv2v_reg <= data_i[389];
      data_o_388_sv2v_reg <= data_i[388];
      data_o_387_sv2v_reg <= data_i[387];
      data_o_386_sv2v_reg <= data_i[386];
      data_o_385_sv2v_reg <= data_i[385];
      data_o_384_sv2v_reg <= data_i[384];
      data_o_383_sv2v_reg <= data_i[383];
      data_o_382_sv2v_reg <= data_i[382];
      data_o_381_sv2v_reg <= data_i[381];
      data_o_380_sv2v_reg <= data_i[380];
      data_o_379_sv2v_reg <= data_i[379];
      data_o_378_sv2v_reg <= data_i[378];
      data_o_377_sv2v_reg <= data_i[377];
      data_o_376_sv2v_reg <= data_i[376];
      data_o_375_sv2v_reg <= data_i[375];
      data_o_374_sv2v_reg <= data_i[374];
      data_o_373_sv2v_reg <= data_i[373];
      data_o_372_sv2v_reg <= data_i[372];
      data_o_371_sv2v_reg <= data_i[371];
      data_o_370_sv2v_reg <= data_i[370];
      data_o_369_sv2v_reg <= data_i[369];
      data_o_368_sv2v_reg <= data_i[368];
      data_o_367_sv2v_reg <= data_i[367];
      data_o_366_sv2v_reg <= data_i[366];
      data_o_365_sv2v_reg <= data_i[365];
      data_o_364_sv2v_reg <= data_i[364];
      data_o_363_sv2v_reg <= data_i[363];
      data_o_362_sv2v_reg <= data_i[362];
      data_o_361_sv2v_reg <= data_i[361];
      data_o_360_sv2v_reg <= data_i[360];
      data_o_359_sv2v_reg <= data_i[359];
      data_o_358_sv2v_reg <= data_i[358];
      data_o_357_sv2v_reg <= data_i[357];
      data_o_356_sv2v_reg <= data_i[356];
      data_o_355_sv2v_reg <= data_i[355];
      data_o_354_sv2v_reg <= data_i[354];
      data_o_353_sv2v_reg <= data_i[353];
      data_o_352_sv2v_reg <= data_i[352];
      data_o_351_sv2v_reg <= data_i[351];
      data_o_350_sv2v_reg <= data_i[350];
      data_o_349_sv2v_reg <= data_i[349];
      data_o_348_sv2v_reg <= data_i[348];
      data_o_347_sv2v_reg <= data_i[347];
      data_o_346_sv2v_reg <= data_i[346];
      data_o_345_sv2v_reg <= data_i[345];
      data_o_344_sv2v_reg <= data_i[344];
      data_o_343_sv2v_reg <= data_i[343];
      data_o_342_sv2v_reg <= data_i[342];
      data_o_341_sv2v_reg <= data_i[341];
      data_o_340_sv2v_reg <= data_i[340];
      data_o_339_sv2v_reg <= data_i[339];
      data_o_338_sv2v_reg <= data_i[338];
      data_o_337_sv2v_reg <= data_i[337];
      data_o_336_sv2v_reg <= data_i[336];
      data_o_335_sv2v_reg <= data_i[335];
      data_o_334_sv2v_reg <= data_i[334];
      data_o_333_sv2v_reg <= data_i[333];
      data_o_332_sv2v_reg <= data_i[332];
      data_o_331_sv2v_reg <= data_i[331];
      data_o_330_sv2v_reg <= data_i[330];
      data_o_329_sv2v_reg <= data_i[329];
      data_o_328_sv2v_reg <= data_i[328];
      data_o_327_sv2v_reg <= data_i[327];
      data_o_326_sv2v_reg <= data_i[326];
      data_o_325_sv2v_reg <= data_i[325];
      data_o_324_sv2v_reg <= data_i[324];
      data_o_323_sv2v_reg <= data_i[323];
      data_o_322_sv2v_reg <= data_i[322];
      data_o_321_sv2v_reg <= data_i[321];
      data_o_320_sv2v_reg <= data_i[320];
      data_o_319_sv2v_reg <= data_i[319];
      data_o_318_sv2v_reg <= data_i[318];
      data_o_317_sv2v_reg <= data_i[317];
      data_o_316_sv2v_reg <= data_i[316];
      data_o_315_sv2v_reg <= data_i[315];
      data_o_314_sv2v_reg <= data_i[314];
      data_o_313_sv2v_reg <= data_i[313];
      data_o_312_sv2v_reg <= data_i[312];
      data_o_311_sv2v_reg <= data_i[311];
      data_o_310_sv2v_reg <= data_i[310];
      data_o_309_sv2v_reg <= data_i[309];
      data_o_308_sv2v_reg <= data_i[308];
      data_o_307_sv2v_reg <= data_i[307];
      data_o_306_sv2v_reg <= data_i[306];
      data_o_305_sv2v_reg <= data_i[305];
      data_o_304_sv2v_reg <= data_i[304];
      data_o_303_sv2v_reg <= data_i[303];
      data_o_302_sv2v_reg <= data_i[302];
      data_o_301_sv2v_reg <= data_i[301];
      data_o_300_sv2v_reg <= data_i[300];
      data_o_299_sv2v_reg <= data_i[299];
      data_o_298_sv2v_reg <= data_i[298];
      data_o_297_sv2v_reg <= data_i[297];
      data_o_296_sv2v_reg <= data_i[296];
      data_o_295_sv2v_reg <= data_i[295];
      data_o_294_sv2v_reg <= data_i[294];
      data_o_293_sv2v_reg <= data_i[293];
      data_o_292_sv2v_reg <= data_i[292];
      data_o_291_sv2v_reg <= data_i[291];
      data_o_290_sv2v_reg <= data_i[290];
      data_o_289_sv2v_reg <= data_i[289];
      data_o_288_sv2v_reg <= data_i[288];
      data_o_287_sv2v_reg <= data_i[287];
      data_o_286_sv2v_reg <= data_i[286];
      data_o_285_sv2v_reg <= data_i[285];
      data_o_284_sv2v_reg <= data_i[284];
      data_o_283_sv2v_reg <= data_i[283];
      data_o_282_sv2v_reg <= data_i[282];
      data_o_281_sv2v_reg <= data_i[281];
      data_o_280_sv2v_reg <= data_i[280];
      data_o_279_sv2v_reg <= data_i[279];
      data_o_278_sv2v_reg <= data_i[278];
      data_o_277_sv2v_reg <= data_i[277];
      data_o_276_sv2v_reg <= data_i[276];
      data_o_275_sv2v_reg <= data_i[275];
      data_o_274_sv2v_reg <= data_i[274];
      data_o_273_sv2v_reg <= data_i[273];
      data_o_272_sv2v_reg <= data_i[272];
      data_o_271_sv2v_reg <= data_i[271];
      data_o_270_sv2v_reg <= data_i[270];
      data_o_269_sv2v_reg <= data_i[269];
      data_o_268_sv2v_reg <= data_i[268];
      data_o_267_sv2v_reg <= data_i[267];
      data_o_266_sv2v_reg <= data_i[266];
      data_o_265_sv2v_reg <= data_i[265];
      data_o_264_sv2v_reg <= data_i[264];
      data_o_263_sv2v_reg <= data_i[263];
      data_o_262_sv2v_reg <= data_i[262];
      data_o_261_sv2v_reg <= data_i[261];
      data_o_260_sv2v_reg <= data_i[260];
      data_o_259_sv2v_reg <= data_i[259];
      data_o_258_sv2v_reg <= data_i[258];
      data_o_257_sv2v_reg <= data_i[257];
      data_o_256_sv2v_reg <= data_i[256];
      data_o_255_sv2v_reg <= data_i[255];
      data_o_254_sv2v_reg <= data_i[254];
      data_o_253_sv2v_reg <= data_i[253];
      data_o_252_sv2v_reg <= data_i[252];
      data_o_251_sv2v_reg <= data_i[251];
      data_o_250_sv2v_reg <= data_i[250];
      data_o_249_sv2v_reg <= data_i[249];
      data_o_248_sv2v_reg <= data_i[248];
      data_o_247_sv2v_reg <= data_i[247];
      data_o_246_sv2v_reg <= data_i[246];
      data_o_245_sv2v_reg <= data_i[245];
      data_o_244_sv2v_reg <= data_i[244];
      data_o_243_sv2v_reg <= data_i[243];
      data_o_242_sv2v_reg <= data_i[242];
      data_o_241_sv2v_reg <= data_i[241];
      data_o_240_sv2v_reg <= data_i[240];
      data_o_239_sv2v_reg <= data_i[239];
      data_o_238_sv2v_reg <= data_i[238];
      data_o_237_sv2v_reg <= data_i[237];
      data_o_236_sv2v_reg <= data_i[236];
      data_o_235_sv2v_reg <= data_i[235];
      data_o_234_sv2v_reg <= data_i[234];
      data_o_233_sv2v_reg <= data_i[233];
      data_o_232_sv2v_reg <= data_i[232];
      data_o_231_sv2v_reg <= data_i[231];
      data_o_230_sv2v_reg <= data_i[230];
      data_o_229_sv2v_reg <= data_i[229];
      data_o_228_sv2v_reg <= data_i[228];
      data_o_227_sv2v_reg <= data_i[227];
      data_o_226_sv2v_reg <= data_i[226];
      data_o_225_sv2v_reg <= data_i[225];
      data_o_224_sv2v_reg <= data_i[224];
      data_o_223_sv2v_reg <= data_i[223];
      data_o_222_sv2v_reg <= data_i[222];
      data_o_221_sv2v_reg <= data_i[221];
      data_o_220_sv2v_reg <= data_i[220];
      data_o_219_sv2v_reg <= data_i[219];
      data_o_218_sv2v_reg <= data_i[218];
      data_o_217_sv2v_reg <= data_i[217];
      data_o_216_sv2v_reg <= data_i[216];
      data_o_215_sv2v_reg <= data_i[215];
      data_o_214_sv2v_reg <= data_i[214];
      data_o_213_sv2v_reg <= data_i[213];
      data_o_212_sv2v_reg <= data_i[212];
      data_o_211_sv2v_reg <= data_i[211];
      data_o_210_sv2v_reg <= data_i[210];
      data_o_209_sv2v_reg <= data_i[209];
      data_o_208_sv2v_reg <= data_i[208];
      data_o_207_sv2v_reg <= data_i[207];
      data_o_206_sv2v_reg <= data_i[206];
      data_o_205_sv2v_reg <= data_i[205];
      data_o_204_sv2v_reg <= data_i[204];
      data_o_203_sv2v_reg <= data_i[203];
      data_o_202_sv2v_reg <= data_i[202];
      data_o_201_sv2v_reg <= data_i[201];
      data_o_200_sv2v_reg <= data_i[200];
      data_o_199_sv2v_reg <= data_i[199];
      data_o_198_sv2v_reg <= data_i[198];
      data_o_197_sv2v_reg <= data_i[197];
      data_o_196_sv2v_reg <= data_i[196];
      data_o_195_sv2v_reg <= data_i[195];
      data_o_194_sv2v_reg <= data_i[194];
      data_o_193_sv2v_reg <= data_i[193];
      data_o_192_sv2v_reg <= data_i[192];
      data_o_191_sv2v_reg <= data_i[191];
      data_o_190_sv2v_reg <= data_i[190];
      data_o_189_sv2v_reg <= data_i[189];
      data_o_188_sv2v_reg <= data_i[188];
      data_o_187_sv2v_reg <= data_i[187];
      data_o_186_sv2v_reg <= data_i[186];
      data_o_185_sv2v_reg <= data_i[185];
      data_o_184_sv2v_reg <= data_i[184];
      data_o_183_sv2v_reg <= data_i[183];
      data_o_182_sv2v_reg <= data_i[182];
      data_o_181_sv2v_reg <= data_i[181];
      data_o_180_sv2v_reg <= data_i[180];
      data_o_179_sv2v_reg <= data_i[179];
      data_o_178_sv2v_reg <= data_i[178];
      data_o_177_sv2v_reg <= data_i[177];
      data_o_176_sv2v_reg <= data_i[176];
      data_o_175_sv2v_reg <= data_i[175];
      data_o_174_sv2v_reg <= data_i[174];
      data_o_173_sv2v_reg <= data_i[173];
      data_o_172_sv2v_reg <= data_i[172];
      data_o_171_sv2v_reg <= data_i[171];
      data_o_170_sv2v_reg <= data_i[170];
      data_o_169_sv2v_reg <= data_i[169];
      data_o_168_sv2v_reg <= data_i[168];
      data_o_167_sv2v_reg <= data_i[167];
      data_o_166_sv2v_reg <= data_i[166];
      data_o_165_sv2v_reg <= data_i[165];
      data_o_164_sv2v_reg <= data_i[164];
      data_o_163_sv2v_reg <= data_i[163];
      data_o_162_sv2v_reg <= data_i[162];
      data_o_161_sv2v_reg <= data_i[161];
      data_o_160_sv2v_reg <= data_i[160];
      data_o_159_sv2v_reg <= data_i[159];
      data_o_158_sv2v_reg <= data_i[158];
      data_o_157_sv2v_reg <= data_i[157];
      data_o_156_sv2v_reg <= data_i[156];
      data_o_155_sv2v_reg <= data_i[155];
      data_o_154_sv2v_reg <= data_i[154];
      data_o_153_sv2v_reg <= data_i[153];
      data_o_152_sv2v_reg <= data_i[152];
      data_o_151_sv2v_reg <= data_i[151];
      data_o_150_sv2v_reg <= data_i[150];
      data_o_149_sv2v_reg <= data_i[149];
      data_o_148_sv2v_reg <= data_i[148];
      data_o_147_sv2v_reg <= data_i[147];
      data_o_146_sv2v_reg <= data_i[146];
      data_o_145_sv2v_reg <= data_i[145];
      data_o_144_sv2v_reg <= data_i[144];
      data_o_143_sv2v_reg <= data_i[143];
      data_o_142_sv2v_reg <= data_i[142];
      data_o_141_sv2v_reg <= data_i[141];
      data_o_140_sv2v_reg <= data_i[140];
      data_o_139_sv2v_reg <= data_i[139];
      data_o_138_sv2v_reg <= data_i[138];
      data_o_137_sv2v_reg <= data_i[137];
      data_o_136_sv2v_reg <= data_i[136];
      data_o_135_sv2v_reg <= data_i[135];
      data_o_134_sv2v_reg <= data_i[134];
      data_o_133_sv2v_reg <= data_i[133];
      data_o_132_sv2v_reg <= data_i[132];
      data_o_131_sv2v_reg <= data_i[131];
      data_o_130_sv2v_reg <= data_i[130];
      data_o_129_sv2v_reg <= data_i[129];
      data_o_128_sv2v_reg <= data_i[128];
      data_o_127_sv2v_reg <= data_i[127];
      data_o_126_sv2v_reg <= data_i[126];
      data_o_125_sv2v_reg <= data_i[125];
      data_o_124_sv2v_reg <= data_i[124];
      data_o_123_sv2v_reg <= data_i[123];
      data_o_122_sv2v_reg <= data_i[122];
      data_o_121_sv2v_reg <= data_i[121];
      data_o_120_sv2v_reg <= data_i[120];
      data_o_119_sv2v_reg <= data_i[119];
      data_o_118_sv2v_reg <= data_i[118];
      data_o_117_sv2v_reg <= data_i[117];
      data_o_116_sv2v_reg <= data_i[116];
      data_o_115_sv2v_reg <= data_i[115];
      data_o_114_sv2v_reg <= data_i[114];
      data_o_113_sv2v_reg <= data_i[113];
      data_o_112_sv2v_reg <= data_i[112];
      data_o_111_sv2v_reg <= data_i[111];
      data_o_110_sv2v_reg <= data_i[110];
      data_o_109_sv2v_reg <= data_i[109];
      data_o_108_sv2v_reg <= data_i[108];
      data_o_107_sv2v_reg <= data_i[107];
      data_o_106_sv2v_reg <= data_i[106];
      data_o_105_sv2v_reg <= data_i[105];
      data_o_104_sv2v_reg <= data_i[104];
      data_o_103_sv2v_reg <= data_i[103];
      data_o_102_sv2v_reg <= data_i[102];
      data_o_101_sv2v_reg <= data_i[101];
      data_o_100_sv2v_reg <= data_i[100];
      data_o_99_sv2v_reg <= data_i[99];
      data_o_98_sv2v_reg <= data_i[98];
      data_o_97_sv2v_reg <= data_i[97];
      data_o_96_sv2v_reg <= data_i[96];
      data_o_95_sv2v_reg <= data_i[95];
      data_o_94_sv2v_reg <= data_i[94];
      data_o_93_sv2v_reg <= data_i[93];
      data_o_92_sv2v_reg <= data_i[92];
      data_o_91_sv2v_reg <= data_i[91];
      data_o_90_sv2v_reg <= data_i[90];
      data_o_89_sv2v_reg <= data_i[89];
      data_o_88_sv2v_reg <= data_i[88];
      data_o_87_sv2v_reg <= data_i[87];
      data_o_86_sv2v_reg <= data_i[86];
      data_o_85_sv2v_reg <= data_i[85];
      data_o_84_sv2v_reg <= data_i[84];
      data_o_83_sv2v_reg <= data_i[83];
      data_o_82_sv2v_reg <= data_i[82];
      data_o_81_sv2v_reg <= data_i[81];
      data_o_80_sv2v_reg <= data_i[80];
      data_o_79_sv2v_reg <= data_i[79];
      data_o_78_sv2v_reg <= data_i[78];
      data_o_77_sv2v_reg <= data_i[77];
      data_o_76_sv2v_reg <= data_i[76];
      data_o_75_sv2v_reg <= data_i[75];
      data_o_74_sv2v_reg <= data_i[74];
      data_o_73_sv2v_reg <= data_i[73];
      data_o_72_sv2v_reg <= data_i[72];
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_adder_one_hot_00000008
(
  a_i,
  b_i,
  o
);

  input [7:0] a_i;
  input [7:0] b_i;
  output [7:0] o;
  wire [7:0] o,\rof_0_.aggregate ,\rof_1_.aggregate ,\rof_2_.aggregate ,\rof_3_.aggregate ,
  \rof_4_.aggregate ,\rof_5_.aggregate ,\rof_6_.aggregate ,\rof_7_.aggregate ;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47;
  assign \rof_0_.aggregate [0] = a_i[0] & b_i[0];
  assign \rof_0_.aggregate [1] = a_i[1] & b_i[7];
  assign \rof_0_.aggregate [2] = a_i[2] & b_i[6];
  assign \rof_0_.aggregate [3] = a_i[3] & b_i[5];
  assign \rof_0_.aggregate [4] = a_i[4] & b_i[4];
  assign \rof_0_.aggregate [5] = a_i[5] & b_i[3];
  assign \rof_0_.aggregate [6] = a_i[6] & b_i[2];
  assign \rof_0_.aggregate [7] = a_i[7] & b_i[1];
  assign o[0] = N5 | \rof_0_.aggregate [0];
  assign N5 = N4 | \rof_0_.aggregate [1];
  assign N4 = N3 | \rof_0_.aggregate [2];
  assign N3 = N2 | \rof_0_.aggregate [3];
  assign N2 = N1 | \rof_0_.aggregate [4];
  assign N1 = N0 | \rof_0_.aggregate [5];
  assign N0 = \rof_0_.aggregate [7] | \rof_0_.aggregate [6];
  assign \rof_1_.aggregate [0] = a_i[0] & b_i[1];
  assign \rof_1_.aggregate [1] = a_i[1] & b_i[0];
  assign \rof_1_.aggregate [2] = a_i[2] & b_i[7];
  assign \rof_1_.aggregate [3] = a_i[3] & b_i[6];
  assign \rof_1_.aggregate [4] = a_i[4] & b_i[5];
  assign \rof_1_.aggregate [5] = a_i[5] & b_i[4];
  assign \rof_1_.aggregate [6] = a_i[6] & b_i[3];
  assign \rof_1_.aggregate [7] = a_i[7] & b_i[2];
  assign o[1] = N11 | \rof_1_.aggregate [0];
  assign N11 = N10 | \rof_1_.aggregate [1];
  assign N10 = N9 | \rof_1_.aggregate [2];
  assign N9 = N8 | \rof_1_.aggregate [3];
  assign N8 = N7 | \rof_1_.aggregate [4];
  assign N7 = N6 | \rof_1_.aggregate [5];
  assign N6 = \rof_1_.aggregate [7] | \rof_1_.aggregate [6];
  assign \rof_2_.aggregate [0] = a_i[0] & b_i[2];
  assign \rof_2_.aggregate [1] = a_i[1] & b_i[1];
  assign \rof_2_.aggregate [2] = a_i[2] & b_i[0];
  assign \rof_2_.aggregate [3] = a_i[3] & b_i[7];
  assign \rof_2_.aggregate [4] = a_i[4] & b_i[6];
  assign \rof_2_.aggregate [5] = a_i[5] & b_i[5];
  assign \rof_2_.aggregate [6] = a_i[6] & b_i[4];
  assign \rof_2_.aggregate [7] = a_i[7] & b_i[3];
  assign o[2] = N17 | \rof_2_.aggregate [0];
  assign N17 = N16 | \rof_2_.aggregate [1];
  assign N16 = N15 | \rof_2_.aggregate [2];
  assign N15 = N14 | \rof_2_.aggregate [3];
  assign N14 = N13 | \rof_2_.aggregate [4];
  assign N13 = N12 | \rof_2_.aggregate [5];
  assign N12 = \rof_2_.aggregate [7] | \rof_2_.aggregate [6];
  assign \rof_3_.aggregate [0] = a_i[0] & b_i[3];
  assign \rof_3_.aggregate [1] = a_i[1] & b_i[2];
  assign \rof_3_.aggregate [2] = a_i[2] & b_i[1];
  assign \rof_3_.aggregate [3] = a_i[3] & b_i[0];
  assign \rof_3_.aggregate [4] = a_i[4] & b_i[7];
  assign \rof_3_.aggregate [5] = a_i[5] & b_i[6];
  assign \rof_3_.aggregate [6] = a_i[6] & b_i[5];
  assign \rof_3_.aggregate [7] = a_i[7] & b_i[4];
  assign o[3] = N23 | \rof_3_.aggregate [0];
  assign N23 = N22 | \rof_3_.aggregate [1];
  assign N22 = N21 | \rof_3_.aggregate [2];
  assign N21 = N20 | \rof_3_.aggregate [3];
  assign N20 = N19 | \rof_3_.aggregate [4];
  assign N19 = N18 | \rof_3_.aggregate [5];
  assign N18 = \rof_3_.aggregate [7] | \rof_3_.aggregate [6];
  assign \rof_4_.aggregate [0] = a_i[0] & b_i[4];
  assign \rof_4_.aggregate [1] = a_i[1] & b_i[3];
  assign \rof_4_.aggregate [2] = a_i[2] & b_i[2];
  assign \rof_4_.aggregate [3] = a_i[3] & b_i[1];
  assign \rof_4_.aggregate [4] = a_i[4] & b_i[0];
  assign \rof_4_.aggregate [5] = a_i[5] & b_i[7];
  assign \rof_4_.aggregate [6] = a_i[6] & b_i[6];
  assign \rof_4_.aggregate [7] = a_i[7] & b_i[5];
  assign o[4] = N29 | \rof_4_.aggregate [0];
  assign N29 = N28 | \rof_4_.aggregate [1];
  assign N28 = N27 | \rof_4_.aggregate [2];
  assign N27 = N26 | \rof_4_.aggregate [3];
  assign N26 = N25 | \rof_4_.aggregate [4];
  assign N25 = N24 | \rof_4_.aggregate [5];
  assign N24 = \rof_4_.aggregate [7] | \rof_4_.aggregate [6];
  assign \rof_5_.aggregate [0] = a_i[0] & b_i[5];
  assign \rof_5_.aggregate [1] = a_i[1] & b_i[4];
  assign \rof_5_.aggregate [2] = a_i[2] & b_i[3];
  assign \rof_5_.aggregate [3] = a_i[3] & b_i[2];
  assign \rof_5_.aggregate [4] = a_i[4] & b_i[1];
  assign \rof_5_.aggregate [5] = a_i[5] & b_i[0];
  assign \rof_5_.aggregate [6] = a_i[6] & b_i[7];
  assign \rof_5_.aggregate [7] = a_i[7] & b_i[6];
  assign o[5] = N35 | \rof_5_.aggregate [0];
  assign N35 = N34 | \rof_5_.aggregate [1];
  assign N34 = N33 | \rof_5_.aggregate [2];
  assign N33 = N32 | \rof_5_.aggregate [3];
  assign N32 = N31 | \rof_5_.aggregate [4];
  assign N31 = N30 | \rof_5_.aggregate [5];
  assign N30 = \rof_5_.aggregate [7] | \rof_5_.aggregate [6];
  assign \rof_6_.aggregate [0] = a_i[0] & b_i[6];
  assign \rof_6_.aggregate [1] = a_i[1] & b_i[5];
  assign \rof_6_.aggregate [2] = a_i[2] & b_i[4];
  assign \rof_6_.aggregate [3] = a_i[3] & b_i[3];
  assign \rof_6_.aggregate [4] = a_i[4] & b_i[2];
  assign \rof_6_.aggregate [5] = a_i[5] & b_i[1];
  assign \rof_6_.aggregate [6] = a_i[6] & b_i[0];
  assign \rof_6_.aggregate [7] = a_i[7] & b_i[7];
  assign o[6] = N41 | \rof_6_.aggregate [0];
  assign N41 = N40 | \rof_6_.aggregate [1];
  assign N40 = N39 | \rof_6_.aggregate [2];
  assign N39 = N38 | \rof_6_.aggregate [3];
  assign N38 = N37 | \rof_6_.aggregate [4];
  assign N37 = N36 | \rof_6_.aggregate [5];
  assign N36 = \rof_6_.aggregate [7] | \rof_6_.aggregate [6];
  assign \rof_7_.aggregate [0] = a_i[0] & b_i[7];
  assign \rof_7_.aggregate [1] = a_i[1] & b_i[6];
  assign \rof_7_.aggregate [2] = a_i[2] & b_i[5];
  assign \rof_7_.aggregate [3] = a_i[3] & b_i[4];
  assign \rof_7_.aggregate [4] = a_i[4] & b_i[3];
  assign \rof_7_.aggregate [5] = a_i[5] & b_i[2];
  assign \rof_7_.aggregate [6] = a_i[6] & b_i[1];
  assign \rof_7_.aggregate [7] = a_i[7] & b_i[0];
  assign o[7] = N47 | \rof_7_.aggregate [0];
  assign N47 = N46 | \rof_7_.aggregate [1];
  assign N46 = N45 | \rof_7_.aggregate [2];
  assign N45 = N44 | \rof_7_.aggregate [3];
  assign N44 = N43 | \rof_7_.aggregate [4];
  assign N43 = N42 | \rof_7_.aggregate [5];
  assign N42 = \rof_7_.aggregate [7] | \rof_7_.aggregate [6];

endmodule



module bsg_mux_one_hot_00000040_00000008
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [511:0] data_i;
  input [7:0] sel_one_hot_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383;
  wire [511:0] data_masked;
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[1];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[1];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[1];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[2];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[2];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[2];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[2];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[2];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[2];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[2];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[2];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[2];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[2];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[2];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[2];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[2];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[2];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[2];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[2];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[2];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[2];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[2];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[2];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[2];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[2];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[2];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[2];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[2];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[2];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[2];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[2];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[2];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[2];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[2];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[2];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[2];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[2];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[2];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[2];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[2];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[2];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[2];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[2];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[2];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[2];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[2];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[2];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[2];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[2];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[2];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[2];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[2];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[2];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[2];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[2];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[2];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[2];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[2];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[2];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[2];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[2];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[2];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[2];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[2];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[2];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[2];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[2];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[3];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[3];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[3];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[3];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[3];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[3];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[3];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[3];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[3];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[3];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[3];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[3];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[3];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[3];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[3];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[3];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[3];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[3];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[3];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[3];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[3];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[3];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[3];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[3];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[3];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[3];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[3];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[3];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[3];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[3];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[3];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[3];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[3];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[3];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[3];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[3];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[3];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[3];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[3];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[3];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[3];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[3];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[3];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[3];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[3];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[3];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[3];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[3];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[3];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[3];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[3];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[3];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[3];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[3];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[3];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[3];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[3];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[3];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[3];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[3];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[3];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[3];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[3];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[3];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[4];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[4];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[4];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[4];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[4];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[4];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[4];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[4];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[4];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[4];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[4];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[4];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[4];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[4];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[4];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[4];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[4];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[4];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[4];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[4];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[4];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[4];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[4];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[4];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[4];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[4];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[4];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[4];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[4];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[4];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[4];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[4];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[4];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[4];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[4];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[4];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[4];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[4];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[4];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[4];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[4];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[4];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[4];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[4];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[4];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[4];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[4];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[4];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[4];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[4];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[4];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[4];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[4];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[4];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[4];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[4];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[4];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[4];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[4];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[4];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[4];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[4];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[4];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[4];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[5];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[5];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[5];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[5];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[5];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[5];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[5];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[5];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[5];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[5];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[5];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[5];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[5];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[5];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[5];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[5];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[5];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[5];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[5];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[5];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[5];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[5];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[5];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[5];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[5];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[5];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[5];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[5];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[5];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[5];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[5];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[5];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[5];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[5];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[5];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[5];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[5];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[5];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[5];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[5];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[5];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[5];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[5];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[5];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[5];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[5];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[5];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[5];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[5];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[5];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[5];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[5];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[5];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[5];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[5];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[5];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[5];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[5];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[5];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[5];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[5];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[5];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[5];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[5];
  assign data_masked[447] = data_i[447] & sel_one_hot_i[6];
  assign data_masked[446] = data_i[446] & sel_one_hot_i[6];
  assign data_masked[445] = data_i[445] & sel_one_hot_i[6];
  assign data_masked[444] = data_i[444] & sel_one_hot_i[6];
  assign data_masked[443] = data_i[443] & sel_one_hot_i[6];
  assign data_masked[442] = data_i[442] & sel_one_hot_i[6];
  assign data_masked[441] = data_i[441] & sel_one_hot_i[6];
  assign data_masked[440] = data_i[440] & sel_one_hot_i[6];
  assign data_masked[439] = data_i[439] & sel_one_hot_i[6];
  assign data_masked[438] = data_i[438] & sel_one_hot_i[6];
  assign data_masked[437] = data_i[437] & sel_one_hot_i[6];
  assign data_masked[436] = data_i[436] & sel_one_hot_i[6];
  assign data_masked[435] = data_i[435] & sel_one_hot_i[6];
  assign data_masked[434] = data_i[434] & sel_one_hot_i[6];
  assign data_masked[433] = data_i[433] & sel_one_hot_i[6];
  assign data_masked[432] = data_i[432] & sel_one_hot_i[6];
  assign data_masked[431] = data_i[431] & sel_one_hot_i[6];
  assign data_masked[430] = data_i[430] & sel_one_hot_i[6];
  assign data_masked[429] = data_i[429] & sel_one_hot_i[6];
  assign data_masked[428] = data_i[428] & sel_one_hot_i[6];
  assign data_masked[427] = data_i[427] & sel_one_hot_i[6];
  assign data_masked[426] = data_i[426] & sel_one_hot_i[6];
  assign data_masked[425] = data_i[425] & sel_one_hot_i[6];
  assign data_masked[424] = data_i[424] & sel_one_hot_i[6];
  assign data_masked[423] = data_i[423] & sel_one_hot_i[6];
  assign data_masked[422] = data_i[422] & sel_one_hot_i[6];
  assign data_masked[421] = data_i[421] & sel_one_hot_i[6];
  assign data_masked[420] = data_i[420] & sel_one_hot_i[6];
  assign data_masked[419] = data_i[419] & sel_one_hot_i[6];
  assign data_masked[418] = data_i[418] & sel_one_hot_i[6];
  assign data_masked[417] = data_i[417] & sel_one_hot_i[6];
  assign data_masked[416] = data_i[416] & sel_one_hot_i[6];
  assign data_masked[415] = data_i[415] & sel_one_hot_i[6];
  assign data_masked[414] = data_i[414] & sel_one_hot_i[6];
  assign data_masked[413] = data_i[413] & sel_one_hot_i[6];
  assign data_masked[412] = data_i[412] & sel_one_hot_i[6];
  assign data_masked[411] = data_i[411] & sel_one_hot_i[6];
  assign data_masked[410] = data_i[410] & sel_one_hot_i[6];
  assign data_masked[409] = data_i[409] & sel_one_hot_i[6];
  assign data_masked[408] = data_i[408] & sel_one_hot_i[6];
  assign data_masked[407] = data_i[407] & sel_one_hot_i[6];
  assign data_masked[406] = data_i[406] & sel_one_hot_i[6];
  assign data_masked[405] = data_i[405] & sel_one_hot_i[6];
  assign data_masked[404] = data_i[404] & sel_one_hot_i[6];
  assign data_masked[403] = data_i[403] & sel_one_hot_i[6];
  assign data_masked[402] = data_i[402] & sel_one_hot_i[6];
  assign data_masked[401] = data_i[401] & sel_one_hot_i[6];
  assign data_masked[400] = data_i[400] & sel_one_hot_i[6];
  assign data_masked[399] = data_i[399] & sel_one_hot_i[6];
  assign data_masked[398] = data_i[398] & sel_one_hot_i[6];
  assign data_masked[397] = data_i[397] & sel_one_hot_i[6];
  assign data_masked[396] = data_i[396] & sel_one_hot_i[6];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[6];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[6];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[6];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[6];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[6];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[6];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[6];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[6];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[6];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[6];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[6];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[6];
  assign data_masked[511] = data_i[511] & sel_one_hot_i[7];
  assign data_masked[510] = data_i[510] & sel_one_hot_i[7];
  assign data_masked[509] = data_i[509] & sel_one_hot_i[7];
  assign data_masked[508] = data_i[508] & sel_one_hot_i[7];
  assign data_masked[507] = data_i[507] & sel_one_hot_i[7];
  assign data_masked[506] = data_i[506] & sel_one_hot_i[7];
  assign data_masked[505] = data_i[505] & sel_one_hot_i[7];
  assign data_masked[504] = data_i[504] & sel_one_hot_i[7];
  assign data_masked[503] = data_i[503] & sel_one_hot_i[7];
  assign data_masked[502] = data_i[502] & sel_one_hot_i[7];
  assign data_masked[501] = data_i[501] & sel_one_hot_i[7];
  assign data_masked[500] = data_i[500] & sel_one_hot_i[7];
  assign data_masked[499] = data_i[499] & sel_one_hot_i[7];
  assign data_masked[498] = data_i[498] & sel_one_hot_i[7];
  assign data_masked[497] = data_i[497] & sel_one_hot_i[7];
  assign data_masked[496] = data_i[496] & sel_one_hot_i[7];
  assign data_masked[495] = data_i[495] & sel_one_hot_i[7];
  assign data_masked[494] = data_i[494] & sel_one_hot_i[7];
  assign data_masked[493] = data_i[493] & sel_one_hot_i[7];
  assign data_masked[492] = data_i[492] & sel_one_hot_i[7];
  assign data_masked[491] = data_i[491] & sel_one_hot_i[7];
  assign data_masked[490] = data_i[490] & sel_one_hot_i[7];
  assign data_masked[489] = data_i[489] & sel_one_hot_i[7];
  assign data_masked[488] = data_i[488] & sel_one_hot_i[7];
  assign data_masked[487] = data_i[487] & sel_one_hot_i[7];
  assign data_masked[486] = data_i[486] & sel_one_hot_i[7];
  assign data_masked[485] = data_i[485] & sel_one_hot_i[7];
  assign data_masked[484] = data_i[484] & sel_one_hot_i[7];
  assign data_masked[483] = data_i[483] & sel_one_hot_i[7];
  assign data_masked[482] = data_i[482] & sel_one_hot_i[7];
  assign data_masked[481] = data_i[481] & sel_one_hot_i[7];
  assign data_masked[480] = data_i[480] & sel_one_hot_i[7];
  assign data_masked[479] = data_i[479] & sel_one_hot_i[7];
  assign data_masked[478] = data_i[478] & sel_one_hot_i[7];
  assign data_masked[477] = data_i[477] & sel_one_hot_i[7];
  assign data_masked[476] = data_i[476] & sel_one_hot_i[7];
  assign data_masked[475] = data_i[475] & sel_one_hot_i[7];
  assign data_masked[474] = data_i[474] & sel_one_hot_i[7];
  assign data_masked[473] = data_i[473] & sel_one_hot_i[7];
  assign data_masked[472] = data_i[472] & sel_one_hot_i[7];
  assign data_masked[471] = data_i[471] & sel_one_hot_i[7];
  assign data_masked[470] = data_i[470] & sel_one_hot_i[7];
  assign data_masked[469] = data_i[469] & sel_one_hot_i[7];
  assign data_masked[468] = data_i[468] & sel_one_hot_i[7];
  assign data_masked[467] = data_i[467] & sel_one_hot_i[7];
  assign data_masked[466] = data_i[466] & sel_one_hot_i[7];
  assign data_masked[465] = data_i[465] & sel_one_hot_i[7];
  assign data_masked[464] = data_i[464] & sel_one_hot_i[7];
  assign data_masked[463] = data_i[463] & sel_one_hot_i[7];
  assign data_masked[462] = data_i[462] & sel_one_hot_i[7];
  assign data_masked[461] = data_i[461] & sel_one_hot_i[7];
  assign data_masked[460] = data_i[460] & sel_one_hot_i[7];
  assign data_masked[459] = data_i[459] & sel_one_hot_i[7];
  assign data_masked[458] = data_i[458] & sel_one_hot_i[7];
  assign data_masked[457] = data_i[457] & sel_one_hot_i[7];
  assign data_masked[456] = data_i[456] & sel_one_hot_i[7];
  assign data_masked[455] = data_i[455] & sel_one_hot_i[7];
  assign data_masked[454] = data_i[454] & sel_one_hot_i[7];
  assign data_masked[453] = data_i[453] & sel_one_hot_i[7];
  assign data_masked[452] = data_i[452] & sel_one_hot_i[7];
  assign data_masked[451] = data_i[451] & sel_one_hot_i[7];
  assign data_masked[450] = data_i[450] & sel_one_hot_i[7];
  assign data_masked[449] = data_i[449] & sel_one_hot_i[7];
  assign data_masked[448] = data_i[448] & sel_one_hot_i[7];
  assign data_o[0] = N5 | data_masked[0];
  assign N5 = N4 | data_masked[64];
  assign N4 = N3 | data_masked[128];
  assign N3 = N2 | data_masked[192];
  assign N2 = N1 | data_masked[256];
  assign N1 = N0 | data_masked[320];
  assign N0 = data_masked[448] | data_masked[384];
  assign data_o[1] = N11 | data_masked[1];
  assign N11 = N10 | data_masked[65];
  assign N10 = N9 | data_masked[129];
  assign N9 = N8 | data_masked[193];
  assign N8 = N7 | data_masked[257];
  assign N7 = N6 | data_masked[321];
  assign N6 = data_masked[449] | data_masked[385];
  assign data_o[2] = N17 | data_masked[2];
  assign N17 = N16 | data_masked[66];
  assign N16 = N15 | data_masked[130];
  assign N15 = N14 | data_masked[194];
  assign N14 = N13 | data_masked[258];
  assign N13 = N12 | data_masked[322];
  assign N12 = data_masked[450] | data_masked[386];
  assign data_o[3] = N23 | data_masked[3];
  assign N23 = N22 | data_masked[67];
  assign N22 = N21 | data_masked[131];
  assign N21 = N20 | data_masked[195];
  assign N20 = N19 | data_masked[259];
  assign N19 = N18 | data_masked[323];
  assign N18 = data_masked[451] | data_masked[387];
  assign data_o[4] = N29 | data_masked[4];
  assign N29 = N28 | data_masked[68];
  assign N28 = N27 | data_masked[132];
  assign N27 = N26 | data_masked[196];
  assign N26 = N25 | data_masked[260];
  assign N25 = N24 | data_masked[324];
  assign N24 = data_masked[452] | data_masked[388];
  assign data_o[5] = N35 | data_masked[5];
  assign N35 = N34 | data_masked[69];
  assign N34 = N33 | data_masked[133];
  assign N33 = N32 | data_masked[197];
  assign N32 = N31 | data_masked[261];
  assign N31 = N30 | data_masked[325];
  assign N30 = data_masked[453] | data_masked[389];
  assign data_o[6] = N41 | data_masked[6];
  assign N41 = N40 | data_masked[70];
  assign N40 = N39 | data_masked[134];
  assign N39 = N38 | data_masked[198];
  assign N38 = N37 | data_masked[262];
  assign N37 = N36 | data_masked[326];
  assign N36 = data_masked[454] | data_masked[390];
  assign data_o[7] = N47 | data_masked[7];
  assign N47 = N46 | data_masked[71];
  assign N46 = N45 | data_masked[135];
  assign N45 = N44 | data_masked[199];
  assign N44 = N43 | data_masked[263];
  assign N43 = N42 | data_masked[327];
  assign N42 = data_masked[455] | data_masked[391];
  assign data_o[8] = N53 | data_masked[8];
  assign N53 = N52 | data_masked[72];
  assign N52 = N51 | data_masked[136];
  assign N51 = N50 | data_masked[200];
  assign N50 = N49 | data_masked[264];
  assign N49 = N48 | data_masked[328];
  assign N48 = data_masked[456] | data_masked[392];
  assign data_o[9] = N59 | data_masked[9];
  assign N59 = N58 | data_masked[73];
  assign N58 = N57 | data_masked[137];
  assign N57 = N56 | data_masked[201];
  assign N56 = N55 | data_masked[265];
  assign N55 = N54 | data_masked[329];
  assign N54 = data_masked[457] | data_masked[393];
  assign data_o[10] = N65 | data_masked[10];
  assign N65 = N64 | data_masked[74];
  assign N64 = N63 | data_masked[138];
  assign N63 = N62 | data_masked[202];
  assign N62 = N61 | data_masked[266];
  assign N61 = N60 | data_masked[330];
  assign N60 = data_masked[458] | data_masked[394];
  assign data_o[11] = N71 | data_masked[11];
  assign N71 = N70 | data_masked[75];
  assign N70 = N69 | data_masked[139];
  assign N69 = N68 | data_masked[203];
  assign N68 = N67 | data_masked[267];
  assign N67 = N66 | data_masked[331];
  assign N66 = data_masked[459] | data_masked[395];
  assign data_o[12] = N77 | data_masked[12];
  assign N77 = N76 | data_masked[76];
  assign N76 = N75 | data_masked[140];
  assign N75 = N74 | data_masked[204];
  assign N74 = N73 | data_masked[268];
  assign N73 = N72 | data_masked[332];
  assign N72 = data_masked[460] | data_masked[396];
  assign data_o[13] = N83 | data_masked[13];
  assign N83 = N82 | data_masked[77];
  assign N82 = N81 | data_masked[141];
  assign N81 = N80 | data_masked[205];
  assign N80 = N79 | data_masked[269];
  assign N79 = N78 | data_masked[333];
  assign N78 = data_masked[461] | data_masked[397];
  assign data_o[14] = N89 | data_masked[14];
  assign N89 = N88 | data_masked[78];
  assign N88 = N87 | data_masked[142];
  assign N87 = N86 | data_masked[206];
  assign N86 = N85 | data_masked[270];
  assign N85 = N84 | data_masked[334];
  assign N84 = data_masked[462] | data_masked[398];
  assign data_o[15] = N95 | data_masked[15];
  assign N95 = N94 | data_masked[79];
  assign N94 = N93 | data_masked[143];
  assign N93 = N92 | data_masked[207];
  assign N92 = N91 | data_masked[271];
  assign N91 = N90 | data_masked[335];
  assign N90 = data_masked[463] | data_masked[399];
  assign data_o[16] = N101 | data_masked[16];
  assign N101 = N100 | data_masked[80];
  assign N100 = N99 | data_masked[144];
  assign N99 = N98 | data_masked[208];
  assign N98 = N97 | data_masked[272];
  assign N97 = N96 | data_masked[336];
  assign N96 = data_masked[464] | data_masked[400];
  assign data_o[17] = N107 | data_masked[17];
  assign N107 = N106 | data_masked[81];
  assign N106 = N105 | data_masked[145];
  assign N105 = N104 | data_masked[209];
  assign N104 = N103 | data_masked[273];
  assign N103 = N102 | data_masked[337];
  assign N102 = data_masked[465] | data_masked[401];
  assign data_o[18] = N113 | data_masked[18];
  assign N113 = N112 | data_masked[82];
  assign N112 = N111 | data_masked[146];
  assign N111 = N110 | data_masked[210];
  assign N110 = N109 | data_masked[274];
  assign N109 = N108 | data_masked[338];
  assign N108 = data_masked[466] | data_masked[402];
  assign data_o[19] = N119 | data_masked[19];
  assign N119 = N118 | data_masked[83];
  assign N118 = N117 | data_masked[147];
  assign N117 = N116 | data_masked[211];
  assign N116 = N115 | data_masked[275];
  assign N115 = N114 | data_masked[339];
  assign N114 = data_masked[467] | data_masked[403];
  assign data_o[20] = N125 | data_masked[20];
  assign N125 = N124 | data_masked[84];
  assign N124 = N123 | data_masked[148];
  assign N123 = N122 | data_masked[212];
  assign N122 = N121 | data_masked[276];
  assign N121 = N120 | data_masked[340];
  assign N120 = data_masked[468] | data_masked[404];
  assign data_o[21] = N131 | data_masked[21];
  assign N131 = N130 | data_masked[85];
  assign N130 = N129 | data_masked[149];
  assign N129 = N128 | data_masked[213];
  assign N128 = N127 | data_masked[277];
  assign N127 = N126 | data_masked[341];
  assign N126 = data_masked[469] | data_masked[405];
  assign data_o[22] = N137 | data_masked[22];
  assign N137 = N136 | data_masked[86];
  assign N136 = N135 | data_masked[150];
  assign N135 = N134 | data_masked[214];
  assign N134 = N133 | data_masked[278];
  assign N133 = N132 | data_masked[342];
  assign N132 = data_masked[470] | data_masked[406];
  assign data_o[23] = N143 | data_masked[23];
  assign N143 = N142 | data_masked[87];
  assign N142 = N141 | data_masked[151];
  assign N141 = N140 | data_masked[215];
  assign N140 = N139 | data_masked[279];
  assign N139 = N138 | data_masked[343];
  assign N138 = data_masked[471] | data_masked[407];
  assign data_o[24] = N149 | data_masked[24];
  assign N149 = N148 | data_masked[88];
  assign N148 = N147 | data_masked[152];
  assign N147 = N146 | data_masked[216];
  assign N146 = N145 | data_masked[280];
  assign N145 = N144 | data_masked[344];
  assign N144 = data_masked[472] | data_masked[408];
  assign data_o[25] = N155 | data_masked[25];
  assign N155 = N154 | data_masked[89];
  assign N154 = N153 | data_masked[153];
  assign N153 = N152 | data_masked[217];
  assign N152 = N151 | data_masked[281];
  assign N151 = N150 | data_masked[345];
  assign N150 = data_masked[473] | data_masked[409];
  assign data_o[26] = N161 | data_masked[26];
  assign N161 = N160 | data_masked[90];
  assign N160 = N159 | data_masked[154];
  assign N159 = N158 | data_masked[218];
  assign N158 = N157 | data_masked[282];
  assign N157 = N156 | data_masked[346];
  assign N156 = data_masked[474] | data_masked[410];
  assign data_o[27] = N167 | data_masked[27];
  assign N167 = N166 | data_masked[91];
  assign N166 = N165 | data_masked[155];
  assign N165 = N164 | data_masked[219];
  assign N164 = N163 | data_masked[283];
  assign N163 = N162 | data_masked[347];
  assign N162 = data_masked[475] | data_masked[411];
  assign data_o[28] = N173 | data_masked[28];
  assign N173 = N172 | data_masked[92];
  assign N172 = N171 | data_masked[156];
  assign N171 = N170 | data_masked[220];
  assign N170 = N169 | data_masked[284];
  assign N169 = N168 | data_masked[348];
  assign N168 = data_masked[476] | data_masked[412];
  assign data_o[29] = N179 | data_masked[29];
  assign N179 = N178 | data_masked[93];
  assign N178 = N177 | data_masked[157];
  assign N177 = N176 | data_masked[221];
  assign N176 = N175 | data_masked[285];
  assign N175 = N174 | data_masked[349];
  assign N174 = data_masked[477] | data_masked[413];
  assign data_o[30] = N185 | data_masked[30];
  assign N185 = N184 | data_masked[94];
  assign N184 = N183 | data_masked[158];
  assign N183 = N182 | data_masked[222];
  assign N182 = N181 | data_masked[286];
  assign N181 = N180 | data_masked[350];
  assign N180 = data_masked[478] | data_masked[414];
  assign data_o[31] = N191 | data_masked[31];
  assign N191 = N190 | data_masked[95];
  assign N190 = N189 | data_masked[159];
  assign N189 = N188 | data_masked[223];
  assign N188 = N187 | data_masked[287];
  assign N187 = N186 | data_masked[351];
  assign N186 = data_masked[479] | data_masked[415];
  assign data_o[32] = N197 | data_masked[32];
  assign N197 = N196 | data_masked[96];
  assign N196 = N195 | data_masked[160];
  assign N195 = N194 | data_masked[224];
  assign N194 = N193 | data_masked[288];
  assign N193 = N192 | data_masked[352];
  assign N192 = data_masked[480] | data_masked[416];
  assign data_o[33] = N203 | data_masked[33];
  assign N203 = N202 | data_masked[97];
  assign N202 = N201 | data_masked[161];
  assign N201 = N200 | data_masked[225];
  assign N200 = N199 | data_masked[289];
  assign N199 = N198 | data_masked[353];
  assign N198 = data_masked[481] | data_masked[417];
  assign data_o[34] = N209 | data_masked[34];
  assign N209 = N208 | data_masked[98];
  assign N208 = N207 | data_masked[162];
  assign N207 = N206 | data_masked[226];
  assign N206 = N205 | data_masked[290];
  assign N205 = N204 | data_masked[354];
  assign N204 = data_masked[482] | data_masked[418];
  assign data_o[35] = N215 | data_masked[35];
  assign N215 = N214 | data_masked[99];
  assign N214 = N213 | data_masked[163];
  assign N213 = N212 | data_masked[227];
  assign N212 = N211 | data_masked[291];
  assign N211 = N210 | data_masked[355];
  assign N210 = data_masked[483] | data_masked[419];
  assign data_o[36] = N221 | data_masked[36];
  assign N221 = N220 | data_masked[100];
  assign N220 = N219 | data_masked[164];
  assign N219 = N218 | data_masked[228];
  assign N218 = N217 | data_masked[292];
  assign N217 = N216 | data_masked[356];
  assign N216 = data_masked[484] | data_masked[420];
  assign data_o[37] = N227 | data_masked[37];
  assign N227 = N226 | data_masked[101];
  assign N226 = N225 | data_masked[165];
  assign N225 = N224 | data_masked[229];
  assign N224 = N223 | data_masked[293];
  assign N223 = N222 | data_masked[357];
  assign N222 = data_masked[485] | data_masked[421];
  assign data_o[38] = N233 | data_masked[38];
  assign N233 = N232 | data_masked[102];
  assign N232 = N231 | data_masked[166];
  assign N231 = N230 | data_masked[230];
  assign N230 = N229 | data_masked[294];
  assign N229 = N228 | data_masked[358];
  assign N228 = data_masked[486] | data_masked[422];
  assign data_o[39] = N239 | data_masked[39];
  assign N239 = N238 | data_masked[103];
  assign N238 = N237 | data_masked[167];
  assign N237 = N236 | data_masked[231];
  assign N236 = N235 | data_masked[295];
  assign N235 = N234 | data_masked[359];
  assign N234 = data_masked[487] | data_masked[423];
  assign data_o[40] = N245 | data_masked[40];
  assign N245 = N244 | data_masked[104];
  assign N244 = N243 | data_masked[168];
  assign N243 = N242 | data_masked[232];
  assign N242 = N241 | data_masked[296];
  assign N241 = N240 | data_masked[360];
  assign N240 = data_masked[488] | data_masked[424];
  assign data_o[41] = N251 | data_masked[41];
  assign N251 = N250 | data_masked[105];
  assign N250 = N249 | data_masked[169];
  assign N249 = N248 | data_masked[233];
  assign N248 = N247 | data_masked[297];
  assign N247 = N246 | data_masked[361];
  assign N246 = data_masked[489] | data_masked[425];
  assign data_o[42] = N257 | data_masked[42];
  assign N257 = N256 | data_masked[106];
  assign N256 = N255 | data_masked[170];
  assign N255 = N254 | data_masked[234];
  assign N254 = N253 | data_masked[298];
  assign N253 = N252 | data_masked[362];
  assign N252 = data_masked[490] | data_masked[426];
  assign data_o[43] = N263 | data_masked[43];
  assign N263 = N262 | data_masked[107];
  assign N262 = N261 | data_masked[171];
  assign N261 = N260 | data_masked[235];
  assign N260 = N259 | data_masked[299];
  assign N259 = N258 | data_masked[363];
  assign N258 = data_masked[491] | data_masked[427];
  assign data_o[44] = N269 | data_masked[44];
  assign N269 = N268 | data_masked[108];
  assign N268 = N267 | data_masked[172];
  assign N267 = N266 | data_masked[236];
  assign N266 = N265 | data_masked[300];
  assign N265 = N264 | data_masked[364];
  assign N264 = data_masked[492] | data_masked[428];
  assign data_o[45] = N275 | data_masked[45];
  assign N275 = N274 | data_masked[109];
  assign N274 = N273 | data_masked[173];
  assign N273 = N272 | data_masked[237];
  assign N272 = N271 | data_masked[301];
  assign N271 = N270 | data_masked[365];
  assign N270 = data_masked[493] | data_masked[429];
  assign data_o[46] = N281 | data_masked[46];
  assign N281 = N280 | data_masked[110];
  assign N280 = N279 | data_masked[174];
  assign N279 = N278 | data_masked[238];
  assign N278 = N277 | data_masked[302];
  assign N277 = N276 | data_masked[366];
  assign N276 = data_masked[494] | data_masked[430];
  assign data_o[47] = N287 | data_masked[47];
  assign N287 = N286 | data_masked[111];
  assign N286 = N285 | data_masked[175];
  assign N285 = N284 | data_masked[239];
  assign N284 = N283 | data_masked[303];
  assign N283 = N282 | data_masked[367];
  assign N282 = data_masked[495] | data_masked[431];
  assign data_o[48] = N293 | data_masked[48];
  assign N293 = N292 | data_masked[112];
  assign N292 = N291 | data_masked[176];
  assign N291 = N290 | data_masked[240];
  assign N290 = N289 | data_masked[304];
  assign N289 = N288 | data_masked[368];
  assign N288 = data_masked[496] | data_masked[432];
  assign data_o[49] = N299 | data_masked[49];
  assign N299 = N298 | data_masked[113];
  assign N298 = N297 | data_masked[177];
  assign N297 = N296 | data_masked[241];
  assign N296 = N295 | data_masked[305];
  assign N295 = N294 | data_masked[369];
  assign N294 = data_masked[497] | data_masked[433];
  assign data_o[50] = N305 | data_masked[50];
  assign N305 = N304 | data_masked[114];
  assign N304 = N303 | data_masked[178];
  assign N303 = N302 | data_masked[242];
  assign N302 = N301 | data_masked[306];
  assign N301 = N300 | data_masked[370];
  assign N300 = data_masked[498] | data_masked[434];
  assign data_o[51] = N311 | data_masked[51];
  assign N311 = N310 | data_masked[115];
  assign N310 = N309 | data_masked[179];
  assign N309 = N308 | data_masked[243];
  assign N308 = N307 | data_masked[307];
  assign N307 = N306 | data_masked[371];
  assign N306 = data_masked[499] | data_masked[435];
  assign data_o[52] = N317 | data_masked[52];
  assign N317 = N316 | data_masked[116];
  assign N316 = N315 | data_masked[180];
  assign N315 = N314 | data_masked[244];
  assign N314 = N313 | data_masked[308];
  assign N313 = N312 | data_masked[372];
  assign N312 = data_masked[500] | data_masked[436];
  assign data_o[53] = N323 | data_masked[53];
  assign N323 = N322 | data_masked[117];
  assign N322 = N321 | data_masked[181];
  assign N321 = N320 | data_masked[245];
  assign N320 = N319 | data_masked[309];
  assign N319 = N318 | data_masked[373];
  assign N318 = data_masked[501] | data_masked[437];
  assign data_o[54] = N329 | data_masked[54];
  assign N329 = N328 | data_masked[118];
  assign N328 = N327 | data_masked[182];
  assign N327 = N326 | data_masked[246];
  assign N326 = N325 | data_masked[310];
  assign N325 = N324 | data_masked[374];
  assign N324 = data_masked[502] | data_masked[438];
  assign data_o[55] = N335 | data_masked[55];
  assign N335 = N334 | data_masked[119];
  assign N334 = N333 | data_masked[183];
  assign N333 = N332 | data_masked[247];
  assign N332 = N331 | data_masked[311];
  assign N331 = N330 | data_masked[375];
  assign N330 = data_masked[503] | data_masked[439];
  assign data_o[56] = N341 | data_masked[56];
  assign N341 = N340 | data_masked[120];
  assign N340 = N339 | data_masked[184];
  assign N339 = N338 | data_masked[248];
  assign N338 = N337 | data_masked[312];
  assign N337 = N336 | data_masked[376];
  assign N336 = data_masked[504] | data_masked[440];
  assign data_o[57] = N347 | data_masked[57];
  assign N347 = N346 | data_masked[121];
  assign N346 = N345 | data_masked[185];
  assign N345 = N344 | data_masked[249];
  assign N344 = N343 | data_masked[313];
  assign N343 = N342 | data_masked[377];
  assign N342 = data_masked[505] | data_masked[441];
  assign data_o[58] = N353 | data_masked[58];
  assign N353 = N352 | data_masked[122];
  assign N352 = N351 | data_masked[186];
  assign N351 = N350 | data_masked[250];
  assign N350 = N349 | data_masked[314];
  assign N349 = N348 | data_masked[378];
  assign N348 = data_masked[506] | data_masked[442];
  assign data_o[59] = N359 | data_masked[59];
  assign N359 = N358 | data_masked[123];
  assign N358 = N357 | data_masked[187];
  assign N357 = N356 | data_masked[251];
  assign N356 = N355 | data_masked[315];
  assign N355 = N354 | data_masked[379];
  assign N354 = data_masked[507] | data_masked[443];
  assign data_o[60] = N365 | data_masked[60];
  assign N365 = N364 | data_masked[124];
  assign N364 = N363 | data_masked[188];
  assign N363 = N362 | data_masked[252];
  assign N362 = N361 | data_masked[316];
  assign N361 = N360 | data_masked[380];
  assign N360 = data_masked[508] | data_masked[444];
  assign data_o[61] = N371 | data_masked[61];
  assign N371 = N370 | data_masked[125];
  assign N370 = N369 | data_masked[189];
  assign N369 = N368 | data_masked[253];
  assign N368 = N367 | data_masked[317];
  assign N367 = N366 | data_masked[381];
  assign N366 = data_masked[509] | data_masked[445];
  assign data_o[62] = N377 | data_masked[62];
  assign N377 = N376 | data_masked[126];
  assign N376 = N375 | data_masked[190];
  assign N375 = N374 | data_masked[254];
  assign N374 = N373 | data_masked[318];
  assign N373 = N372 | data_masked[382];
  assign N372 = data_masked[510] | data_masked[446];
  assign data_o[63] = N383 | data_masked[63];
  assign N383 = N382 | data_masked[127];
  assign N382 = N381 | data_masked[191];
  assign N381 = N380 | data_masked[255];
  assign N380 = N379 | data_masked[319];
  assign N379 = N378 | data_masked[383];
  assign N378 = data_masked[511] | data_masked[447];

endmodule



module bsg_mux_00000040_00000001
(
  data_i,
  sel_i,
  data_o
);

  input [63:0] data_i;
  input [0:0] sel_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  assign data_o[63] = data_i[63];
  assign data_o[62] = data_i[62];
  assign data_o[61] = data_i[61];
  assign data_o[60] = data_i[60];
  assign data_o[59] = data_i[59];
  assign data_o[58] = data_i[58];
  assign data_o[57] = data_i[57];
  assign data_o[56] = data_i[56];
  assign data_o[55] = data_i[55];
  assign data_o[54] = data_i[54];
  assign data_o[53] = data_i[53];
  assign data_o[52] = data_i[52];
  assign data_o[51] = data_i[51];
  assign data_o[50] = data_i[50];
  assign data_o[49] = data_i[49];
  assign data_o[48] = data_i[48];
  assign data_o[47] = data_i[47];
  assign data_o[46] = data_i[46];
  assign data_o[45] = data_i[45];
  assign data_o[44] = data_i[44];
  assign data_o[43] = data_i[43];
  assign data_o[42] = data_i[42];
  assign data_o[41] = data_i[41];
  assign data_o[40] = data_i[40];
  assign data_o[39] = data_i[39];
  assign data_o[38] = data_i[38];
  assign data_o[37] = data_i[37];
  assign data_o[36] = data_i[36];
  assign data_o[35] = data_i[35];
  assign data_o[34] = data_i[34];
  assign data_o[33] = data_i[33];
  assign data_o[32] = data_i[32];
  assign data_o[31] = data_i[31];
  assign data_o[30] = data_i[30];
  assign data_o[29] = data_i[29];
  assign data_o[28] = data_i[28];
  assign data_o[27] = data_i[27];
  assign data_o[26] = data_i[26];
  assign data_o[25] = data_i[25];
  assign data_o[24] = data_i[24];
  assign data_o[23] = data_i[23];
  assign data_o[22] = data_i[22];
  assign data_o[21] = data_i[21];
  assign data_o[20] = data_i[20];
  assign data_o[19] = data_i[19];
  assign data_o[18] = data_i[18];
  assign data_o[17] = data_i[17];
  assign data_o[16] = data_i[16];
  assign data_o[15] = data_i[15];
  assign data_o[14] = data_i[14];
  assign data_o[13] = data_i[13];
  assign data_o[12] = data_i[12];
  assign data_o[11] = data_i[11];
  assign data_o[10] = data_i[10];
  assign data_o[9] = data_i[9];
  assign data_o[8] = data_i[8];
  assign data_o[7] = data_i[7];
  assign data_o[6] = data_i[6];
  assign data_o[5] = data_i[5];
  assign data_o[4] = data_i[4];
  assign data_o[3] = data_i[3];
  assign data_o[2] = data_i[2];
  assign data_o[1] = data_i[1];
  assign data_o[0] = data_i[0];

endmodule



module bsg_mem_1rw_sync_mask_write_bit_0000000f_00000040_1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [14:0] data_i;
  input [5:0] addr_i;
  input [14:0] w_mask_i;
  output [14:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [14:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_expand_bitmask_in_width_p8_expand_p1
(
  i,
  o
);

  input [7:0] i;
  output [7:0] o;
  wire [7:0] o;
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_decode_num_out_p4
(
  i,
  o
);

  input [1:0] i;
  output [3:0] o;
  wire [3:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_expand_bitmask_in_width_p4_expand_p2
(
  i,
  o
);

  input [3:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire o_7_,o_5_,o_3_,o_1_;
  assign o_7_ = i[3];
  assign o[6] = o_7_;
  assign o[7] = o_7_;
  assign o_5_ = i[2];
  assign o[4] = o_5_;
  assign o[5] = o_5_;
  assign o_3_ = i[1];
  assign o[2] = o_3_;
  assign o[3] = o_3_;
  assign o_1_ = i[0];
  assign o[0] = o_1_;
  assign o[1] = o_1_;

endmodule



module bsg_expand_bitmask_in_width_p2_expand_p4
(
  i,
  o
);

  input [1:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire o_7_,o_3_;
  assign o_7_ = i[1];
  assign o[4] = o_7_;
  assign o[5] = o_7_;
  assign o[6] = o_7_;
  assign o[7] = o_7_;
  assign o_3_ = i[0];
  assign o[0] = o_3_;
  assign o[1] = o_3_;
  assign o[2] = o_3_;
  assign o[3] = o_3_;

endmodule



module bsg_decode_num_out_p1
(
  i,
  o
);

  input [0:0] i;
  output [0:0] o;
  wire [0:0] o;
  assign o[0] = 1'b1;

endmodule



module bsg_expand_bitmask_in_width_p1_expand_p8
(
  i,
  o
);

  input [0:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire o_7_;
  assign o_7_ = i[0];
  assign o[0] = o_7_;
  assign o[1] = o_7_;
  assign o[2] = o_7_;
  assign o[3] = o_7_;
  assign o[4] = o_7_;
  assign o[5] = o_7_;
  assign o[6] = o_7_;
  assign o[7] = o_7_;

endmodule



module bsg_mux_one_hot_width_p64_els_p4
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [255:0] data_i;
  input [3:0] sel_one_hot_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127;
  wire [255:0] data_masked;
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[1];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[1];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[1];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[2];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[2];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[2];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[2];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[2];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[2];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[2];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[2];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[2];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[2];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[2];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[2];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[2];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[2];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[2];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[2];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[2];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[2];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[2];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[2];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[2];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[2];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[2];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[2];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[2];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[2];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[2];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[2];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[2];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[2];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[2];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[2];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[2];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[2];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[2];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[2];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[2];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[2];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[2];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[2];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[2];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[2];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[2];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[2];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[2];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[2];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[2];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[2];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[2];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[2];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[2];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[2];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[2];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[2];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[2];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[2];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[2];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[2];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[2];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[2];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[2];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[2];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[2];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[2];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[3];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[3];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[3];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[3];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[3];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[3];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[3];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[3];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[3];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[3];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[3];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[3];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[3];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[3];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[3];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[3];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[3];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[3];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[3];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[3];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[3];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[3];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[3];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[3];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[3];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[3];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[3];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[3];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[3];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[3];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[3];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[3];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[3];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[3];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[3];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[3];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[3];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[3];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[3];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[3];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[3];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[3];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[3];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[3];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[3];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[3];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[3];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[3];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[3];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[3];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[3];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[3];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[3];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[3];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[3];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[3];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[3];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[3];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[3];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[3];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[3];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[3];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[3];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[3];
  assign data_o[0] = N1 | data_masked[0];
  assign N1 = N0 | data_masked[64];
  assign N0 = data_masked[192] | data_masked[128];
  assign data_o[1] = N3 | data_masked[1];
  assign N3 = N2 | data_masked[65];
  assign N2 = data_masked[193] | data_masked[129];
  assign data_o[2] = N5 | data_masked[2];
  assign N5 = N4 | data_masked[66];
  assign N4 = data_masked[194] | data_masked[130];
  assign data_o[3] = N7 | data_masked[3];
  assign N7 = N6 | data_masked[67];
  assign N6 = data_masked[195] | data_masked[131];
  assign data_o[4] = N9 | data_masked[4];
  assign N9 = N8 | data_masked[68];
  assign N8 = data_masked[196] | data_masked[132];
  assign data_o[5] = N11 | data_masked[5];
  assign N11 = N10 | data_masked[69];
  assign N10 = data_masked[197] | data_masked[133];
  assign data_o[6] = N13 | data_masked[6];
  assign N13 = N12 | data_masked[70];
  assign N12 = data_masked[198] | data_masked[134];
  assign data_o[7] = N15 | data_masked[7];
  assign N15 = N14 | data_masked[71];
  assign N14 = data_masked[199] | data_masked[135];
  assign data_o[8] = N17 | data_masked[8];
  assign N17 = N16 | data_masked[72];
  assign N16 = data_masked[200] | data_masked[136];
  assign data_o[9] = N19 | data_masked[9];
  assign N19 = N18 | data_masked[73];
  assign N18 = data_masked[201] | data_masked[137];
  assign data_o[10] = N21 | data_masked[10];
  assign N21 = N20 | data_masked[74];
  assign N20 = data_masked[202] | data_masked[138];
  assign data_o[11] = N23 | data_masked[11];
  assign N23 = N22 | data_masked[75];
  assign N22 = data_masked[203] | data_masked[139];
  assign data_o[12] = N25 | data_masked[12];
  assign N25 = N24 | data_masked[76];
  assign N24 = data_masked[204] | data_masked[140];
  assign data_o[13] = N27 | data_masked[13];
  assign N27 = N26 | data_masked[77];
  assign N26 = data_masked[205] | data_masked[141];
  assign data_o[14] = N29 | data_masked[14];
  assign N29 = N28 | data_masked[78];
  assign N28 = data_masked[206] | data_masked[142];
  assign data_o[15] = N31 | data_masked[15];
  assign N31 = N30 | data_masked[79];
  assign N30 = data_masked[207] | data_masked[143];
  assign data_o[16] = N33 | data_masked[16];
  assign N33 = N32 | data_masked[80];
  assign N32 = data_masked[208] | data_masked[144];
  assign data_o[17] = N35 | data_masked[17];
  assign N35 = N34 | data_masked[81];
  assign N34 = data_masked[209] | data_masked[145];
  assign data_o[18] = N37 | data_masked[18];
  assign N37 = N36 | data_masked[82];
  assign N36 = data_masked[210] | data_masked[146];
  assign data_o[19] = N39 | data_masked[19];
  assign N39 = N38 | data_masked[83];
  assign N38 = data_masked[211] | data_masked[147];
  assign data_o[20] = N41 | data_masked[20];
  assign N41 = N40 | data_masked[84];
  assign N40 = data_masked[212] | data_masked[148];
  assign data_o[21] = N43 | data_masked[21];
  assign N43 = N42 | data_masked[85];
  assign N42 = data_masked[213] | data_masked[149];
  assign data_o[22] = N45 | data_masked[22];
  assign N45 = N44 | data_masked[86];
  assign N44 = data_masked[214] | data_masked[150];
  assign data_o[23] = N47 | data_masked[23];
  assign N47 = N46 | data_masked[87];
  assign N46 = data_masked[215] | data_masked[151];
  assign data_o[24] = N49 | data_masked[24];
  assign N49 = N48 | data_masked[88];
  assign N48 = data_masked[216] | data_masked[152];
  assign data_o[25] = N51 | data_masked[25];
  assign N51 = N50 | data_masked[89];
  assign N50 = data_masked[217] | data_masked[153];
  assign data_o[26] = N53 | data_masked[26];
  assign N53 = N52 | data_masked[90];
  assign N52 = data_masked[218] | data_masked[154];
  assign data_o[27] = N55 | data_masked[27];
  assign N55 = N54 | data_masked[91];
  assign N54 = data_masked[219] | data_masked[155];
  assign data_o[28] = N57 | data_masked[28];
  assign N57 = N56 | data_masked[92];
  assign N56 = data_masked[220] | data_masked[156];
  assign data_o[29] = N59 | data_masked[29];
  assign N59 = N58 | data_masked[93];
  assign N58 = data_masked[221] | data_masked[157];
  assign data_o[30] = N61 | data_masked[30];
  assign N61 = N60 | data_masked[94];
  assign N60 = data_masked[222] | data_masked[158];
  assign data_o[31] = N63 | data_masked[31];
  assign N63 = N62 | data_masked[95];
  assign N62 = data_masked[223] | data_masked[159];
  assign data_o[32] = N65 | data_masked[32];
  assign N65 = N64 | data_masked[96];
  assign N64 = data_masked[224] | data_masked[160];
  assign data_o[33] = N67 | data_masked[33];
  assign N67 = N66 | data_masked[97];
  assign N66 = data_masked[225] | data_masked[161];
  assign data_o[34] = N69 | data_masked[34];
  assign N69 = N68 | data_masked[98];
  assign N68 = data_masked[226] | data_masked[162];
  assign data_o[35] = N71 | data_masked[35];
  assign N71 = N70 | data_masked[99];
  assign N70 = data_masked[227] | data_masked[163];
  assign data_o[36] = N73 | data_masked[36];
  assign N73 = N72 | data_masked[100];
  assign N72 = data_masked[228] | data_masked[164];
  assign data_o[37] = N75 | data_masked[37];
  assign N75 = N74 | data_masked[101];
  assign N74 = data_masked[229] | data_masked[165];
  assign data_o[38] = N77 | data_masked[38];
  assign N77 = N76 | data_masked[102];
  assign N76 = data_masked[230] | data_masked[166];
  assign data_o[39] = N79 | data_masked[39];
  assign N79 = N78 | data_masked[103];
  assign N78 = data_masked[231] | data_masked[167];
  assign data_o[40] = N81 | data_masked[40];
  assign N81 = N80 | data_masked[104];
  assign N80 = data_masked[232] | data_masked[168];
  assign data_o[41] = N83 | data_masked[41];
  assign N83 = N82 | data_masked[105];
  assign N82 = data_masked[233] | data_masked[169];
  assign data_o[42] = N85 | data_masked[42];
  assign N85 = N84 | data_masked[106];
  assign N84 = data_masked[234] | data_masked[170];
  assign data_o[43] = N87 | data_masked[43];
  assign N87 = N86 | data_masked[107];
  assign N86 = data_masked[235] | data_masked[171];
  assign data_o[44] = N89 | data_masked[44];
  assign N89 = N88 | data_masked[108];
  assign N88 = data_masked[236] | data_masked[172];
  assign data_o[45] = N91 | data_masked[45];
  assign N91 = N90 | data_masked[109];
  assign N90 = data_masked[237] | data_masked[173];
  assign data_o[46] = N93 | data_masked[46];
  assign N93 = N92 | data_masked[110];
  assign N92 = data_masked[238] | data_masked[174];
  assign data_o[47] = N95 | data_masked[47];
  assign N95 = N94 | data_masked[111];
  assign N94 = data_masked[239] | data_masked[175];
  assign data_o[48] = N97 | data_masked[48];
  assign N97 = N96 | data_masked[112];
  assign N96 = data_masked[240] | data_masked[176];
  assign data_o[49] = N99 | data_masked[49];
  assign N99 = N98 | data_masked[113];
  assign N98 = data_masked[241] | data_masked[177];
  assign data_o[50] = N101 | data_masked[50];
  assign N101 = N100 | data_masked[114];
  assign N100 = data_masked[242] | data_masked[178];
  assign data_o[51] = N103 | data_masked[51];
  assign N103 = N102 | data_masked[115];
  assign N102 = data_masked[243] | data_masked[179];
  assign data_o[52] = N105 | data_masked[52];
  assign N105 = N104 | data_masked[116];
  assign N104 = data_masked[244] | data_masked[180];
  assign data_o[53] = N107 | data_masked[53];
  assign N107 = N106 | data_masked[117];
  assign N106 = data_masked[245] | data_masked[181];
  assign data_o[54] = N109 | data_masked[54];
  assign N109 = N108 | data_masked[118];
  assign N108 = data_masked[246] | data_masked[182];
  assign data_o[55] = N111 | data_masked[55];
  assign N111 = N110 | data_masked[119];
  assign N110 = data_masked[247] | data_masked[183];
  assign data_o[56] = N113 | data_masked[56];
  assign N113 = N112 | data_masked[120];
  assign N112 = data_masked[248] | data_masked[184];
  assign data_o[57] = N115 | data_masked[57];
  assign N115 = N114 | data_masked[121];
  assign N114 = data_masked[249] | data_masked[185];
  assign data_o[58] = N117 | data_masked[58];
  assign N117 = N116 | data_masked[122];
  assign N116 = data_masked[250] | data_masked[186];
  assign data_o[59] = N119 | data_masked[59];
  assign N119 = N118 | data_masked[123];
  assign N118 = data_masked[251] | data_masked[187];
  assign data_o[60] = N121 | data_masked[60];
  assign N121 = N120 | data_masked[124];
  assign N120 = data_masked[252] | data_masked[188];
  assign data_o[61] = N123 | data_masked[61];
  assign N123 = N122 | data_masked[125];
  assign N122 = data_masked[253] | data_masked[189];
  assign data_o[62] = N125 | data_masked[62];
  assign N125 = N124 | data_masked[126];
  assign N124 = data_masked[254] | data_masked[190];
  assign data_o[63] = N127 | data_masked[63];
  assign N127 = N126 | data_masked[127];
  assign N126 = data_masked[255] | data_masked[191];

endmodule



module bsg_mux_one_hot_00000008_4
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [31:0] data_i;
  input [3:0] sel_one_hot_i;
  output [7:0] data_o;
  wire [7:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;
  wire [31:0] data_masked;
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[1];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[1];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[1];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[1];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[1];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[1];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[1];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[1];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[2];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[2];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[2];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[2];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[2];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[2];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[2];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[2];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[3];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[3];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[3];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[3];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[3];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[3];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[3];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[3];
  assign data_o[0] = N1 | data_masked[0];
  assign N1 = N0 | data_masked[8];
  assign N0 = data_masked[24] | data_masked[16];
  assign data_o[1] = N3 | data_masked[1];
  assign N3 = N2 | data_masked[9];
  assign N2 = data_masked[25] | data_masked[17];
  assign data_o[2] = N5 | data_masked[2];
  assign N5 = N4 | data_masked[10];
  assign N4 = data_masked[26] | data_masked[18];
  assign data_o[3] = N7 | data_masked[3];
  assign N7 = N6 | data_masked[11];
  assign N6 = data_masked[27] | data_masked[19];
  assign data_o[4] = N9 | data_masked[4];
  assign N9 = N8 | data_masked[12];
  assign N8 = data_masked[28] | data_masked[20];
  assign data_o[5] = N11 | data_masked[5];
  assign N11 = N10 | data_masked[13];
  assign N10 = data_masked[29] | data_masked[21];
  assign data_o[6] = N13 | data_masked[6];
  assign N13 = N12 | data_masked[14];
  assign N12 = data_masked[30] | data_masked[22];
  assign data_o[7] = N15 | data_masked[7];
  assign N15 = N14 | data_masked[15];
  assign N14 = data_masked[31] | data_masked[23];

endmodule



module bsg_counter_up_down_max_val_p2_init_val_p0_max_step_p1
(
  clk_i,
  reset_i,
  up_i,
  down_i,
  count_o
);

  input [0:0] up_i;
  input [0:0] down_i;
  output [1:0] count_o;
  input clk_i;
  input reset_i;
  wire [1:0] count_o;
  wire N0,N1,N2,N3,N4;
  reg count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign { N2, N1 } = count_o - down_i[0];
  assign { N4, N3 } = { N2, N1 } + up_i[0];
  assign N0 = ~reset_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      count_o_1_sv2v_reg <= 1'b0;
      count_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      count_o_1_sv2v_reg <= N4;
      count_o_0_sv2v_reg <= N3;
    end 
  end


endmodule



module bsg_dff_en_width_p113
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [112:0] data_i;
  output [112:0] data_o;
  input clk_i;
  input en_i;
  wire [112:0] data_o;
  reg data_o_112_sv2v_reg,data_o_111_sv2v_reg,data_o_110_sv2v_reg,data_o_109_sv2v_reg,
  data_o_108_sv2v_reg,data_o_107_sv2v_reg,data_o_106_sv2v_reg,data_o_105_sv2v_reg,
  data_o_104_sv2v_reg,data_o_103_sv2v_reg,data_o_102_sv2v_reg,data_o_101_sv2v_reg,
  data_o_100_sv2v_reg,data_o_99_sv2v_reg,data_o_98_sv2v_reg,data_o_97_sv2v_reg,
  data_o_96_sv2v_reg,data_o_95_sv2v_reg,data_o_94_sv2v_reg,data_o_93_sv2v_reg,
  data_o_92_sv2v_reg,data_o_91_sv2v_reg,data_o_90_sv2v_reg,data_o_89_sv2v_reg,
  data_o_88_sv2v_reg,data_o_87_sv2v_reg,data_o_86_sv2v_reg,data_o_85_sv2v_reg,
  data_o_84_sv2v_reg,data_o_83_sv2v_reg,data_o_82_sv2v_reg,data_o_81_sv2v_reg,data_o_80_sv2v_reg,
  data_o_79_sv2v_reg,data_o_78_sv2v_reg,data_o_77_sv2v_reg,data_o_76_sv2v_reg,
  data_o_75_sv2v_reg,data_o_74_sv2v_reg,data_o_73_sv2v_reg,data_o_72_sv2v_reg,
  data_o_71_sv2v_reg,data_o_70_sv2v_reg,data_o_69_sv2v_reg,data_o_68_sv2v_reg,
  data_o_67_sv2v_reg,data_o_66_sv2v_reg,data_o_65_sv2v_reg,data_o_64_sv2v_reg,
  data_o_63_sv2v_reg,data_o_62_sv2v_reg,data_o_61_sv2v_reg,data_o_60_sv2v_reg,data_o_59_sv2v_reg,
  data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,data_o_55_sv2v_reg,
  data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,data_o_51_sv2v_reg,
  data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,data_o_47_sv2v_reg,
  data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,data_o_43_sv2v_reg,
  data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,
  data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,
  data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,
  data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,
  data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,
  data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,
  data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,
  data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,
  data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[112] = data_o_112_sv2v_reg;
  assign data_o[111] = data_o_111_sv2v_reg;
  assign data_o[110] = data_o_110_sv2v_reg;
  assign data_o[109] = data_o_109_sv2v_reg;
  assign data_o[108] = data_o_108_sv2v_reg;
  assign data_o[107] = data_o_107_sv2v_reg;
  assign data_o[106] = data_o_106_sv2v_reg;
  assign data_o[105] = data_o_105_sv2v_reg;
  assign data_o[104] = data_o_104_sv2v_reg;
  assign data_o[103] = data_o_103_sv2v_reg;
  assign data_o[102] = data_o_102_sv2v_reg;
  assign data_o[101] = data_o_101_sv2v_reg;
  assign data_o[100] = data_o_100_sv2v_reg;
  assign data_o[99] = data_o_99_sv2v_reg;
  assign data_o[98] = data_o_98_sv2v_reg;
  assign data_o[97] = data_o_97_sv2v_reg;
  assign data_o[96] = data_o_96_sv2v_reg;
  assign data_o[95] = data_o_95_sv2v_reg;
  assign data_o[94] = data_o_94_sv2v_reg;
  assign data_o[93] = data_o_93_sv2v_reg;
  assign data_o[92] = data_o_92_sv2v_reg;
  assign data_o[91] = data_o_91_sv2v_reg;
  assign data_o[90] = data_o_90_sv2v_reg;
  assign data_o[89] = data_o_89_sv2v_reg;
  assign data_o[88] = data_o_88_sv2v_reg;
  assign data_o[87] = data_o_87_sv2v_reg;
  assign data_o[86] = data_o_86_sv2v_reg;
  assign data_o[85] = data_o_85_sv2v_reg;
  assign data_o[84] = data_o_84_sv2v_reg;
  assign data_o[83] = data_o_83_sv2v_reg;
  assign data_o[82] = data_o_82_sv2v_reg;
  assign data_o[81] = data_o_81_sv2v_reg;
  assign data_o[80] = data_o_80_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_112_sv2v_reg <= data_i[112];
      data_o_111_sv2v_reg <= data_i[111];
      data_o_110_sv2v_reg <= data_i[110];
      data_o_109_sv2v_reg <= data_i[109];
      data_o_108_sv2v_reg <= data_i[108];
      data_o_107_sv2v_reg <= data_i[107];
      data_o_106_sv2v_reg <= data_i[106];
      data_o_105_sv2v_reg <= data_i[105];
      data_o_104_sv2v_reg <= data_i[104];
      data_o_103_sv2v_reg <= data_i[103];
      data_o_102_sv2v_reg <= data_i[102];
      data_o_101_sv2v_reg <= data_i[101];
      data_o_100_sv2v_reg <= data_i[100];
      data_o_99_sv2v_reg <= data_i[99];
      data_o_98_sv2v_reg <= data_i[98];
      data_o_97_sv2v_reg <= data_i[97];
      data_o_96_sv2v_reg <= data_i[96];
      data_o_95_sv2v_reg <= data_i[95];
      data_o_94_sv2v_reg <= data_i[94];
      data_o_93_sv2v_reg <= data_i[93];
      data_o_92_sv2v_reg <= data_i[92];
      data_o_91_sv2v_reg <= data_i[91];
      data_o_90_sv2v_reg <= data_i[90];
      data_o_89_sv2v_reg <= data_i[89];
      data_o_88_sv2v_reg <= data_i[88];
      data_o_87_sv2v_reg <= data_i[87];
      data_o_86_sv2v_reg <= data_i[86];
      data_o_85_sv2v_reg <= data_i[85];
      data_o_84_sv2v_reg <= data_i[84];
      data_o_83_sv2v_reg <= data_i[83];
      data_o_82_sv2v_reg <= data_i[82];
      data_o_81_sv2v_reg <= data_i[81];
      data_o_80_sv2v_reg <= data_i[80];
      data_o_79_sv2v_reg <= data_i[79];
      data_o_78_sv2v_reg <= data_i[78];
      data_o_77_sv2v_reg <= data_i[77];
      data_o_76_sv2v_reg <= data_i[76];
      data_o_75_sv2v_reg <= data_i[75];
      data_o_74_sv2v_reg <= data_i[74];
      data_o_73_sv2v_reg <= data_i[73];
      data_o_72_sv2v_reg <= data_i[72];
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mux_segmented_segments_p8_segment_width_p8
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [63:0] data0_i;
  input [63:0] data1_i;
  input [7:0] sel_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;
  assign data_o[7:0] = (N0)? data1_i[7:0] : 
                       (N8)? data0_i[7:0] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[15:8] = (N1)? data1_i[15:8] : 
                        (N9)? data0_i[15:8] : 1'b0;
  assign N1 = sel_i[1];
  assign data_o[23:16] = (N2)? data1_i[23:16] : 
                         (N10)? data0_i[23:16] : 1'b0;
  assign N2 = sel_i[2];
  assign data_o[31:24] = (N3)? data1_i[31:24] : 
                         (N11)? data0_i[31:24] : 1'b0;
  assign N3 = sel_i[3];
  assign data_o[39:32] = (N4)? data1_i[39:32] : 
                         (N12)? data0_i[39:32] : 1'b0;
  assign N4 = sel_i[4];
  assign data_o[47:40] = (N5)? data1_i[47:40] : 
                         (N13)? data0_i[47:40] : 1'b0;
  assign N5 = sel_i[5];
  assign data_o[55:48] = (N6)? data1_i[55:48] : 
                         (N14)? data0_i[55:48] : 1'b0;
  assign N6 = sel_i[6];
  assign data_o[63:56] = (N7)? data1_i[63:56] : 
                         (N15)? data0_i[63:56] : 1'b0;
  assign N7 = sel_i[7];
  assign N8 = ~sel_i[0];
  assign N9 = ~sel_i[1];
  assign N10 = ~sel_i[2];
  assign N11 = ~sel_i[3];
  assign N12 = ~sel_i[4];
  assign N13 = ~sel_i[5];
  assign N14 = ~sel_i[6];
  assign N15 = ~sel_i[7];

endmodule



module bsg_dff_reset_width_p72
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [71:0] data_i;
  output [71:0] data_o;
  input clk_i;
  input reset_i;
  wire [71:0] data_o;
  reg data_o_71_sv2v_reg,data_o_70_sv2v_reg,data_o_69_sv2v_reg,data_o_68_sv2v_reg,
  data_o_67_sv2v_reg,data_o_66_sv2v_reg,data_o_65_sv2v_reg,data_o_64_sv2v_reg,
  data_o_63_sv2v_reg,data_o_62_sv2v_reg,data_o_61_sv2v_reg,data_o_60_sv2v_reg,
  data_o_59_sv2v_reg,data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,
  data_o_55_sv2v_reg,data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,data_o_51_sv2v_reg,
  data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,data_o_47_sv2v_reg,
  data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,data_o_43_sv2v_reg,
  data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,
  data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,
  data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,
  data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,
  data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,
  data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,
  data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,
  data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_71_sv2v_reg <= 1'b0;
      data_o_70_sv2v_reg <= 1'b0;
      data_o_69_sv2v_reg <= 1'b0;
      data_o_68_sv2v_reg <= 1'b0;
      data_o_67_sv2v_reg <= 1'b0;
      data_o_66_sv2v_reg <= 1'b0;
      data_o_65_sv2v_reg <= 1'b0;
      data_o_64_sv2v_reg <= 1'b0;
      data_o_63_sv2v_reg <= 1'b0;
      data_o_62_sv2v_reg <= 1'b0;
      data_o_61_sv2v_reg <= 1'b0;
      data_o_60_sv2v_reg <= 1'b0;
      data_o_59_sv2v_reg <= 1'b0;
      data_o_58_sv2v_reg <= 1'b0;
      data_o_57_sv2v_reg <= 1'b0;
      data_o_56_sv2v_reg <= 1'b0;
      data_o_55_sv2v_reg <= 1'b0;
      data_o_54_sv2v_reg <= 1'b0;
      data_o_53_sv2v_reg <= 1'b0;
      data_o_52_sv2v_reg <= 1'b0;
      data_o_51_sv2v_reg <= 1'b0;
      data_o_50_sv2v_reg <= 1'b0;
      data_o_49_sv2v_reg <= 1'b0;
      data_o_48_sv2v_reg <= 1'b0;
      data_o_47_sv2v_reg <= 1'b0;
      data_o_46_sv2v_reg <= 1'b0;
      data_o_45_sv2v_reg <= 1'b0;
      data_o_44_sv2v_reg <= 1'b0;
      data_o_43_sv2v_reg <= 1'b0;
      data_o_42_sv2v_reg <= 1'b0;
      data_o_41_sv2v_reg <= 1'b0;
      data_o_40_sv2v_reg <= 1'b0;
      data_o_39_sv2v_reg <= 1'b0;
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bp_be_dcache_wbuf_00_00000040_00000008_00000200_00000080_00000014
(
  clk_i,
  reset_i,
  wbuf_entry_i,
  v_i,
  wbuf_entry_o,
  v_o,
  force_o,
  yumi_i,
  data_mem_pkt_i,
  data_mem_pkt_v_i,
  tag_mem_pkt_i,
  tag_mem_pkt_v_i,
  stat_mem_pkt_i,
  stat_mem_pkt_v_i,
  snoop_match_o,
  v_tl_i,
  addr_tl_i,
  data_tv_i,
  data_merged_o
);

  input [112:0] wbuf_entry_i;
  output [112:0] wbuf_entry_o;
  input [142:0] data_mem_pkt_i;
  input [34:0] tag_mem_pkt_i;
  input [10:0] stat_mem_pkt_i;
  input [31:0] addr_tl_i;
  input [63:0] data_tv_i;
  output [63:0] data_merged_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input data_mem_pkt_v_i;
  input tag_mem_pkt_v_i;
  input stat_mem_pkt_v_i;
  input v_tl_i;
  output v_o;
  output force_o;
  output snoop_match_o;
  wire [112:0] wbuf_entry_o,wbuf_entry_el0_r,wbuf_entry_el1_n,wbuf_entry_el1_r;
  wire [63:0] data_merged_o,el0or1_data,bypass_data_n,bypass_data_r;
  wire v_o,force_o,snoop_match_o,N0,N1,N2,N3,N4,N5,N6,N7,el0_valid,el1_valid,
  el0_enable,N8,el1_enable,mux1_sel,N9,N10,N11,N12,N13,N14,N15,N16,tag_hit0_n,tag_hit1_n,
  tag_hit2_n,_2_net__7_,_2_net__6_,_2_net__5_,_2_net__4_,_2_net__3_,_2_net__2_,
  _2_net__1_,_2_net__0_,_4_net__7_,_4_net__6_,_4_net__5_,_4_net__4_,_4_net__3_,
  _4_net__2_,_4_net__1_,_4_net__0_,N17,snoop_tag_match,N18,snoop_stat_match,N19,
  snoop_el0_match,N20,snoop_el1_match,N21,snoop_el2_match,N22,N23,N24,N25,N26,N27,N28,N29,
  N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,
  N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,
  N70,N71,N72,N73,N74,N75;
  wire [1:0] num_els_r;
  wire [7:7] tag_hit0x4,tag_hit1x4,tag_hit2x4;
  wire [7:0] bypass_mask_n,bypass_mask_r;

  bsg_counter_up_down_max_val_p2_init_val_p0_max_step_p1
  num_els_counter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .up_i(v_i),
    .down_i(yumi_i),
    .count_o(num_els_r)
  );


  bsg_dff_en_width_p113
  wbuf_entry0_reg
  (
    .clk_i(clk_i),
    .data_i(wbuf_entry_i),
    .en_i(el0_enable),
    .data_o(wbuf_entry_el0_r)
  );


  bsg_dff_en_width_p113
  wbuf_entry1_reg
  (
    .clk_i(clk_i),
    .data_i(wbuf_entry_el1_n),
    .en_i(el1_enable),
    .data_o(wbuf_entry_el1_r)
  );

  assign tag_hit0_n = addr_tl_i[31:3] == wbuf_entry_el0_r[31:3];
  assign tag_hit1_n = addr_tl_i[31:3] == wbuf_entry_el1_r[31:3];
  assign tag_hit2_n = addr_tl_i[31:3] == wbuf_entry_i[31:3];

  bsg_mux_segmented_segments_p8_segment_width_p8
  mux_segmented_merge0
  (
    .data0_i(wbuf_entry_el1_r[95:32]),
    .data1_i(wbuf_entry_el0_r[95:32]),
    .sel_i({ _2_net__7_, _2_net__6_, _2_net__5_, _2_net__4_, _2_net__3_, _2_net__2_, _2_net__1_, _2_net__0_ }),
    .data_o(el0or1_data)
  );


  bsg_mux_segmented_segments_p8_segment_width_p8
  mux_segmented_merge1
  (
    .data0_i(el0or1_data),
    .data1_i(wbuf_entry_i[95:32]),
    .sel_i({ _4_net__7_, _4_net__6_, _4_net__5_, _4_net__4_, _4_net__3_, _4_net__2_, _4_net__1_, _4_net__0_ }),
    .data_o(bypass_data_n)
  );


  bsg_dff_reset_width_p72
  bypass_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ bypass_mask_n, bypass_data_n }),
    .data_o({ bypass_mask_r, bypass_data_r })
  );


  bsg_mux_segmented_segments_p8_segment_width_p8
  bypass_mux_segmented
  (
    .data0_i(data_tv_i),
    .data1_i(bypass_data_r),
    .sel_i(bypass_mask_r),
    .data_o(data_merged_o)
  );

  assign N17 = addr_tl_i[11:6] == tag_mem_pkt_i[34:29];
  assign N18 = addr_tl_i[11:6] == stat_mem_pkt_i[10:5];
  assign N19 = wbuf_entry_el0_r[11:6] == data_mem_pkt_i[142:137];
  assign N20 = wbuf_entry_el1_r[11:6] == data_mem_pkt_i[142:137];
  assign N21 = wbuf_entry_i[11:6] == data_mem_pkt_i[142:137];
  assign N22 = ~num_els_r[1];
  assign N23 = num_els_r[0] | N22;
  assign N24 = ~N23;
  assign N11 = (N0)? v_i : 
               (N1)? 1'b1 : 1'b0;
  assign N0 = N7;
  assign N1 = num_els_r[0];
  assign N12 = (N0)? 1'b0 : 
               (N1)? N9 : 1'b0;
  assign N13 = (N0)? N8 : 
               (N1)? N10 : 1'b0;
  assign mux1_sel = (N2)? num_els_r[0] : 
                    (N3)? 1'b1 : 1'b0;
  assign N2 = N22;
  assign N3 = el0_valid;
  assign v_o = (N2)? N11 : 
               (N3)? 1'b1 : 1'b0;
  assign el1_valid = (N2)? num_els_r[0] : 
                     (N3)? 1'b1 : 1'b0;
  assign el0_enable = (N2)? N12 : 
                      (N3)? N14 : 1'b0;
  assign el1_enable = (N2)? N13 : 
                      (N3)? yumi_i : 1'b0;
  assign wbuf_entry_el1_n = (N3)? wbuf_entry_el0_r : 
                            (N4)? wbuf_entry_i : 1'b0;
  assign N4 = N15;
  assign wbuf_entry_o = (N5)? wbuf_entry_el1_r : 
                        (N6)? wbuf_entry_i : 1'b0;
  assign N5 = mux1_sel;
  assign N6 = N16;
  assign el0_valid = num_els_r[1];
  assign N7 = ~num_els_r[0];
  assign N8 = v_i & N25;
  assign N25 = ~yumi_i;
  assign N9 = v_i & N26;
  assign N26 = ~yumi_i;
  assign N10 = v_i & yumi_i;
  assign N14 = v_i & yumi_i;
  assign force_o = v_i & N24;
  assign N15 = ~el0_valid;
  assign N16 = ~mux1_sel;
  assign tag_hit0x4[7] = N27 & el0_valid;
  assign N27 = v_tl_i & tag_hit0_n;
  assign tag_hit1x4[7] = N28 & el1_valid;
  assign N28 = v_tl_i & tag_hit1_n;
  assign tag_hit2x4[7] = N29 & v_i;
  assign N29 = v_tl_i & tag_hit2_n;
  assign _2_net__7_ = tag_hit0x4[7] & wbuf_entry_el0_r[103];
  assign _2_net__6_ = tag_hit0x4[7] & wbuf_entry_el0_r[102];
  assign _2_net__5_ = tag_hit0x4[7] & wbuf_entry_el0_r[101];
  assign _2_net__4_ = tag_hit0x4[7] & wbuf_entry_el0_r[100];
  assign _2_net__3_ = tag_hit0x4[7] & wbuf_entry_el0_r[99];
  assign _2_net__2_ = tag_hit0x4[7] & wbuf_entry_el0_r[98];
  assign _2_net__1_ = tag_hit0x4[7] & wbuf_entry_el0_r[97];
  assign _2_net__0_ = tag_hit0x4[7] & wbuf_entry_el0_r[96];
  assign _4_net__7_ = tag_hit2x4[7] & wbuf_entry_i[103];
  assign _4_net__6_ = tag_hit2x4[7] & wbuf_entry_i[102];
  assign _4_net__5_ = tag_hit2x4[7] & wbuf_entry_i[101];
  assign _4_net__4_ = tag_hit2x4[7] & wbuf_entry_i[100];
  assign _4_net__3_ = tag_hit2x4[7] & wbuf_entry_i[99];
  assign _4_net__2_ = tag_hit2x4[7] & wbuf_entry_i[98];
  assign _4_net__1_ = tag_hit2x4[7] & wbuf_entry_i[97];
  assign _4_net__0_ = tag_hit2x4[7] & wbuf_entry_i[96];
  assign bypass_mask_n[7] = N32 | N33;
  assign N32 = N30 | N31;
  assign N30 = tag_hit0x4[7] & wbuf_entry_el0_r[103];
  assign N31 = tag_hit1x4[7] & wbuf_entry_el1_r[103];
  assign N33 = tag_hit2x4[7] & wbuf_entry_i[103];
  assign bypass_mask_n[6] = N36 | N37;
  assign N36 = N34 | N35;
  assign N34 = tag_hit0x4[7] & wbuf_entry_el0_r[102];
  assign N35 = tag_hit1x4[7] & wbuf_entry_el1_r[102];
  assign N37 = tag_hit2x4[7] & wbuf_entry_i[102];
  assign bypass_mask_n[5] = N40 | N41;
  assign N40 = N38 | N39;
  assign N38 = tag_hit0x4[7] & wbuf_entry_el0_r[101];
  assign N39 = tag_hit1x4[7] & wbuf_entry_el1_r[101];
  assign N41 = tag_hit2x4[7] & wbuf_entry_i[101];
  assign bypass_mask_n[4] = N44 | N45;
  assign N44 = N42 | N43;
  assign N42 = tag_hit0x4[7] & wbuf_entry_el0_r[100];
  assign N43 = tag_hit1x4[7] & wbuf_entry_el1_r[100];
  assign N45 = tag_hit2x4[7] & wbuf_entry_i[100];
  assign bypass_mask_n[3] = N48 | N49;
  assign N48 = N46 | N47;
  assign N46 = tag_hit0x4[7] & wbuf_entry_el0_r[99];
  assign N47 = tag_hit1x4[7] & wbuf_entry_el1_r[99];
  assign N49 = tag_hit2x4[7] & wbuf_entry_i[99];
  assign bypass_mask_n[2] = N52 | N53;
  assign N52 = N50 | N51;
  assign N50 = tag_hit0x4[7] & wbuf_entry_el0_r[98];
  assign N51 = tag_hit1x4[7] & wbuf_entry_el1_r[98];
  assign N53 = tag_hit2x4[7] & wbuf_entry_i[98];
  assign bypass_mask_n[1] = N56 | N57;
  assign N56 = N54 | N55;
  assign N54 = tag_hit0x4[7] & wbuf_entry_el0_r[97];
  assign N55 = tag_hit1x4[7] & wbuf_entry_el1_r[97];
  assign N57 = tag_hit2x4[7] & wbuf_entry_i[97];
  assign bypass_mask_n[0] = N60 | N61;
  assign N60 = N58 | N59;
  assign N58 = tag_hit0x4[7] & wbuf_entry_el0_r[96];
  assign N59 = tag_hit1x4[7] & wbuf_entry_el1_r[96];
  assign N61 = tag_hit2x4[7] & wbuf_entry_i[96];
  assign snoop_tag_match = N62 & N17;
  assign N62 = v_tl_i & tag_mem_pkt_v_i;
  assign snoop_stat_match = N63 & N18;
  assign N63 = v_tl_i & stat_mem_pkt_v_i;
  assign snoop_el0_match = N66 & N19;
  assign N66 = N65 & data_mem_pkt_v_i;
  assign N65 = el0_valid & N64;
  assign N64 = ~wbuf_entry_i[112];
  assign snoop_el1_match = N69 & N20;
  assign N69 = N68 & data_mem_pkt_v_i;
  assign N68 = el1_valid & N67;
  assign N67 = ~wbuf_entry_el1_r[112];
  assign snoop_el2_match = N72 & N21;
  assign N72 = N71 & data_mem_pkt_v_i;
  assign N71 = v_i & N70;
  assign N70 = ~wbuf_entry_i[112];
  assign snoop_match_o = N75 | snoop_el2_match;
  assign N75 = N74 | snoop_el1_match;
  assign N74 = N73 | snoop_el0_match;
  assign N73 = snoop_tag_match | snoop_stat_match;

endmodule



module bsg_dff_0000000c
(
  clk_i,
  data_i,
  data_o
);

  input [11:0] data_i;
  output [11:0] data_o;
  input clk_i;
  wire [11:0] data_o;
  reg data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,
  data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_rotate_left_00000008
(
  data_i,
  rot_i,
  o
);

  input [7:0] data_i;
  input [2:0] rot_i;
  output [7:0] o;
  wire [7:0] o;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7;
  assign { o, sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7 } = { data_i, data_i[7:1] } << rot_i;

endmodule



module bsg_rotate_left_00000080
(
  data_i,
  rot_i,
  o
);

  input [127:0] data_i;
  input [6:0] rot_i;
  output [127:0] o;
  wire [127:0] o;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,
  sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,
  sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,sv2v_dc_21,sv2v_dc_22,
  sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,sv2v_dc_27,sv2v_dc_28,sv2v_dc_29,
  sv2v_dc_30,sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,sv2v_dc_34,sv2v_dc_35,sv2v_dc_36,sv2v_dc_37,
  sv2v_dc_38,sv2v_dc_39,sv2v_dc_40,sv2v_dc_41,sv2v_dc_42,sv2v_dc_43,sv2v_dc_44,
  sv2v_dc_45,sv2v_dc_46,sv2v_dc_47,sv2v_dc_48,sv2v_dc_49,sv2v_dc_50,sv2v_dc_51,
  sv2v_dc_52,sv2v_dc_53,sv2v_dc_54,sv2v_dc_55,sv2v_dc_56,sv2v_dc_57,sv2v_dc_58,sv2v_dc_59,
  sv2v_dc_60,sv2v_dc_61,sv2v_dc_62,sv2v_dc_63,sv2v_dc_64,sv2v_dc_65,sv2v_dc_66,
  sv2v_dc_67,sv2v_dc_68,sv2v_dc_69,sv2v_dc_70,sv2v_dc_71,sv2v_dc_72,sv2v_dc_73,
  sv2v_dc_74,sv2v_dc_75,sv2v_dc_76,sv2v_dc_77,sv2v_dc_78,sv2v_dc_79,sv2v_dc_80,
  sv2v_dc_81,sv2v_dc_82,sv2v_dc_83,sv2v_dc_84,sv2v_dc_85,sv2v_dc_86,sv2v_dc_87,sv2v_dc_88,
  sv2v_dc_89,sv2v_dc_90,sv2v_dc_91,sv2v_dc_92,sv2v_dc_93,sv2v_dc_94,sv2v_dc_95,
  sv2v_dc_96,sv2v_dc_97,sv2v_dc_98,sv2v_dc_99,sv2v_dc_100,sv2v_dc_101,sv2v_dc_102,
  sv2v_dc_103,sv2v_dc_104,sv2v_dc_105,sv2v_dc_106,sv2v_dc_107,sv2v_dc_108,sv2v_dc_109,
  sv2v_dc_110,sv2v_dc_111,sv2v_dc_112,sv2v_dc_113,sv2v_dc_114,sv2v_dc_115,
  sv2v_dc_116,sv2v_dc_117,sv2v_dc_118,sv2v_dc_119,sv2v_dc_120,sv2v_dc_121,sv2v_dc_122,
  sv2v_dc_123,sv2v_dc_124,sv2v_dc_125,sv2v_dc_126,sv2v_dc_127;
  assign { o, sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36, sv2v_dc_37, sv2v_dc_38, sv2v_dc_39, sv2v_dc_40, sv2v_dc_41, sv2v_dc_42, sv2v_dc_43, sv2v_dc_44, sv2v_dc_45, sv2v_dc_46, sv2v_dc_47, sv2v_dc_48, sv2v_dc_49, sv2v_dc_50, sv2v_dc_51, sv2v_dc_52, sv2v_dc_53, sv2v_dc_54, sv2v_dc_55, sv2v_dc_56, sv2v_dc_57, sv2v_dc_58, sv2v_dc_59, sv2v_dc_60, sv2v_dc_61, sv2v_dc_62, sv2v_dc_63, sv2v_dc_64, sv2v_dc_65, sv2v_dc_66, sv2v_dc_67, sv2v_dc_68, sv2v_dc_69, sv2v_dc_70, sv2v_dc_71, sv2v_dc_72, sv2v_dc_73, sv2v_dc_74, sv2v_dc_75, sv2v_dc_76, sv2v_dc_77, sv2v_dc_78, sv2v_dc_79, sv2v_dc_80, sv2v_dc_81, sv2v_dc_82, sv2v_dc_83, sv2v_dc_84, sv2v_dc_85, sv2v_dc_86, sv2v_dc_87, sv2v_dc_88, sv2v_dc_89, sv2v_dc_90, sv2v_dc_91, sv2v_dc_92, sv2v_dc_93, sv2v_dc_94, sv2v_dc_95, sv2v_dc_96, sv2v_dc_97, sv2v_dc_98, sv2v_dc_99, sv2v_dc_100, sv2v_dc_101, sv2v_dc_102, sv2v_dc_103, sv2v_dc_104, sv2v_dc_105, sv2v_dc_106, sv2v_dc_107, sv2v_dc_108, sv2v_dc_109, sv2v_dc_110, sv2v_dc_111, sv2v_dc_112, sv2v_dc_113, sv2v_dc_114, sv2v_dc_115, sv2v_dc_116, sv2v_dc_117, sv2v_dc_118, sv2v_dc_119, sv2v_dc_120, sv2v_dc_121, sv2v_dc_122, sv2v_dc_123, sv2v_dc_124, sv2v_dc_125, sv2v_dc_126, sv2v_dc_127 } = { data_i, data_i[127:1] } << rot_i;

endmodule



module bsg_rotate_right_00000200
(
  data_i,
  rot_i,
  o
);

  input [511:0] data_i;
  input [8:0] rot_i;
  output [511:0] o;
  wire [511:0] o;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,
  sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,
  sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,sv2v_dc_21,sv2v_dc_22,
  sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,sv2v_dc_27,sv2v_dc_28,sv2v_dc_29,
  sv2v_dc_30,sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,sv2v_dc_34,sv2v_dc_35,sv2v_dc_36,sv2v_dc_37,
  sv2v_dc_38,sv2v_dc_39,sv2v_dc_40,sv2v_dc_41,sv2v_dc_42,sv2v_dc_43,sv2v_dc_44,
  sv2v_dc_45,sv2v_dc_46,sv2v_dc_47,sv2v_dc_48,sv2v_dc_49,sv2v_dc_50,sv2v_dc_51,
  sv2v_dc_52,sv2v_dc_53,sv2v_dc_54,sv2v_dc_55,sv2v_dc_56,sv2v_dc_57,sv2v_dc_58,sv2v_dc_59,
  sv2v_dc_60,sv2v_dc_61,sv2v_dc_62,sv2v_dc_63,sv2v_dc_64,sv2v_dc_65,sv2v_dc_66,
  sv2v_dc_67,sv2v_dc_68,sv2v_dc_69,sv2v_dc_70,sv2v_dc_71,sv2v_dc_72,sv2v_dc_73,
  sv2v_dc_74,sv2v_dc_75,sv2v_dc_76,sv2v_dc_77,sv2v_dc_78,sv2v_dc_79,sv2v_dc_80,
  sv2v_dc_81,sv2v_dc_82,sv2v_dc_83,sv2v_dc_84,sv2v_dc_85,sv2v_dc_86,sv2v_dc_87,sv2v_dc_88,
  sv2v_dc_89,sv2v_dc_90,sv2v_dc_91,sv2v_dc_92,sv2v_dc_93,sv2v_dc_94,sv2v_dc_95,
  sv2v_dc_96,sv2v_dc_97,sv2v_dc_98,sv2v_dc_99,sv2v_dc_100,sv2v_dc_101,sv2v_dc_102,
  sv2v_dc_103,sv2v_dc_104,sv2v_dc_105,sv2v_dc_106,sv2v_dc_107,sv2v_dc_108,sv2v_dc_109,
  sv2v_dc_110,sv2v_dc_111,sv2v_dc_112,sv2v_dc_113,sv2v_dc_114,sv2v_dc_115,
  sv2v_dc_116,sv2v_dc_117,sv2v_dc_118,sv2v_dc_119,sv2v_dc_120,sv2v_dc_121,sv2v_dc_122,
  sv2v_dc_123,sv2v_dc_124,sv2v_dc_125,sv2v_dc_126,sv2v_dc_127,sv2v_dc_128,sv2v_dc_129,
  sv2v_dc_130,sv2v_dc_131,sv2v_dc_132,sv2v_dc_133,sv2v_dc_134,sv2v_dc_135,
  sv2v_dc_136,sv2v_dc_137,sv2v_dc_138,sv2v_dc_139,sv2v_dc_140,sv2v_dc_141,sv2v_dc_142,
  sv2v_dc_143,sv2v_dc_144,sv2v_dc_145,sv2v_dc_146,sv2v_dc_147,sv2v_dc_148,sv2v_dc_149,
  sv2v_dc_150,sv2v_dc_151,sv2v_dc_152,sv2v_dc_153,sv2v_dc_154,sv2v_dc_155,
  sv2v_dc_156,sv2v_dc_157,sv2v_dc_158,sv2v_dc_159,sv2v_dc_160,sv2v_dc_161,sv2v_dc_162,
  sv2v_dc_163,sv2v_dc_164,sv2v_dc_165,sv2v_dc_166,sv2v_dc_167,sv2v_dc_168,sv2v_dc_169,
  sv2v_dc_170,sv2v_dc_171,sv2v_dc_172,sv2v_dc_173,sv2v_dc_174,sv2v_dc_175,
  sv2v_dc_176,sv2v_dc_177,sv2v_dc_178,sv2v_dc_179,sv2v_dc_180,sv2v_dc_181,sv2v_dc_182,
  sv2v_dc_183,sv2v_dc_184,sv2v_dc_185,sv2v_dc_186,sv2v_dc_187,sv2v_dc_188,sv2v_dc_189,
  sv2v_dc_190,sv2v_dc_191,sv2v_dc_192,sv2v_dc_193,sv2v_dc_194,sv2v_dc_195,
  sv2v_dc_196,sv2v_dc_197,sv2v_dc_198,sv2v_dc_199,sv2v_dc_200,sv2v_dc_201,sv2v_dc_202,
  sv2v_dc_203,sv2v_dc_204,sv2v_dc_205,sv2v_dc_206,sv2v_dc_207,sv2v_dc_208,sv2v_dc_209,
  sv2v_dc_210,sv2v_dc_211,sv2v_dc_212,sv2v_dc_213,sv2v_dc_214,sv2v_dc_215,
  sv2v_dc_216,sv2v_dc_217,sv2v_dc_218,sv2v_dc_219,sv2v_dc_220,sv2v_dc_221,sv2v_dc_222,
  sv2v_dc_223,sv2v_dc_224,sv2v_dc_225,sv2v_dc_226,sv2v_dc_227,sv2v_dc_228,sv2v_dc_229,
  sv2v_dc_230,sv2v_dc_231,sv2v_dc_232,sv2v_dc_233,sv2v_dc_234,sv2v_dc_235,
  sv2v_dc_236,sv2v_dc_237,sv2v_dc_238,sv2v_dc_239,sv2v_dc_240,sv2v_dc_241,sv2v_dc_242,
  sv2v_dc_243,sv2v_dc_244,sv2v_dc_245,sv2v_dc_246,sv2v_dc_247,sv2v_dc_248,sv2v_dc_249,
  sv2v_dc_250,sv2v_dc_251,sv2v_dc_252,sv2v_dc_253,sv2v_dc_254,sv2v_dc_255,
  sv2v_dc_256,sv2v_dc_257,sv2v_dc_258,sv2v_dc_259,sv2v_dc_260,sv2v_dc_261,sv2v_dc_262,
  sv2v_dc_263,sv2v_dc_264,sv2v_dc_265,sv2v_dc_266,sv2v_dc_267,sv2v_dc_268,sv2v_dc_269,
  sv2v_dc_270,sv2v_dc_271,sv2v_dc_272,sv2v_dc_273,sv2v_dc_274,sv2v_dc_275,
  sv2v_dc_276,sv2v_dc_277,sv2v_dc_278,sv2v_dc_279,sv2v_dc_280,sv2v_dc_281,sv2v_dc_282,
  sv2v_dc_283,sv2v_dc_284,sv2v_dc_285,sv2v_dc_286,sv2v_dc_287,sv2v_dc_288,sv2v_dc_289,
  sv2v_dc_290,sv2v_dc_291,sv2v_dc_292,sv2v_dc_293,sv2v_dc_294,sv2v_dc_295,
  sv2v_dc_296,sv2v_dc_297,sv2v_dc_298,sv2v_dc_299,sv2v_dc_300,sv2v_dc_301,sv2v_dc_302,
  sv2v_dc_303,sv2v_dc_304,sv2v_dc_305,sv2v_dc_306,sv2v_dc_307,sv2v_dc_308,sv2v_dc_309,
  sv2v_dc_310,sv2v_dc_311,sv2v_dc_312,sv2v_dc_313,sv2v_dc_314,sv2v_dc_315,
  sv2v_dc_316,sv2v_dc_317,sv2v_dc_318,sv2v_dc_319,sv2v_dc_320,sv2v_dc_321,sv2v_dc_322,
  sv2v_dc_323,sv2v_dc_324,sv2v_dc_325,sv2v_dc_326,sv2v_dc_327,sv2v_dc_328,sv2v_dc_329,
  sv2v_dc_330,sv2v_dc_331,sv2v_dc_332,sv2v_dc_333,sv2v_dc_334,sv2v_dc_335,
  sv2v_dc_336,sv2v_dc_337,sv2v_dc_338,sv2v_dc_339,sv2v_dc_340,sv2v_dc_341,sv2v_dc_342,
  sv2v_dc_343,sv2v_dc_344,sv2v_dc_345,sv2v_dc_346,sv2v_dc_347,sv2v_dc_348,sv2v_dc_349,
  sv2v_dc_350,sv2v_dc_351,sv2v_dc_352,sv2v_dc_353,sv2v_dc_354,sv2v_dc_355,
  sv2v_dc_356,sv2v_dc_357,sv2v_dc_358,sv2v_dc_359,sv2v_dc_360,sv2v_dc_361,sv2v_dc_362,
  sv2v_dc_363,sv2v_dc_364,sv2v_dc_365,sv2v_dc_366,sv2v_dc_367,sv2v_dc_368,sv2v_dc_369,
  sv2v_dc_370,sv2v_dc_371,sv2v_dc_372,sv2v_dc_373,sv2v_dc_374,sv2v_dc_375,
  sv2v_dc_376,sv2v_dc_377,sv2v_dc_378,sv2v_dc_379,sv2v_dc_380,sv2v_dc_381,sv2v_dc_382,
  sv2v_dc_383,sv2v_dc_384,sv2v_dc_385,sv2v_dc_386,sv2v_dc_387,sv2v_dc_388,sv2v_dc_389,
  sv2v_dc_390,sv2v_dc_391,sv2v_dc_392,sv2v_dc_393,sv2v_dc_394,sv2v_dc_395,
  sv2v_dc_396,sv2v_dc_397,sv2v_dc_398,sv2v_dc_399,sv2v_dc_400,sv2v_dc_401,sv2v_dc_402,
  sv2v_dc_403,sv2v_dc_404,sv2v_dc_405,sv2v_dc_406,sv2v_dc_407,sv2v_dc_408,sv2v_dc_409,
  sv2v_dc_410,sv2v_dc_411,sv2v_dc_412,sv2v_dc_413,sv2v_dc_414,sv2v_dc_415,
  sv2v_dc_416,sv2v_dc_417,sv2v_dc_418,sv2v_dc_419,sv2v_dc_420,sv2v_dc_421,sv2v_dc_422,
  sv2v_dc_423,sv2v_dc_424,sv2v_dc_425,sv2v_dc_426,sv2v_dc_427,sv2v_dc_428,sv2v_dc_429,
  sv2v_dc_430,sv2v_dc_431,sv2v_dc_432,sv2v_dc_433,sv2v_dc_434,sv2v_dc_435,
  sv2v_dc_436,sv2v_dc_437,sv2v_dc_438,sv2v_dc_439,sv2v_dc_440,sv2v_dc_441,sv2v_dc_442,
  sv2v_dc_443,sv2v_dc_444,sv2v_dc_445,sv2v_dc_446,sv2v_dc_447,sv2v_dc_448,sv2v_dc_449,
  sv2v_dc_450,sv2v_dc_451,sv2v_dc_452,sv2v_dc_453,sv2v_dc_454,sv2v_dc_455,
  sv2v_dc_456,sv2v_dc_457,sv2v_dc_458,sv2v_dc_459,sv2v_dc_460,sv2v_dc_461,sv2v_dc_462,
  sv2v_dc_463,sv2v_dc_464,sv2v_dc_465,sv2v_dc_466,sv2v_dc_467,sv2v_dc_468,sv2v_dc_469,
  sv2v_dc_470,sv2v_dc_471,sv2v_dc_472,sv2v_dc_473,sv2v_dc_474,sv2v_dc_475,
  sv2v_dc_476,sv2v_dc_477,sv2v_dc_478,sv2v_dc_479,sv2v_dc_480,sv2v_dc_481,sv2v_dc_482,
  sv2v_dc_483,sv2v_dc_484,sv2v_dc_485,sv2v_dc_486,sv2v_dc_487,sv2v_dc_488,sv2v_dc_489,
  sv2v_dc_490,sv2v_dc_491,sv2v_dc_492,sv2v_dc_493,sv2v_dc_494,sv2v_dc_495,
  sv2v_dc_496,sv2v_dc_497,sv2v_dc_498,sv2v_dc_499,sv2v_dc_500,sv2v_dc_501,sv2v_dc_502,
  sv2v_dc_503,sv2v_dc_504,sv2v_dc_505,sv2v_dc_506,sv2v_dc_507,sv2v_dc_508,sv2v_dc_509,
  sv2v_dc_510,sv2v_dc_511;
  assign { sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36, sv2v_dc_37, sv2v_dc_38, sv2v_dc_39, sv2v_dc_40, sv2v_dc_41, sv2v_dc_42, sv2v_dc_43, sv2v_dc_44, sv2v_dc_45, sv2v_dc_46, sv2v_dc_47, sv2v_dc_48, sv2v_dc_49, sv2v_dc_50, sv2v_dc_51, sv2v_dc_52, sv2v_dc_53, sv2v_dc_54, sv2v_dc_55, sv2v_dc_56, sv2v_dc_57, sv2v_dc_58, sv2v_dc_59, sv2v_dc_60, sv2v_dc_61, sv2v_dc_62, sv2v_dc_63, sv2v_dc_64, sv2v_dc_65, sv2v_dc_66, sv2v_dc_67, sv2v_dc_68, sv2v_dc_69, sv2v_dc_70, sv2v_dc_71, sv2v_dc_72, sv2v_dc_73, sv2v_dc_74, sv2v_dc_75, sv2v_dc_76, sv2v_dc_77, sv2v_dc_78, sv2v_dc_79, sv2v_dc_80, sv2v_dc_81, sv2v_dc_82, sv2v_dc_83, sv2v_dc_84, sv2v_dc_85, sv2v_dc_86, sv2v_dc_87, sv2v_dc_88, sv2v_dc_89, sv2v_dc_90, sv2v_dc_91, sv2v_dc_92, sv2v_dc_93, sv2v_dc_94, sv2v_dc_95, sv2v_dc_96, sv2v_dc_97, sv2v_dc_98, sv2v_dc_99, sv2v_dc_100, sv2v_dc_101, sv2v_dc_102, sv2v_dc_103, sv2v_dc_104, sv2v_dc_105, sv2v_dc_106, sv2v_dc_107, sv2v_dc_108, sv2v_dc_109, sv2v_dc_110, sv2v_dc_111, sv2v_dc_112, sv2v_dc_113, sv2v_dc_114, sv2v_dc_115, sv2v_dc_116, sv2v_dc_117, sv2v_dc_118, sv2v_dc_119, sv2v_dc_120, sv2v_dc_121, sv2v_dc_122, sv2v_dc_123, sv2v_dc_124, sv2v_dc_125, sv2v_dc_126, sv2v_dc_127, sv2v_dc_128, sv2v_dc_129, sv2v_dc_130, sv2v_dc_131, sv2v_dc_132, sv2v_dc_133, sv2v_dc_134, sv2v_dc_135, sv2v_dc_136, sv2v_dc_137, sv2v_dc_138, sv2v_dc_139, sv2v_dc_140, sv2v_dc_141, sv2v_dc_142, sv2v_dc_143, sv2v_dc_144, sv2v_dc_145, sv2v_dc_146, sv2v_dc_147, sv2v_dc_148, sv2v_dc_149, sv2v_dc_150, sv2v_dc_151, sv2v_dc_152, sv2v_dc_153, sv2v_dc_154, sv2v_dc_155, sv2v_dc_156, sv2v_dc_157, sv2v_dc_158, sv2v_dc_159, sv2v_dc_160, sv2v_dc_161, sv2v_dc_162, sv2v_dc_163, sv2v_dc_164, sv2v_dc_165, sv2v_dc_166, sv2v_dc_167, sv2v_dc_168, sv2v_dc_169, sv2v_dc_170, sv2v_dc_171, sv2v_dc_172, sv2v_dc_173, sv2v_dc_174, sv2v_dc_175, sv2v_dc_176, sv2v_dc_177, sv2v_dc_178, sv2v_dc_179, sv2v_dc_180, sv2v_dc_181, sv2v_dc_182, sv2v_dc_183, sv2v_dc_184, sv2v_dc_185, sv2v_dc_186, sv2v_dc_187, sv2v_dc_188, sv2v_dc_189, sv2v_dc_190, sv2v_dc_191, sv2v_dc_192, sv2v_dc_193, sv2v_dc_194, sv2v_dc_195, sv2v_dc_196, sv2v_dc_197, sv2v_dc_198, sv2v_dc_199, sv2v_dc_200, sv2v_dc_201, sv2v_dc_202, sv2v_dc_203, sv2v_dc_204, sv2v_dc_205, sv2v_dc_206, sv2v_dc_207, sv2v_dc_208, sv2v_dc_209, sv2v_dc_210, sv2v_dc_211, sv2v_dc_212, sv2v_dc_213, sv2v_dc_214, sv2v_dc_215, sv2v_dc_216, sv2v_dc_217, sv2v_dc_218, sv2v_dc_219, sv2v_dc_220, sv2v_dc_221, sv2v_dc_222, sv2v_dc_223, sv2v_dc_224, sv2v_dc_225, sv2v_dc_226, sv2v_dc_227, sv2v_dc_228, sv2v_dc_229, sv2v_dc_230, sv2v_dc_231, sv2v_dc_232, sv2v_dc_233, sv2v_dc_234, sv2v_dc_235, sv2v_dc_236, sv2v_dc_237, sv2v_dc_238, sv2v_dc_239, sv2v_dc_240, sv2v_dc_241, sv2v_dc_242, sv2v_dc_243, sv2v_dc_244, sv2v_dc_245, sv2v_dc_246, sv2v_dc_247, sv2v_dc_248, sv2v_dc_249, sv2v_dc_250, sv2v_dc_251, sv2v_dc_252, sv2v_dc_253, sv2v_dc_254, sv2v_dc_255, sv2v_dc_256, sv2v_dc_257, sv2v_dc_258, sv2v_dc_259, sv2v_dc_260, sv2v_dc_261, sv2v_dc_262, sv2v_dc_263, sv2v_dc_264, sv2v_dc_265, sv2v_dc_266, sv2v_dc_267, sv2v_dc_268, sv2v_dc_269, sv2v_dc_270, sv2v_dc_271, sv2v_dc_272, sv2v_dc_273, sv2v_dc_274, sv2v_dc_275, sv2v_dc_276, sv2v_dc_277, sv2v_dc_278, sv2v_dc_279, sv2v_dc_280, sv2v_dc_281, sv2v_dc_282, sv2v_dc_283, sv2v_dc_284, sv2v_dc_285, sv2v_dc_286, sv2v_dc_287, sv2v_dc_288, sv2v_dc_289, sv2v_dc_290, sv2v_dc_291, sv2v_dc_292, sv2v_dc_293, sv2v_dc_294, sv2v_dc_295, sv2v_dc_296, sv2v_dc_297, sv2v_dc_298, sv2v_dc_299, sv2v_dc_300, sv2v_dc_301, sv2v_dc_302, sv2v_dc_303, sv2v_dc_304, sv2v_dc_305, sv2v_dc_306, sv2v_dc_307, sv2v_dc_308, sv2v_dc_309, sv2v_dc_310, sv2v_dc_311, sv2v_dc_312, sv2v_dc_313, sv2v_dc_314, sv2v_dc_315, sv2v_dc_316, sv2v_dc_317, sv2v_dc_318, sv2v_dc_319, sv2v_dc_320, sv2v_dc_321, sv2v_dc_322, sv2v_dc_323, sv2v_dc_324, sv2v_dc_325, sv2v_dc_326, sv2v_dc_327, sv2v_dc_328, sv2v_dc_329, sv2v_dc_330, sv2v_dc_331, sv2v_dc_332, sv2v_dc_333, sv2v_dc_334, sv2v_dc_335, sv2v_dc_336, sv2v_dc_337, sv2v_dc_338, sv2v_dc_339, sv2v_dc_340, sv2v_dc_341, sv2v_dc_342, sv2v_dc_343, sv2v_dc_344, sv2v_dc_345, sv2v_dc_346, sv2v_dc_347, sv2v_dc_348, sv2v_dc_349, sv2v_dc_350, sv2v_dc_351, sv2v_dc_352, sv2v_dc_353, sv2v_dc_354, sv2v_dc_355, sv2v_dc_356, sv2v_dc_357, sv2v_dc_358, sv2v_dc_359, sv2v_dc_360, sv2v_dc_361, sv2v_dc_362, sv2v_dc_363, sv2v_dc_364, sv2v_dc_365, sv2v_dc_366, sv2v_dc_367, sv2v_dc_368, sv2v_dc_369, sv2v_dc_370, sv2v_dc_371, sv2v_dc_372, sv2v_dc_373, sv2v_dc_374, sv2v_dc_375, sv2v_dc_376, sv2v_dc_377, sv2v_dc_378, sv2v_dc_379, sv2v_dc_380, sv2v_dc_381, sv2v_dc_382, sv2v_dc_383, sv2v_dc_384, sv2v_dc_385, sv2v_dc_386, sv2v_dc_387, sv2v_dc_388, sv2v_dc_389, sv2v_dc_390, sv2v_dc_391, sv2v_dc_392, sv2v_dc_393, sv2v_dc_394, sv2v_dc_395, sv2v_dc_396, sv2v_dc_397, sv2v_dc_398, sv2v_dc_399, sv2v_dc_400, sv2v_dc_401, sv2v_dc_402, sv2v_dc_403, sv2v_dc_404, sv2v_dc_405, sv2v_dc_406, sv2v_dc_407, sv2v_dc_408, sv2v_dc_409, sv2v_dc_410, sv2v_dc_411, sv2v_dc_412, sv2v_dc_413, sv2v_dc_414, sv2v_dc_415, sv2v_dc_416, sv2v_dc_417, sv2v_dc_418, sv2v_dc_419, sv2v_dc_420, sv2v_dc_421, sv2v_dc_422, sv2v_dc_423, sv2v_dc_424, sv2v_dc_425, sv2v_dc_426, sv2v_dc_427, sv2v_dc_428, sv2v_dc_429, sv2v_dc_430, sv2v_dc_431, sv2v_dc_432, sv2v_dc_433, sv2v_dc_434, sv2v_dc_435, sv2v_dc_436, sv2v_dc_437, sv2v_dc_438, sv2v_dc_439, sv2v_dc_440, sv2v_dc_441, sv2v_dc_442, sv2v_dc_443, sv2v_dc_444, sv2v_dc_445, sv2v_dc_446, sv2v_dc_447, sv2v_dc_448, sv2v_dc_449, sv2v_dc_450, sv2v_dc_451, sv2v_dc_452, sv2v_dc_453, sv2v_dc_454, sv2v_dc_455, sv2v_dc_456, sv2v_dc_457, sv2v_dc_458, sv2v_dc_459, sv2v_dc_460, sv2v_dc_461, sv2v_dc_462, sv2v_dc_463, sv2v_dc_464, sv2v_dc_465, sv2v_dc_466, sv2v_dc_467, sv2v_dc_468, sv2v_dc_469, sv2v_dc_470, sv2v_dc_471, sv2v_dc_472, sv2v_dc_473, sv2v_dc_474, sv2v_dc_475, sv2v_dc_476, sv2v_dc_477, sv2v_dc_478, sv2v_dc_479, sv2v_dc_480, sv2v_dc_481, sv2v_dc_482, sv2v_dc_483, sv2v_dc_484, sv2v_dc_485, sv2v_dc_486, sv2v_dc_487, sv2v_dc_488, sv2v_dc_489, sv2v_dc_490, sv2v_dc_491, sv2v_dc_492, sv2v_dc_493, sv2v_dc_494, sv2v_dc_495, sv2v_dc_496, sv2v_dc_497, sv2v_dc_498, sv2v_dc_499, sv2v_dc_500, sv2v_dc_501, sv2v_dc_502, sv2v_dc_503, sv2v_dc_504, sv2v_dc_505, sv2v_dc_506, sv2v_dc_507, sv2v_dc_508, sv2v_dc_509, sv2v_dc_510, sv2v_dc_511, o } = { data_i[510:0], data_i } >> rot_i;

endmodule



module bsg_decode_with_v_00000008
(
  i,
  v_i,
  o
);

  input [2:0] i;
  output [7:0] o;
  input v_i;
  wire [7:0] o,lo;

  bsg_decode_00000008
  bd
  (
    .i(i),
    .o(lo)
  );

  assign o[7] = v_i & lo[7];
  assign o[6] = v_i & lo[6];
  assign o[5] = v_i & lo[5];
  assign o[4] = v_i & lo[4];
  assign o[3] = v_i & lo[3];
  assign o[2] = v_i & lo[2];
  assign o[1] = v_i & lo[1];
  assign o[0] = v_i & lo[0];

endmodule



module bsg_dff_reset_set_clear_width_p1_clear_over_set_p1
(
  clk_i,
  reset_i,
  set_i,
  clear_i,
  data_o
);

  input [0:0] set_i;
  input [0:0] clear_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  wire [0:0] data_o;
  wire N0,N1,N2;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N0 = N1 & N2;
  assign N1 = data_o[0] | set_i[0];
  assign N2 = ~clear_i[0];

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_0_sv2v_reg <= N0;
    end 
  end


endmodule



module bsg_dff_en_0000001a
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [25:0] data_i;
  output [25:0] data_o;
  input clk_i;
  input en_i;
  wire [25:0] data_o;
  reg data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,
  data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,
  data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_counter_clear_up_max_val_p15_init_val_p0_disable_overflow_warning_p1
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [3:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire [3:0] count_o;
  wire N0,N1,N4,N5,N6,N8,N9,N10,N11,N12,N13,N14,N15,N16,N2,N3,N7,N30,N17;
  reg count_o_3_sv2v_reg,count_o_2_sv2v_reg,count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[3] = count_o_3_sv2v_reg;
  assign count_o[2] = count_o_2_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign N17 = reset_i | clear_i;
  assign { N9, N8, N6, N5 } = count_o + 1'b1;
  assign N10 = (N0)? 1'b1 : 
               (N7)? 1'b1 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = clear_i;
  assign N12 = (N1)? 1'b1 : 
               (N30)? 1'b0 : 1'b0;
  assign N1 = up_i;
  assign N11 = (N0)? up_i : 
               (N7)? N5 : 1'b0;
  assign N4 = N16;
  assign N13 = ~reset_i;
  assign N14 = ~clear_i;
  assign N15 = N13 & N14;
  assign N16 = up_i & N15;
  assign N2 = up_i | clear_i;
  assign N3 = ~N2;
  assign N7 = up_i & N14;
  assign N30 = ~up_i;

  always @(posedge clk_i) begin
    if(N17) begin
      count_o_3_sv2v_reg <= 1'b0;
      count_o_2_sv2v_reg <= 1'b0;
      count_o_1_sv2v_reg <= 1'b0;
    end else if(N12) begin
      count_o_3_sv2v_reg <= N9;
      count_o_2_sv2v_reg <= N8;
      count_o_1_sv2v_reg <= N6;
    end 
    if(reset_i) begin
      count_o_0_sv2v_reg <= 1'b0;
    end else if(N10) begin
      count_o_0_sv2v_reg <= N11;
    end 
  end


endmodule



module bsg_dff_en_0000008a
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [137:0] data_i;
  output [137:0] data_o;
  input clk_i;
  input en_i;
  wire [137:0] data_o;
  reg data_o_137_sv2v_reg,data_o_136_sv2v_reg,data_o_135_sv2v_reg,data_o_134_sv2v_reg,
  data_o_133_sv2v_reg,data_o_132_sv2v_reg,data_o_131_sv2v_reg,data_o_130_sv2v_reg,
  data_o_129_sv2v_reg,data_o_128_sv2v_reg,data_o_127_sv2v_reg,data_o_126_sv2v_reg,
  data_o_125_sv2v_reg,data_o_124_sv2v_reg,data_o_123_sv2v_reg,data_o_122_sv2v_reg,
  data_o_121_sv2v_reg,data_o_120_sv2v_reg,data_o_119_sv2v_reg,data_o_118_sv2v_reg,
  data_o_117_sv2v_reg,data_o_116_sv2v_reg,data_o_115_sv2v_reg,data_o_114_sv2v_reg,
  data_o_113_sv2v_reg,data_o_112_sv2v_reg,data_o_111_sv2v_reg,data_o_110_sv2v_reg,
  data_o_109_sv2v_reg,data_o_108_sv2v_reg,data_o_107_sv2v_reg,data_o_106_sv2v_reg,
  data_o_105_sv2v_reg,data_o_104_sv2v_reg,data_o_103_sv2v_reg,data_o_102_sv2v_reg,
  data_o_101_sv2v_reg,data_o_100_sv2v_reg,data_o_99_sv2v_reg,data_o_98_sv2v_reg,
  data_o_97_sv2v_reg,data_o_96_sv2v_reg,data_o_95_sv2v_reg,data_o_94_sv2v_reg,
  data_o_93_sv2v_reg,data_o_92_sv2v_reg,data_o_91_sv2v_reg,data_o_90_sv2v_reg,
  data_o_89_sv2v_reg,data_o_88_sv2v_reg,data_o_87_sv2v_reg,data_o_86_sv2v_reg,
  data_o_85_sv2v_reg,data_o_84_sv2v_reg,data_o_83_sv2v_reg,data_o_82_sv2v_reg,
  data_o_81_sv2v_reg,data_o_80_sv2v_reg,data_o_79_sv2v_reg,data_o_78_sv2v_reg,data_o_77_sv2v_reg,
  data_o_76_sv2v_reg,data_o_75_sv2v_reg,data_o_74_sv2v_reg,data_o_73_sv2v_reg,
  data_o_72_sv2v_reg,data_o_71_sv2v_reg,data_o_70_sv2v_reg,data_o_69_sv2v_reg,
  data_o_68_sv2v_reg,data_o_67_sv2v_reg,data_o_66_sv2v_reg,data_o_65_sv2v_reg,
  data_o_64_sv2v_reg,data_o_63_sv2v_reg,data_o_62_sv2v_reg,data_o_61_sv2v_reg,data_o_60_sv2v_reg,
  data_o_59_sv2v_reg,data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,
  data_o_55_sv2v_reg,data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,
  data_o_51_sv2v_reg,data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,
  data_o_47_sv2v_reg,data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,
  data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,
  data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,
  data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,
  data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,
  data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,
  data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,
  data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[137] = data_o_137_sv2v_reg;
  assign data_o[136] = data_o_136_sv2v_reg;
  assign data_o[135] = data_o_135_sv2v_reg;
  assign data_o[134] = data_o_134_sv2v_reg;
  assign data_o[133] = data_o_133_sv2v_reg;
  assign data_o[132] = data_o_132_sv2v_reg;
  assign data_o[131] = data_o_131_sv2v_reg;
  assign data_o[130] = data_o_130_sv2v_reg;
  assign data_o[129] = data_o_129_sv2v_reg;
  assign data_o[128] = data_o_128_sv2v_reg;
  assign data_o[127] = data_o_127_sv2v_reg;
  assign data_o[126] = data_o_126_sv2v_reg;
  assign data_o[125] = data_o_125_sv2v_reg;
  assign data_o[124] = data_o_124_sv2v_reg;
  assign data_o[123] = data_o_123_sv2v_reg;
  assign data_o[122] = data_o_122_sv2v_reg;
  assign data_o[121] = data_o_121_sv2v_reg;
  assign data_o[120] = data_o_120_sv2v_reg;
  assign data_o[119] = data_o_119_sv2v_reg;
  assign data_o[118] = data_o_118_sv2v_reg;
  assign data_o[117] = data_o_117_sv2v_reg;
  assign data_o[116] = data_o_116_sv2v_reg;
  assign data_o[115] = data_o_115_sv2v_reg;
  assign data_o[114] = data_o_114_sv2v_reg;
  assign data_o[113] = data_o_113_sv2v_reg;
  assign data_o[112] = data_o_112_sv2v_reg;
  assign data_o[111] = data_o_111_sv2v_reg;
  assign data_o[110] = data_o_110_sv2v_reg;
  assign data_o[109] = data_o_109_sv2v_reg;
  assign data_o[108] = data_o_108_sv2v_reg;
  assign data_o[107] = data_o_107_sv2v_reg;
  assign data_o[106] = data_o_106_sv2v_reg;
  assign data_o[105] = data_o_105_sv2v_reg;
  assign data_o[104] = data_o_104_sv2v_reg;
  assign data_o[103] = data_o_103_sv2v_reg;
  assign data_o[102] = data_o_102_sv2v_reg;
  assign data_o[101] = data_o_101_sv2v_reg;
  assign data_o[100] = data_o_100_sv2v_reg;
  assign data_o[99] = data_o_99_sv2v_reg;
  assign data_o[98] = data_o_98_sv2v_reg;
  assign data_o[97] = data_o_97_sv2v_reg;
  assign data_o[96] = data_o_96_sv2v_reg;
  assign data_o[95] = data_o_95_sv2v_reg;
  assign data_o[94] = data_o_94_sv2v_reg;
  assign data_o[93] = data_o_93_sv2v_reg;
  assign data_o[92] = data_o_92_sv2v_reg;
  assign data_o[91] = data_o_91_sv2v_reg;
  assign data_o[90] = data_o_90_sv2v_reg;
  assign data_o[89] = data_o_89_sv2v_reg;
  assign data_o[88] = data_o_88_sv2v_reg;
  assign data_o[87] = data_o_87_sv2v_reg;
  assign data_o[86] = data_o_86_sv2v_reg;
  assign data_o[85] = data_o_85_sv2v_reg;
  assign data_o[84] = data_o_84_sv2v_reg;
  assign data_o[83] = data_o_83_sv2v_reg;
  assign data_o[82] = data_o_82_sv2v_reg;
  assign data_o[81] = data_o_81_sv2v_reg;
  assign data_o[80] = data_o_80_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_137_sv2v_reg <= data_i[137];
      data_o_136_sv2v_reg <= data_i[136];
      data_o_135_sv2v_reg <= data_i[135];
      data_o_134_sv2v_reg <= data_i[134];
      data_o_133_sv2v_reg <= data_i[133];
      data_o_132_sv2v_reg <= data_i[132];
      data_o_131_sv2v_reg <= data_i[131];
      data_o_130_sv2v_reg <= data_i[130];
      data_o_129_sv2v_reg <= data_i[129];
      data_o_128_sv2v_reg <= data_i[128];
      data_o_127_sv2v_reg <= data_i[127];
      data_o_126_sv2v_reg <= data_i[126];
      data_o_125_sv2v_reg <= data_i[125];
      data_o_124_sv2v_reg <= data_i[124];
      data_o_123_sv2v_reg <= data_i[123];
      data_o_122_sv2v_reg <= data_i[122];
      data_o_121_sv2v_reg <= data_i[121];
      data_o_120_sv2v_reg <= data_i[120];
      data_o_119_sv2v_reg <= data_i[119];
      data_o_118_sv2v_reg <= data_i[118];
      data_o_117_sv2v_reg <= data_i[117];
      data_o_116_sv2v_reg <= data_i[116];
      data_o_115_sv2v_reg <= data_i[115];
      data_o_114_sv2v_reg <= data_i[114];
      data_o_113_sv2v_reg <= data_i[113];
      data_o_112_sv2v_reg <= data_i[112];
      data_o_111_sv2v_reg <= data_i[111];
      data_o_110_sv2v_reg <= data_i[110];
      data_o_109_sv2v_reg <= data_i[109];
      data_o_108_sv2v_reg <= data_i[108];
      data_o_107_sv2v_reg <= data_i[107];
      data_o_106_sv2v_reg <= data_i[106];
      data_o_105_sv2v_reg <= data_i[105];
      data_o_104_sv2v_reg <= data_i[104];
      data_o_103_sv2v_reg <= data_i[103];
      data_o_102_sv2v_reg <= data_i[102];
      data_o_101_sv2v_reg <= data_i[101];
      data_o_100_sv2v_reg <= data_i[100];
      data_o_99_sv2v_reg <= data_i[99];
      data_o_98_sv2v_reg <= data_i[98];
      data_o_97_sv2v_reg <= data_i[97];
      data_o_96_sv2v_reg <= data_i[96];
      data_o_95_sv2v_reg <= data_i[95];
      data_o_94_sv2v_reg <= data_i[94];
      data_o_93_sv2v_reg <= data_i[93];
      data_o_92_sv2v_reg <= data_i[92];
      data_o_91_sv2v_reg <= data_i[91];
      data_o_90_sv2v_reg <= data_i[90];
      data_o_89_sv2v_reg <= data_i[89];
      data_o_88_sv2v_reg <= data_i[88];
      data_o_87_sv2v_reg <= data_i[87];
      data_o_86_sv2v_reg <= data_i[86];
      data_o_85_sv2v_reg <= data_i[85];
      data_o_84_sv2v_reg <= data_i[84];
      data_o_83_sv2v_reg <= data_i[83];
      data_o_82_sv2v_reg <= data_i[82];
      data_o_81_sv2v_reg <= data_i[81];
      data_o_80_sv2v_reg <= data_i[80];
      data_o_79_sv2v_reg <= data_i[79];
      data_o_78_sv2v_reg <= data_i[78];
      data_o_77_sv2v_reg <= data_i[77];
      data_o_76_sv2v_reg <= data_i[76];
      data_o_75_sv2v_reg <= data_i[75];
      data_o_74_sv2v_reg <= data_i[74];
      data_o_73_sv2v_reg <= data_i[73];
      data_o_72_sv2v_reg <= data_i[72];
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_en_00000010
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [15:0] data_i;
  output [15:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [15:0] data_o;
  wire N0,N1,N2;
  reg data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,
  data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,
  data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bp_be_dcache_00
(
  clk_i,
  reset_i,
  cfg_bus_i,
  busy_o,
  ordered_o,
  dcache_pkt_i,
  v_i,
  ptag_i,
  ptag_v_i,
  ptag_uncached_i,
  ptag_dram_i,
  st_data_i,
  flush_i,
  v_o,
  data_o,
  rd_addr_o,
  tag_o,
  unsigned_o,
  int_o,
  float_o,
  ptw_o,
  ret_o,
  late_o,
  cache_req_o,
  cache_req_v_o,
  cache_req_yumi_i,
  cache_req_lock_i,
  cache_req_metadata_o,
  cache_req_metadata_v_o,
  cache_req_id_i,
  cache_req_critical_i,
  cache_req_last_i,
  cache_req_credits_full_i,
  cache_req_credits_empty_i,
  data_mem_pkt_v_i,
  data_mem_pkt_i,
  data_mem_pkt_yumi_o,
  data_mem_o,
  tag_mem_pkt_v_i,
  tag_mem_pkt_i,
  tag_mem_pkt_yumi_o,
  tag_mem_o,
  stat_mem_pkt_v_i,
  stat_mem_pkt_i,
  stat_mem_pkt_yumi_o,
  stat_mem_o
);

  input [60:0] cfg_bus_i;
  input [22:0] dcache_pkt_i;
  input [27:0] ptag_i;
  input [63:0] st_data_i;
  output [63:0] data_o;
  output [4:0] rd_addr_o;
  output [1:0] tag_o;
  output [116:0] cache_req_o;
  output [3:0] cache_req_metadata_o;
  input [0:0] cache_req_id_i;
  input [142:0] data_mem_pkt_i;
  output [511:0] data_mem_o;
  input [34:0] tag_mem_pkt_i;
  output [22:0] tag_mem_o;
  input [10:0] stat_mem_pkt_i;
  output [14:0] stat_mem_o;
  input clk_i;
  input reset_i;
  input v_i;
  input ptag_v_i;
  input ptag_uncached_i;
  input ptag_dram_i;
  input flush_i;
  input cache_req_yumi_i;
  input cache_req_lock_i;
  input cache_req_critical_i;
  input cache_req_last_i;
  input cache_req_credits_full_i;
  input cache_req_credits_empty_i;
  input data_mem_pkt_v_i;
  input tag_mem_pkt_v_i;
  input stat_mem_pkt_v_i;
  output busy_o;
  output ordered_o;
  output v_o;
  output unsigned_o;
  output int_o;
  output float_o;
  output ptw_o;
  output ret_o;
  output late_o;
  output cache_req_v_o;
  output cache_req_metadata_v_o;
  output data_mem_pkt_yumi_o;
  output tag_mem_pkt_yumi_o;
  output stat_mem_pkt_yumi_o;
  wire [63:0] data_o,data_mem_mask_li,st_data_tv_n,snoop_st_data,ld_data_way_picked,
  ld_data_dword_raw,ld_data_dword_merged,final_data_tv,atomic_reg_data,atomic_mem_data,
  atomic_alu_result,atomic_result,\wbuf_in_3_.slice_data ;
  wire [4:0] rd_addr_o;
  wire [1:0] tag_o,state_r,\wbuf_in_2_.addr_dec ,state_n;
  wire [116:0] cache_req_o;
  wire [3:0] cache_req_metadata_o,\wbuf_in_1_.addr_dec ,\l1_lrsc.lrsc_lock_cnt ;
  wire [511:0] data_mem_o,data_mem_data_li,data_mem_data_lo,ld_data_tv_n,ld_data_tv_r;
  wire [22:0] tag_mem_o;
  wire [14:0] stat_mem_o,stat_mem_data_li,stat_mem_mask_li;
  wire busy_o,ordered_o,v_o,unsigned_o,int_o,float_o,ptw_o,ret_o,late_o,cache_req_v_o,
  cache_req_metadata_v_o,data_mem_pkt_yumi_o,tag_mem_pkt_yumi_o,
  stat_mem_pkt_yumi_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,blocking_hazard,nonblocking_hazard,fill_hazard,
  flush_tv,data_mem_write_hazard,flush_tl,critical_recv,complete_recv,tag_mem_v_li,
  tag_mem_w_li,safe_tl_we,tl_we,v_tl_r,N89,\tag_comp_tl_0_.tag_match_tl ,N90,N91,N92,
  N93,N94,N95,N96,N97,N98,N99,\tag_comp_tl_1_.tag_match_tl ,N100,N101,N102,N103,
  N104,N105,N106,N107,N108,N109,\tag_comp_tl_2_.tag_match_tl ,N110,N111,N112,N113,
  N114,N115,N116,N117,N118,N119,\tag_comp_tl_3_.tag_match_tl ,N120,N121,N122,N123,
  N124,N125,N126,N127,N128,N129,\tag_comp_tl_4_.tag_match_tl ,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,\tag_comp_tl_5_.tag_match_tl ,N140,N141,N142,N143,
  N144,N145,N146,N147,N148,N149,\tag_comp_tl_6_.tag_match_tl ,N150,N151,N152,N153,
  N154,N155,N156,N157,N158,N159,\tag_comp_tl_7_.tag_match_tl ,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,uncached_tl,safe_tv_we,tv_we,_2_net_,v_tv_r,uncached_tv_n,
  snoop_paddr_5,snoop_paddr_4,snoop_paddr_3,snoop_paddr_2,snoop_paddr_1,
  snoop_paddr_0,snoop_uncached,decode_tv_r_load_op_,decode_tv_r_store_op_,
  decode_tv_r_signed_op_,decode_tv_r_cache_op_,decode_tv_r_block_op_,decode_tv_r_double_op_,
  decode_tv_r_word_op_,decode_tv_r_half_op_,decode_tv_r_byte_op_,decode_tv_r_uncached_op_,
  decode_tv_r_lr_op_,decode_tv_r_sc_op_,decode_tv_r_amo_op_,decode_tv_r_clean_op_,
  decode_tv_r_inval_op_,decode_tv_r_bclean_op_,decode_tv_r_binval_op_,
  decode_tv_r_bzero_op_,decode_tv_r_amo_subop__3_,decode_tv_r_amo_subop__2_,
  decode_tv_r_amo_subop__1_,decode_tv_r_amo_subop__0_,uncached_tv_r,store_hit_tv,sc_fail_tv,
  nonblocking_req,store_miss_tv,load_miss_tv,blocking_miss_tv,nonblocking_miss_tv,
  engine_miss_tv,any_miss_tv,sc_success_tv,N169,N170,N171,N172,N173,stat_mem_v_li,
  stat_mem_w_li,wbuf_v_li,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
  N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,
  N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,
  N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,
  N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,
  N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,
  N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,
  N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,
  N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,
  N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,
  N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,
  N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,
  N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,
  N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,
  N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,
  N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,
  N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,
  N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,
  N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,
  N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,
  N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,
  N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,
  N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,
  N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,
  N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,
  N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,
  N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,
  N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,
  N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,
  N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,
  N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,
  N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,
  N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,
  N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,
  N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,
  N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,
  N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,
  N763,N764,N765,N766,N767,N768,wbuf_entry_in_bank_sel__7_,
  wbuf_entry_in_bank_sel__6_,wbuf_entry_in_bank_sel__5_,wbuf_entry_in_bank_sel__4_,
  wbuf_entry_in_bank_sel__3_,wbuf_entry_in_bank_sel__2_,wbuf_entry_in_bank_sel__1_,
  wbuf_entry_in_bank_sel__0_,wbuf_entry_in_mask__7_,wbuf_entry_in_mask__6_,wbuf_entry_in_mask__5_,
  wbuf_entry_in_mask__4_,wbuf_entry_in_mask__3_,wbuf_entry_in_mask__2_,
  wbuf_entry_in_mask__1_,wbuf_entry_in_mask__0_,wbuf_entry_in_data__63_,wbuf_entry_in_data__62_,
  wbuf_entry_in_data__61_,wbuf_entry_in_data__60_,wbuf_entry_in_data__59_,
  wbuf_entry_in_data__58_,wbuf_entry_in_data__57_,wbuf_entry_in_data__56_,
  wbuf_entry_in_data__55_,wbuf_entry_in_data__54_,wbuf_entry_in_data__53_,wbuf_entry_in_data__52_,
  wbuf_entry_in_data__51_,wbuf_entry_in_data__50_,wbuf_entry_in_data__49_,
  wbuf_entry_in_data__48_,wbuf_entry_in_data__47_,wbuf_entry_in_data__46_,
  wbuf_entry_in_data__45_,wbuf_entry_in_data__44_,wbuf_entry_in_data__43_,wbuf_entry_in_data__42_,
  wbuf_entry_in_data__41_,wbuf_entry_in_data__40_,wbuf_entry_in_data__39_,
  wbuf_entry_in_data__38_,wbuf_entry_in_data__37_,wbuf_entry_in_data__36_,
  wbuf_entry_in_data__35_,wbuf_entry_in_data__34_,wbuf_entry_in_data__33_,wbuf_entry_in_data__32_,
  wbuf_entry_in_data__31_,wbuf_entry_in_data__30_,wbuf_entry_in_data__29_,
  wbuf_entry_in_data__28_,wbuf_entry_in_data__27_,wbuf_entry_in_data__26_,
  wbuf_entry_in_data__25_,wbuf_entry_in_data__24_,wbuf_entry_in_data__23_,wbuf_entry_in_data__22_,
  wbuf_entry_in_data__21_,wbuf_entry_in_data__20_,wbuf_entry_in_data__19_,
  wbuf_entry_in_data__18_,wbuf_entry_in_data__17_,wbuf_entry_in_data__16_,
  wbuf_entry_in_data__15_,wbuf_entry_in_data__14_,wbuf_entry_in_data__13_,wbuf_entry_in_data__12_,
  wbuf_entry_in_data__11_,wbuf_entry_in_data__10_,wbuf_entry_in_data__9_,
  wbuf_entry_in_data__8_,wbuf_entry_in_data__7_,wbuf_entry_in_data__6_,
  wbuf_entry_in_data__5_,wbuf_entry_in_data__4_,wbuf_entry_in_data__3_,wbuf_entry_in_data__2_,
  wbuf_entry_in_data__1_,wbuf_entry_in_data__0_,wbuf_v_lo,wbuf_force_lo,wbuf_yumi_li,
  wbuf_entry_out_snoop_,wbuf_entry_out_bank_sel__7_,wbuf_entry_out_bank_sel__6_,
  wbuf_entry_out_bank_sel__5_,wbuf_entry_out_bank_sel__4_,wbuf_entry_out_bank_sel__3_,
  wbuf_entry_out_bank_sel__2_,wbuf_entry_out_bank_sel__1_,wbuf_entry_out_bank_sel__0_,
  wbuf_entry_out_data__63_,wbuf_entry_out_data__62_,wbuf_entry_out_data__61_,
  wbuf_entry_out_data__60_,wbuf_entry_out_data__59_,wbuf_entry_out_data__58_,
  wbuf_entry_out_data__57_,wbuf_entry_out_data__56_,wbuf_entry_out_data__55_,
  wbuf_entry_out_data__54_,wbuf_entry_out_data__53_,wbuf_entry_out_data__52_,
  wbuf_entry_out_data__51_,wbuf_entry_out_data__50_,wbuf_entry_out_data__49_,wbuf_entry_out_data__48_,
  wbuf_entry_out_data__47_,wbuf_entry_out_data__46_,wbuf_entry_out_data__45_,
  wbuf_entry_out_data__44_,wbuf_entry_out_data__43_,wbuf_entry_out_data__42_,
  wbuf_entry_out_data__41_,wbuf_entry_out_data__40_,wbuf_entry_out_data__39_,
  wbuf_entry_out_data__38_,wbuf_entry_out_data__37_,wbuf_entry_out_data__36_,
  wbuf_entry_out_data__35_,wbuf_entry_out_data__34_,wbuf_entry_out_data__33_,wbuf_entry_out_data__32_,
  wbuf_entry_out_data__31_,wbuf_entry_out_data__30_,wbuf_entry_out_data__29_,
  wbuf_entry_out_data__28_,wbuf_entry_out_data__27_,wbuf_entry_out_data__26_,
  wbuf_entry_out_data__25_,wbuf_entry_out_data__24_,wbuf_entry_out_data__23_,
  wbuf_entry_out_data__22_,wbuf_entry_out_data__21_,wbuf_entry_out_data__20_,
  wbuf_entry_out_data__19_,wbuf_entry_out_data__18_,wbuf_entry_out_data__17_,wbuf_entry_out_data__16_,
  wbuf_entry_out_data__15_,wbuf_entry_out_data__14_,wbuf_entry_out_data__13_,
  wbuf_entry_out_data__12_,wbuf_entry_out_data__11_,wbuf_entry_out_data__10_,
  wbuf_entry_out_data__9_,wbuf_entry_out_data__8_,wbuf_entry_out_data__7_,
  wbuf_entry_out_data__6_,wbuf_entry_out_data__5_,wbuf_entry_out_data__4_,wbuf_entry_out_data__3_,
  wbuf_entry_out_data__2_,wbuf_entry_out_data__1_,wbuf_entry_out_data__0_,
  wbuf_entry_out_caddr__31_,wbuf_entry_out_caddr__30_,wbuf_entry_out_caddr__29_,
  wbuf_entry_out_caddr__28_,wbuf_entry_out_caddr__27_,wbuf_entry_out_caddr__26_,
  wbuf_entry_out_caddr__25_,wbuf_entry_out_caddr__24_,wbuf_entry_out_caddr__23_,
  wbuf_entry_out_caddr__22_,wbuf_entry_out_caddr__21_,wbuf_entry_out_caddr__20_,
  wbuf_entry_out_caddr__19_,wbuf_entry_out_caddr__18_,wbuf_entry_out_caddr__17_,
  wbuf_entry_out_caddr__16_,wbuf_entry_out_caddr__15_,wbuf_entry_out_caddr__14_,
  wbuf_entry_out_caddr__13_,wbuf_entry_out_caddr__12_,wbuf_entry_out_caddr__11_,
  wbuf_entry_out_caddr__10_,wbuf_entry_out_caddr__9_,wbuf_entry_out_caddr__8_,wbuf_entry_out_caddr__7_,
  wbuf_entry_out_caddr__6_,wbuf_entry_out_caddr__5_,wbuf_entry_out_caddr__4_,
  wbuf_entry_out_caddr__3_,wbuf_entry_out_caddr__2_,wbuf_entry_out_caddr__1_,
  wbuf_entry_out_caddr__0_,wbuf_snoop_match_lo,load_req,store_req,uncached_amo_req,
  uncached_load_req,uncached_store_req,bclean_req,inval_req,clean_req,flush_req,blocking_sent,
  N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,
  N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,
  N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,
  N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,
  N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,
  N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,
  N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,
  metadata_hit_r,_14_net__7_,_14_net__6_,_14_net__5_,_14_net__4_,_14_net__3_,
  _14_net__2_,_14_net__1_,_14_net__0_,metadata_invalid_exist,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,tag_mem_fast_read,
  tag_mem_slow_read,tag_mem_slow_write,tag_mem_fast_write,N897,N898,N899,N900,N901,N902,
  N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,N918,
  N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,N934,
  N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,N950,
  N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,N966,
  N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,N982,
  N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,N998,
  N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012,
  N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,N1025,
  N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038,
  N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,
  N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,N1065,
  N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,
  N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091,N1092,
  N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,N1105,
  N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118,
  N1119,N1120,N1121,N1122,N1123,stat_mem_fast_read,stat_mem_fast_write,
  stat_mem_slow_write,stat_mem_slow_read,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  \tdm.dirty_mask_v_li ,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,
  N1143,\l1_lrsc.set_reservation ,\l1_lrsc.load_reserved_v_r ,N1144,N1145,
  \l1_lrsc.clear_reservation ,N1146,N1147,\l1_lrsc.load_reservation_match_tv ,
  \l1_lrsc.lrsc_lock_up ,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,
  N1159,N1160,\hum.fill_v ,\hum.fill_recv ,N1161,N1162,N1163,N1164,N1165,N1166,N1167,
  N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,_25_net_,N1178,
  N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,
  N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,
  N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,
  N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,
  N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,
  N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,
  N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,
  N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,
  N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,
  N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,
  N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,
  N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,
  N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,
  N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,
  N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,
  N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,
  N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,
  N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,
  N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,
  N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,
  N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,
  N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,
  N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,
  N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,
  N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,
  N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,
  N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
  N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,
  N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,
  N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,
  N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,
  N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,
  N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,
  N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,
  N1633,N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,
  N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,
  N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,
  N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,
  N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,
  N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,
  N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,
  N1726,N1727,N1728,N1729,N1730;
  wire [32:0] decode_lo,decode_tl_r,decode_tv_n,snoop_decode;
  wire [5:0] tag_mem_addr_li,stat_mem_addr_li,\l1_lrsc.load_reserved_index_r ,
  \hum.fill_index ;
  wire [183:0] tag_mem_data_li,tag_mem_mask_li,tag_mem_data_lo;
  wire [7:0] data_mem_v_li,data_mem_w_li,load_hit_tl,store_hit_tl,bank_sel_one_hot_tl,
  way_v_tv_n,store_hit_tv_n,load_hit_tv_n,bank_sel_one_hot_tv_n,snoop_bank_sel_one_hot,
  way_v_tv_r,store_hit_v_tv_r,load_hit_v_tv_r,bank_sel_one_hot_tv_r,
  ld_data_way_select_tv,\wbuf_in_0_.addr_dec ,metadata_way_v_r,tag_mem_way_one_hot,
  data_mem_pkt_fill_mask_expanded,data_mem_write_bank_mask,wbuf_data_mem_mask,
  data_mem_force_write,data_mem_slow_write,data_mem_slow_read,data_mem_fast_write,dirty_mask_lo,
  \hum.fill_bank_mask_r ,\hum.fill_bank_mask_n ,\hum.fill_hit_n ,\hum.fill_hit_r ,
  pseudo_hit;
  wire [71:0] data_mem_addr_li;
  wire [11:0] paddr_tl;
  wire [39:0] paddr_tv_n;
  wire [39:12] snoop_paddr;
  wire [2:0] store_hit_way_tv,load_hit_way_tv,lru_encode,metadata_hit_index_r,
  metadata_invalid_way,lru_way_li,tag_mem_pkt_way_r,\data_mem_lines_0_.data_mem_pkt_offset ,
  \data_mem_lines_1_.data_mem_pkt_offset ,\data_mem_lines_2_.data_mem_pkt_offset ,
  \data_mem_lines_3_.data_mem_pkt_offset ,\data_mem_lines_4_.data_mem_pkt_offset ,
  \data_mem_lines_5_.data_mem_pkt_offset ,\data_mem_lines_6_.data_mem_pkt_offset ,
  \data_mem_lines_7_.data_mem_pkt_offset ,data_mem_pkt_way_r,lru_decode_way_li,
  \tdm.dirty_mask_way_li ,stat_mem_pkt_way_r;
  wire [63:32] amo32_reg_in,amo64_reg_in;
  wire [31:0] wbuf_data_mem_mask_in,\wbuf_in_2_.slice_data ;
  wire [0:0] \wbuf_in_3_.addr_dec ,data_mem_fast_read;
  wire [127:0] data_mem_pkt_fill_data_li;
  wire [6:0] lru_decode_data_lo,lru_decode_mask_lo;
  wire [19:0] \l1_lrsc.load_reserved_tag_r ;
  reg state_r_1_sv2v_reg,state_r_0_sv2v_reg;
  assign state_r[1] = state_r_1_sv2v_reg;
  assign state_r[0] = state_r_0_sv2v_reg;
  assign cache_req_o[116] = 1'b0;

  bp_be_dcache_decoder_00_00000ffe
  pkt_decoder
  (
    .pkt_i(dcache_pkt_i),
    .decode_o(decode_lo)
  );


  bsg_mem_1rw_sync_mask_write_bit_000000b8_00000040_1
  tag_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(tag_mem_data_li),
    .addr_i(tag_mem_addr_li),
    .v_i(tag_mem_v_li),
    .w_mask_i(tag_mem_mask_li),
    .w_i(tag_mem_w_li),
    .data_o(tag_mem_data_lo)
  );


  bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
  \d_0_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li[0]),
    .w_i(data_mem_w_li[0]),
    .addr_i(data_mem_addr_li[8:0]),
    .data_i(data_mem_data_li[63:0]),
    .write_mask_i(data_mem_mask_li[7:0]),
    .data_o(data_mem_data_lo[63:0])
  );


  bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
  \d_1_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li[1]),
    .w_i(data_mem_w_li[1]),
    .addr_i(data_mem_addr_li[17:9]),
    .data_i(data_mem_data_li[127:64]),
    .write_mask_i(data_mem_mask_li[15:8]),
    .data_o(data_mem_data_lo[127:64])
  );


  bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
  \d_2_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li[2]),
    .w_i(data_mem_w_li[2]),
    .addr_i(data_mem_addr_li[26:18]),
    .data_i(data_mem_data_li[191:128]),
    .write_mask_i(data_mem_mask_li[23:16]),
    .data_o(data_mem_data_lo[191:128])
  );


  bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
  \d_3_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li[3]),
    .w_i(data_mem_w_li[3]),
    .addr_i(data_mem_addr_li[35:27]),
    .data_i(data_mem_data_li[255:192]),
    .write_mask_i(data_mem_mask_li[31:24]),
    .data_o(data_mem_data_lo[255:192])
  );


  bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
  \d_4_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li[4]),
    .w_i(data_mem_w_li[4]),
    .addr_i(data_mem_addr_li[44:36]),
    .data_i(data_mem_data_li[319:256]),
    .write_mask_i(data_mem_mask_li[39:32]),
    .data_o(data_mem_data_lo[319:256])
  );


  bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
  \d_5_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li[5]),
    .w_i(data_mem_w_li[5]),
    .addr_i(data_mem_addr_li[53:45]),
    .data_i(data_mem_data_li[383:320]),
    .write_mask_i(data_mem_mask_li[47:40]),
    .data_o(data_mem_data_lo[383:320])
  );


  bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
  \d_6_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li[6]),
    .w_i(data_mem_w_li[6]),
    .addr_i(data_mem_addr_li[62:54]),
    .data_i(data_mem_data_li[447:384]),
    .write_mask_i(data_mem_mask_li[55:48]),
    .data_o(data_mem_data_lo[447:384])
  );


  bsg_mem_1rw_sync_mask_write_byte_00000200_00000040_1
  \d_7_.data_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li[7]),
    .w_i(data_mem_w_li[7]),
    .addr_i(data_mem_addr_li[71:63]),
    .data_i(data_mem_data_li[511:448]),
    .write_mask_i(data_mem_mask_li[63:56]),
    .data_o(data_mem_data_lo[511:448])
  );


  bsg_dff_reset_width_p1
  v_tl_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(tl_we),
    .data_o(v_tl_r)
  );


  bsg_dff_width_p45
  tl_stage_reg
  (
    .clk_i(clk_i),
    .data_i({ dcache_pkt_i[11:0], decode_lo }),
    .data_o({ paddr_tl, decode_tl_r })
  );

  assign N89 = ptag_i[19:0] == tag_mem_data_lo[19:0];
  assign N90 = ~tag_mem_data_lo[22];
  assign N91 = ~tag_mem_data_lo[21];
  assign N92 = N91 | N90;
  assign N93 = tag_mem_data_lo[20] | N92;
  assign N94 = ~N93;
  assign N95 = N91 | tag_mem_data_lo[22];
  assign N96 = tag_mem_data_lo[20] | N95;
  assign N97 = ~N96;
  assign N98 = N94 | N97;
  assign N99 = ptag_i[19:0] == tag_mem_data_lo[42:23];
  assign N100 = ~tag_mem_data_lo[45];
  assign N101 = ~tag_mem_data_lo[44];
  assign N102 = N101 | N100;
  assign N103 = tag_mem_data_lo[43] | N102;
  assign N104 = ~N103;
  assign N105 = N101 | tag_mem_data_lo[45];
  assign N106 = tag_mem_data_lo[43] | N105;
  assign N107 = ~N106;
  assign N108 = N104 | N107;
  assign N109 = ptag_i[19:0] == tag_mem_data_lo[65:46];
  assign N110 = ~tag_mem_data_lo[68];
  assign N111 = ~tag_mem_data_lo[67];
  assign N112 = N111 | N110;
  assign N113 = tag_mem_data_lo[66] | N112;
  assign N114 = ~N113;
  assign N115 = N111 | tag_mem_data_lo[68];
  assign N116 = tag_mem_data_lo[66] | N115;
  assign N117 = ~N116;
  assign N118 = N114 | N117;
  assign N119 = ptag_i[19:0] == tag_mem_data_lo[88:69];
  assign N120 = ~tag_mem_data_lo[91];
  assign N121 = ~tag_mem_data_lo[90];
  assign N122 = N121 | N120;
  assign N123 = tag_mem_data_lo[89] | N122;
  assign N124 = ~N123;
  assign N125 = N121 | tag_mem_data_lo[91];
  assign N126 = tag_mem_data_lo[89] | N125;
  assign N127 = ~N126;
  assign N128 = N124 | N127;
  assign N129 = ptag_i[19:0] == tag_mem_data_lo[111:92];
  assign N130 = ~tag_mem_data_lo[114];
  assign N131 = ~tag_mem_data_lo[113];
  assign N132 = N131 | N130;
  assign N133 = tag_mem_data_lo[112] | N132;
  assign N134 = ~N133;
  assign N135 = N131 | tag_mem_data_lo[114];
  assign N136 = tag_mem_data_lo[112] | N135;
  assign N137 = ~N136;
  assign N138 = N134 | N137;
  assign N139 = ptag_i[19:0] == tag_mem_data_lo[134:115];
  assign N140 = ~tag_mem_data_lo[137];
  assign N141 = ~tag_mem_data_lo[136];
  assign N142 = N141 | N140;
  assign N143 = tag_mem_data_lo[135] | N142;
  assign N144 = ~N143;
  assign N145 = N141 | tag_mem_data_lo[137];
  assign N146 = tag_mem_data_lo[135] | N145;
  assign N147 = ~N146;
  assign N148 = N144 | N147;
  assign N149 = ptag_i[19:0] == tag_mem_data_lo[157:138];
  assign N150 = ~tag_mem_data_lo[160];
  assign N151 = ~tag_mem_data_lo[159];
  assign N152 = N151 | N150;
  assign N153 = tag_mem_data_lo[158] | N152;
  assign N154 = ~N153;
  assign N155 = N151 | tag_mem_data_lo[160];
  assign N156 = tag_mem_data_lo[158] | N155;
  assign N157 = ~N156;
  assign N158 = N154 | N157;
  assign N159 = ptag_i[19:0] == tag_mem_data_lo[180:161];
  assign N160 = ~tag_mem_data_lo[183];
  assign N161 = ~tag_mem_data_lo[182];
  assign N162 = N161 | N160;
  assign N163 = tag_mem_data_lo[181] | N162;
  assign N164 = ~N163;
  assign N165 = N161 | tag_mem_data_lo[183];
  assign N166 = tag_mem_data_lo[181] | N165;
  assign N167 = ~N166;
  assign N168 = N164 | N167;

  bsg_decode_00000008
  offset_decode
  (
    .i(paddr_tl[5:3]),
    .o(bank_sel_one_hot_tl)
  );


  bsg_dff_reset_width_p1
  v_tv_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(_2_net_),
    .data_o(v_tv_r)
  );


  bsg_mux_000002aa_2
  tv_snoop_mux
  (
    .data_i({ pseudo_hit, pseudo_hit, pseudo_hit, data_mem_data_li, snoop_st_data, snoop_paddr, \hum.fill_index , snoop_paddr_5, snoop_paddr_4, snoop_paddr_3, snoop_paddr_2, snoop_paddr_1, snoop_paddr_0, snoop_bank_sel_one_hot, snoop_uncached, snoop_decode, N1196, N1198, N1200, N1202, N1204, N1206, N1208, N1210, store_hit_tl, load_hit_tl, data_mem_data_lo, st_data_i, ptag_i, paddr_tl, bank_sel_one_hot_tl, uncached_tl, decode_tl_r }),
    .sel_i(critical_recv),
    .data_o({ way_v_tv_n, store_hit_tv_n, load_hit_tv_n, ld_data_tv_n, st_data_tv_n, paddr_tv_n, bank_sel_one_hot_tv_n, uncached_tv_n, decode_tv_n })
  );


  bsg_dff_000002ab
  tv_stage_reg
  (
    .clk_i(clk_i),
    .data_i({ critical_recv, way_v_tv_n, store_hit_tv_n, load_hit_tv_n, paddr_tv_n, ld_data_tv_n, st_data_tv_n, bank_sel_one_hot_tv_n, uncached_tv_n, decode_tv_n }),
    .data_o({ late_o, way_v_tv_r, store_hit_v_tv_r, load_hit_v_tv_r, cache_req_o[47:8], ld_data_tv_r, amo64_reg_in, amo32_reg_in, bank_sel_one_hot_tv_r, uncached_tv_r, tag_o, decode_tv_r_load_op_, ret_o, decode_tv_r_store_op_, decode_tv_r_signed_op_, float_o, int_o, ptw_o, decode_tv_r_cache_op_, decode_tv_r_block_op_, decode_tv_r_double_op_, decode_tv_r_word_op_, decode_tv_r_half_op_, decode_tv_r_byte_op_, decode_tv_r_uncached_op_, decode_tv_r_lr_op_, decode_tv_r_sc_op_, decode_tv_r_amo_op_, decode_tv_r_clean_op_, decode_tv_r_inval_op_, decode_tv_r_bclean_op_, decode_tv_r_binval_op_, decode_tv_r_bzero_op_, decode_tv_r_amo_subop__3_, decode_tv_r_amo_subop__2_, decode_tv_r_amo_subop__1_, decode_tv_r_amo_subop__0_, rd_addr_o })
  );


  bsg_encode_one_hot_00000008_1
  store_hit_index_encoder
  (
    .i(store_hit_v_tv_r),
    .addr_o(store_hit_way_tv),
    .v_o(store_hit_tv)
  );


  bsg_encode_one_hot_00000008_1
  load_hit_index_encoder
  (
    .i(load_hit_v_tv_r),
    .addr_o(load_hit_way_tv),
    .v_o(cache_req_o[115])
  );


  bsg_adder_one_hot_00000008
  select_adder
  (
    .a_i(load_hit_v_tv_r),
    .b_i(bank_sel_one_hot_tv_r),
    .o(ld_data_way_select_tv)
  );


  bsg_mux_one_hot_00000040_00000008
  ld_data_set_select_mux
  (
    .data_i(ld_data_tv_r),
    .sel_one_hot_i(ld_data_way_select_tv),
    .data_o(ld_data_way_picked)
  );


  bsg_mux_00000040_00000001
  dword_mux
  (
    .data_i(ld_data_way_picked),
    .sel_i(cache_req_o[11]),
    .data_o(ld_data_dword_raw)
  );

  assign final_data_tv = ld_data_dword_merged >> { cache_req_o[10:8], 1'b0, 1'b0, 1'b0 };

  bsg_mem_1rw_sync_mask_write_bit_0000000f_00000040_1
  stat_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(stat_mem_data_li),
    .addr_i(stat_mem_addr_li),
    .v_i(stat_mem_v_li),
    .w_mask_i(stat_mem_mask_li),
    .w_i(stat_mem_w_li),
    .data_o(stat_mem_o)
  );


  bsg_lru_pseudo_tree_encode_00000008
  lru_encoder
  (
    .lru_i(stat_mem_o[14:8]),
    .way_id_o(lru_encode)
  );

  assign N438 = $signed(atomic_reg_data) < $signed(atomic_mem_data);
  assign N504 = $signed(atomic_reg_data) > $signed(atomic_mem_data);
  assign N570 = atomic_reg_data < atomic_mem_data;
  assign N636 = atomic_reg_data > atomic_mem_data;

  bsg_decode_00000008
  \wbuf_in_0_.decode 
  (
    .i(cache_req_o[10:8]),
    .o(\wbuf_in_0_.addr_dec )
  );


  bsg_expand_bitmask_in_width_p8_expand_p1
  \wbuf_in_0_.expand 
  (
    .i(\wbuf_in_0_.addr_dec ),
    .o(wbuf_data_mem_mask_in[7:0])
  );


  bsg_decode_num_out_p4
  \wbuf_in_1_.decode 
  (
    .i(cache_req_o[10:9]),
    .o(\wbuf_in_1_.addr_dec )
  );


  bsg_expand_bitmask_in_width_p4_expand_p2
  \wbuf_in_1_.expand 
  (
    .i(\wbuf_in_1_.addr_dec ),
    .o(wbuf_data_mem_mask_in[15:8])
  );


  bsg_decode_num_out_p2
  \wbuf_in_2_.decode 
  (
    .i(cache_req_o[10]),
    .o(\wbuf_in_2_.addr_dec )
  );


  bsg_expand_bitmask_in_width_p2_expand_p4
  \wbuf_in_2_.expand 
  (
    .i(\wbuf_in_2_.addr_dec ),
    .o(wbuf_data_mem_mask_in[23:16])
  );


  bsg_decode_num_out_p1
  \wbuf_in_3_.decode 
  (
    .i(cache_req_o[11]),
    .o(\wbuf_in_3_.addr_dec [0])
  );


  bsg_expand_bitmask_in_width_p1_expand_p8
  \wbuf_in_3_.expand 
  (
    .i(\wbuf_in_3_.addr_dec [0]),
    .o(wbuf_data_mem_mask_in[31:24])
  );


  bsg_mux_one_hot_width_p64_els_p4
  wbuf_data_in_mux
  (
    .data_i({ \wbuf_in_3_.slice_data , \wbuf_in_2_.slice_data , \wbuf_in_2_.slice_data , amo32_reg_in[47:32], amo32_reg_in[47:32], amo32_reg_in[47:32], amo32_reg_in[47:32], amo32_reg_in[39:32], amo32_reg_in[39:32], amo32_reg_in[39:32], amo32_reg_in[39:32], amo32_reg_in[39:32], amo32_reg_in[39:32], amo32_reg_in[39:32], amo32_reg_in[39:32] }),
    .sel_one_hot_i({ decode_tv_r_double_op_, decode_tv_r_word_op_, decode_tv_r_half_op_, decode_tv_r_byte_op_ }),
    .data_o({ wbuf_entry_in_data__63_, wbuf_entry_in_data__62_, wbuf_entry_in_data__61_, wbuf_entry_in_data__60_, wbuf_entry_in_data__59_, wbuf_entry_in_data__58_, wbuf_entry_in_data__57_, wbuf_entry_in_data__56_, wbuf_entry_in_data__55_, wbuf_entry_in_data__54_, wbuf_entry_in_data__53_, wbuf_entry_in_data__52_, wbuf_entry_in_data__51_, wbuf_entry_in_data__50_, wbuf_entry_in_data__49_, wbuf_entry_in_data__48_, wbuf_entry_in_data__47_, wbuf_entry_in_data__46_, wbuf_entry_in_data__45_, wbuf_entry_in_data__44_, wbuf_entry_in_data__43_, wbuf_entry_in_data__42_, wbuf_entry_in_data__41_, wbuf_entry_in_data__40_, wbuf_entry_in_data__39_, wbuf_entry_in_data__38_, wbuf_entry_in_data__37_, wbuf_entry_in_data__36_, wbuf_entry_in_data__35_, wbuf_entry_in_data__34_, wbuf_entry_in_data__33_, wbuf_entry_in_data__32_, wbuf_entry_in_data__31_, wbuf_entry_in_data__30_, wbuf_entry_in_data__29_, wbuf_entry_in_data__28_, wbuf_entry_in_data__27_, wbuf_entry_in_data__26_, wbuf_entry_in_data__25_, wbuf_entry_in_data__24_, wbuf_entry_in_data__23_, wbuf_entry_in_data__22_, wbuf_entry_in_data__21_, wbuf_entry_in_data__20_, wbuf_entry_in_data__19_, wbuf_entry_in_data__18_, wbuf_entry_in_data__17_, wbuf_entry_in_data__16_, wbuf_entry_in_data__15_, wbuf_entry_in_data__14_, wbuf_entry_in_data__13_, wbuf_entry_in_data__12_, wbuf_entry_in_data__11_, wbuf_entry_in_data__10_, wbuf_entry_in_data__9_, wbuf_entry_in_data__8_, wbuf_entry_in_data__7_, wbuf_entry_in_data__6_, wbuf_entry_in_data__5_, wbuf_entry_in_data__4_, wbuf_entry_in_data__3_, wbuf_entry_in_data__2_, wbuf_entry_in_data__1_, wbuf_entry_in_data__0_ })
  );


  bsg_mux_one_hot_00000008_4
  wbuf_data_mem_mask_in_mux
  (
    .data_i(wbuf_data_mem_mask_in),
    .sel_one_hot_i({ decode_tv_r_double_op_, decode_tv_r_word_op_, decode_tv_r_half_op_, decode_tv_r_byte_op_ }),
    .data_o({ wbuf_entry_in_mask__7_, wbuf_entry_in_mask__6_, wbuf_entry_in_mask__5_, wbuf_entry_in_mask__4_, wbuf_entry_in_mask__3_, wbuf_entry_in_mask__2_, wbuf_entry_in_mask__1_, wbuf_entry_in_mask__0_ })
  );


  bp_be_dcache_wbuf_00_00000040_00000008_00000200_00000080_00000014
  wbuf
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .wbuf_entry_i({ late_o, wbuf_entry_in_bank_sel__7_, wbuf_entry_in_bank_sel__6_, wbuf_entry_in_bank_sel__5_, wbuf_entry_in_bank_sel__4_, wbuf_entry_in_bank_sel__3_, wbuf_entry_in_bank_sel__2_, wbuf_entry_in_bank_sel__1_, wbuf_entry_in_bank_sel__0_, wbuf_entry_in_mask__7_, wbuf_entry_in_mask__6_, wbuf_entry_in_mask__5_, wbuf_entry_in_mask__4_, wbuf_entry_in_mask__3_, wbuf_entry_in_mask__2_, wbuf_entry_in_mask__1_, wbuf_entry_in_mask__0_, wbuf_entry_in_data__63_, wbuf_entry_in_data__62_, wbuf_entry_in_data__61_, wbuf_entry_in_data__60_, wbuf_entry_in_data__59_, wbuf_entry_in_data__58_, wbuf_entry_in_data__57_, wbuf_entry_in_data__56_, wbuf_entry_in_data__55_, wbuf_entry_in_data__54_, wbuf_entry_in_data__53_, wbuf_entry_in_data__52_, wbuf_entry_in_data__51_, wbuf_entry_in_data__50_, wbuf_entry_in_data__49_, wbuf_entry_in_data__48_, wbuf_entry_in_data__47_, wbuf_entry_in_data__46_, wbuf_entry_in_data__45_, wbuf_entry_in_data__44_, wbuf_entry_in_data__43_, wbuf_entry_in_data__42_, wbuf_entry_in_data__41_, wbuf_entry_in_data__40_, wbuf_entry_in_data__39_, wbuf_entry_in_data__38_, wbuf_entry_in_data__37_, wbuf_entry_in_data__36_, wbuf_entry_in_data__35_, wbuf_entry_in_data__34_, wbuf_entry_in_data__33_, wbuf_entry_in_data__32_, wbuf_entry_in_data__31_, wbuf_entry_in_data__30_, wbuf_entry_in_data__29_, wbuf_entry_in_data__28_, wbuf_entry_in_data__27_, wbuf_entry_in_data__26_, wbuf_entry_in_data__25_, wbuf_entry_in_data__24_, wbuf_entry_in_data__23_, wbuf_entry_in_data__22_, wbuf_entry_in_data__21_, wbuf_entry_in_data__20_, wbuf_entry_in_data__19_, wbuf_entry_in_data__18_, wbuf_entry_in_data__17_, wbuf_entry_in_data__16_, wbuf_entry_in_data__15_, wbuf_entry_in_data__14_, wbuf_entry_in_data__13_, wbuf_entry_in_data__12_, wbuf_entry_in_data__11_, wbuf_entry_in_data__10_, wbuf_entry_in_data__9_, wbuf_entry_in_data__8_, wbuf_entry_in_data__7_, wbuf_entry_in_data__6_, wbuf_entry_in_data__5_, wbuf_entry_in_data__4_, wbuf_entry_in_data__3_, wbuf_entry_in_data__2_, wbuf_entry_in_data__1_, wbuf_entry_in_data__0_, cache_req_o[39:8] }),
    .v_i(wbuf_v_li),
    .wbuf_entry_o({ wbuf_entry_out_snoop_, wbuf_entry_out_bank_sel__7_, wbuf_entry_out_bank_sel__6_, wbuf_entry_out_bank_sel__5_, wbuf_entry_out_bank_sel__4_, wbuf_entry_out_bank_sel__3_, wbuf_entry_out_bank_sel__2_, wbuf_entry_out_bank_sel__1_, wbuf_entry_out_bank_sel__0_, wbuf_data_mem_mask, wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_, wbuf_entry_out_caddr__31_, wbuf_entry_out_caddr__30_, wbuf_entry_out_caddr__29_, wbuf_entry_out_caddr__28_, wbuf_entry_out_caddr__27_, wbuf_entry_out_caddr__26_, wbuf_entry_out_caddr__25_, wbuf_entry_out_caddr__24_, wbuf_entry_out_caddr__23_, wbuf_entry_out_caddr__22_, wbuf_entry_out_caddr__21_, wbuf_entry_out_caddr__20_, wbuf_entry_out_caddr__19_, wbuf_entry_out_caddr__18_, wbuf_entry_out_caddr__17_, wbuf_entry_out_caddr__16_, wbuf_entry_out_caddr__15_, wbuf_entry_out_caddr__14_, wbuf_entry_out_caddr__13_, wbuf_entry_out_caddr__12_, wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_, wbuf_entry_out_caddr__2_, wbuf_entry_out_caddr__1_, wbuf_entry_out_caddr__0_ }),
    .v_o(wbuf_v_lo),
    .force_o(wbuf_force_lo),
    .yumi_i(wbuf_yumi_li),
    .data_mem_pkt_i(data_mem_pkt_i),
    .data_mem_pkt_v_i(data_mem_pkt_v_i),
    .tag_mem_pkt_i(tag_mem_pkt_i),
    .tag_mem_pkt_v_i(tag_mem_pkt_v_i),
    .stat_mem_pkt_i(stat_mem_pkt_i),
    .stat_mem_pkt_v_i(stat_mem_pkt_v_i),
    .snoop_match_o(wbuf_snoop_match_lo),
    .v_tl_i(v_tl_r),
    .addr_tl_i({ ptag_i[19:0], paddr_tl }),
    .data_tv_i(ld_data_dword_raw),
    .data_merged_o(ld_data_dword_merged)
  );

  assign N784 = decode_tv_r_amo_subop__3_ | decode_tv_r_amo_subop__2_;
  assign N785 = decode_tv_r_amo_subop__1_ | N783;
  assign N786 = N784 | N785;
  assign N789 = N788 | decode_tv_r_amo_subop__0_;
  assign N790 = N784 | N789;
  assign N792 = N788 | N783;
  assign N793 = N784 | N792;
  assign N796 = decode_tv_r_amo_subop__3_ | N795;
  assign N797 = decode_tv_r_amo_subop__1_ | decode_tv_r_amo_subop__0_;
  assign N798 = N796 | N797;
  assign N800 = N796 | N785;
  assign N802 = N796 | N789;
  assign N804 = N796 | N792;
  assign N807 = N806 | decode_tv_r_amo_subop__2_;
  assign N808 = N807 | N797;
  assign N810 = N807 | N785;
  assign N812 = N807 | N789;
  assign N814 = N807 | N792;
  assign N816 = decode_tv_r_amo_subop__3_ & decode_tv_r_amo_subop__2_;
  assign N817 = N806 & N795;
  assign N818 = N788 & N783;
  assign N819 = N817 & N818;

  bsg_dff_reset_width_p1
  cache_req_v_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(cache_req_yumi_i),
    .data_o(cache_req_metadata_v_o)
  );


  bsg_dff_0000000c
  cached_hit_reg
  (
    .clk_i(clk_i),
    .data_i({ way_v_tv_r, cache_req_o[115:115], load_hit_way_tv }),
    .data_o({ metadata_way_v_r, metadata_hit_r, metadata_hit_index_r })
  );


  bsg_priority_encode_00000008_1
  pe_invalid
  (
    .i({ _14_net__7_, _14_net__6_, _14_net__5_, _14_net__4_, _14_net__3_, _14_net__2_, _14_net__1_, _14_net__0_ }),
    .addr_o(metadata_invalid_way),
    .v_o(metadata_invalid_exist)
  );

  assign cache_req_metadata_o[0] = (N889)? stat_mem_o[0] : 
                                   (N891)? stat_mem_o[1] : 
                                   (N893)? stat_mem_o[2] : 
                                   (N895)? stat_mem_o[3] : 
                                   (N890)? stat_mem_o[4] : 
                                   (N892)? stat_mem_o[5] : 
                                   (N894)? stat_mem_o[6] : 
                                   (N896)? stat_mem_o[7] : 1'b0;

  bsg_decode_00000008
  tag_mem_way_decode
  (
    .i(tag_mem_pkt_i[28:26]),
    .o(tag_mem_way_one_hot)
  );

  assign N902 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N903 = tag_mem_pkt_i[1] | N901;
  assign N904 = N902 | N903;
  assign N907 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N908 = N906 | tag_mem_pkt_i[0];
  assign N909 = N907 | N908;
  assign N913 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N914 = N911 | N912;
  assign N915 = N913 | N914;
  assign N917 = N1529 & tag_mem_pkt_i[2];
  assign N920 = N1529 & N918;
  assign N921 = N920 & N919;
  assign N924 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N925 = tag_mem_pkt_i[1] | N923;
  assign N926 = N924 | N925;
  assign N929 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N930 = N928 | tag_mem_pkt_i[0];
  assign N931 = N929 | N930;
  assign N935 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N936 = N933 | N934;
  assign N937 = N935 | N936;
  assign N939 = N1529 & tag_mem_pkt_i[2];
  assign N942 = N1529 & N940;
  assign N943 = N942 & N941;
  assign N946 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N947 = tag_mem_pkt_i[1] | N945;
  assign N948 = N946 | N947;
  assign N951 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N952 = N950 | tag_mem_pkt_i[0];
  assign N953 = N951 | N952;
  assign N957 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N958 = N955 | N956;
  assign N959 = N957 | N958;
  assign N961 = N1529 & tag_mem_pkt_i[2];
  assign N964 = N1529 & N962;
  assign N965 = N964 & N963;
  assign N968 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N969 = tag_mem_pkt_i[1] | N967;
  assign N970 = N968 | N969;
  assign N973 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N974 = N972 | tag_mem_pkt_i[0];
  assign N975 = N973 | N974;
  assign N979 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N980 = N977 | N978;
  assign N981 = N979 | N980;
  assign N983 = N1529 & tag_mem_pkt_i[2];
  assign N986 = N1529 & N984;
  assign N987 = N986 & N985;
  assign N990 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N991 = tag_mem_pkt_i[1] | N989;
  assign N992 = N990 | N991;
  assign N995 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N996 = N994 | tag_mem_pkt_i[0];
  assign N997 = N995 | N996;
  assign N1001 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1002 = N999 | N1000;
  assign N1003 = N1001 | N1002;
  assign N1005 = N1529 & tag_mem_pkt_i[2];
  assign N1008 = N1529 & N1006;
  assign N1009 = N1008 & N1007;
  assign N1012 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1013 = tag_mem_pkt_i[1] | N1011;
  assign N1014 = N1012 | N1013;
  assign N1017 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1018 = N1016 | tag_mem_pkt_i[0];
  assign N1019 = N1017 | N1018;
  assign N1023 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1024 = N1021 | N1022;
  assign N1025 = N1023 | N1024;
  assign N1027 = N1529 & tag_mem_pkt_i[2];
  assign N1030 = N1529 & N1028;
  assign N1031 = N1030 & N1029;
  assign N1034 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1035 = tag_mem_pkt_i[1] | N1033;
  assign N1036 = N1034 | N1035;
  assign N1039 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1040 = N1038 | tag_mem_pkt_i[0];
  assign N1041 = N1039 | N1040;
  assign N1045 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1046 = N1043 | N1044;
  assign N1047 = N1045 | N1046;
  assign N1049 = N1529 & tag_mem_pkt_i[2];
  assign N1052 = N1529 & N1050;
  assign N1053 = N1052 & N1051;
  assign N1056 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1057 = tag_mem_pkt_i[1] | N1055;
  assign N1058 = N1056 | N1057;
  assign N1061 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1062 = N1060 | tag_mem_pkt_i[0];
  assign N1063 = N1061 | N1062;
  assign N1067 = tag_mem_fast_write | tag_mem_pkt_i[2];
  assign N1068 = N1065 | N1066;
  assign N1069 = N1067 | N1068;
  assign N1071 = N1529 & tag_mem_pkt_i[2];
  assign N1074 = N1529 & N1072;
  assign N1075 = N1074 & N1073;

  bsg_dff_width_p3
  tag_mem_pkt_way_reg
  (
    .clk_i(clk_i),
    .data_i(tag_mem_pkt_i[28:26]),
    .data_o(tag_mem_pkt_way_r)
  );

  assign tag_mem_o[22] = (N1084)? tag_mem_data_lo[22] : 
                         (N1086)? tag_mem_data_lo[45] : 
                         (N1088)? tag_mem_data_lo[68] : 
                         (N1090)? tag_mem_data_lo[91] : 
                         (N1085)? tag_mem_data_lo[114] : 
                         (N1087)? tag_mem_data_lo[137] : 
                         (N1089)? tag_mem_data_lo[160] : 
                         (N1091)? tag_mem_data_lo[183] : 1'b0;
  assign tag_mem_o[21] = (N1084)? tag_mem_data_lo[21] : 
                         (N1086)? tag_mem_data_lo[44] : 
                         (N1088)? tag_mem_data_lo[67] : 
                         (N1090)? tag_mem_data_lo[90] : 
                         (N1085)? tag_mem_data_lo[113] : 
                         (N1087)? tag_mem_data_lo[136] : 
                         (N1089)? tag_mem_data_lo[159] : 
                         (N1091)? tag_mem_data_lo[182] : 1'b0;
  assign tag_mem_o[20] = (N1084)? tag_mem_data_lo[20] : 
                         (N1086)? tag_mem_data_lo[43] : 
                         (N1088)? tag_mem_data_lo[66] : 
                         (N1090)? tag_mem_data_lo[89] : 
                         (N1085)? tag_mem_data_lo[112] : 
                         (N1087)? tag_mem_data_lo[135] : 
                         (N1089)? tag_mem_data_lo[158] : 
                         (N1091)? tag_mem_data_lo[181] : 1'b0;
  assign tag_mem_o[19] = (N1084)? tag_mem_data_lo[19] : 
                         (N1086)? tag_mem_data_lo[42] : 
                         (N1088)? tag_mem_data_lo[65] : 
                         (N1090)? tag_mem_data_lo[88] : 
                         (N1085)? tag_mem_data_lo[111] : 
                         (N1087)? tag_mem_data_lo[134] : 
                         (N1089)? tag_mem_data_lo[157] : 
                         (N1091)? tag_mem_data_lo[180] : 1'b0;
  assign tag_mem_o[18] = (N1084)? tag_mem_data_lo[18] : 
                         (N1086)? tag_mem_data_lo[41] : 
                         (N1088)? tag_mem_data_lo[64] : 
                         (N1090)? tag_mem_data_lo[87] : 
                         (N1085)? tag_mem_data_lo[110] : 
                         (N1087)? tag_mem_data_lo[133] : 
                         (N1089)? tag_mem_data_lo[156] : 
                         (N1091)? tag_mem_data_lo[179] : 1'b0;
  assign tag_mem_o[17] = (N1084)? tag_mem_data_lo[17] : 
                         (N1086)? tag_mem_data_lo[40] : 
                         (N1088)? tag_mem_data_lo[63] : 
                         (N1090)? tag_mem_data_lo[86] : 
                         (N1085)? tag_mem_data_lo[109] : 
                         (N1087)? tag_mem_data_lo[132] : 
                         (N1089)? tag_mem_data_lo[155] : 
                         (N1091)? tag_mem_data_lo[178] : 1'b0;
  assign tag_mem_o[16] = (N1084)? tag_mem_data_lo[16] : 
                         (N1086)? tag_mem_data_lo[39] : 
                         (N1088)? tag_mem_data_lo[62] : 
                         (N1090)? tag_mem_data_lo[85] : 
                         (N1085)? tag_mem_data_lo[108] : 
                         (N1087)? tag_mem_data_lo[131] : 
                         (N1089)? tag_mem_data_lo[154] : 
                         (N1091)? tag_mem_data_lo[177] : 1'b0;
  assign tag_mem_o[15] = (N1084)? tag_mem_data_lo[15] : 
                         (N1086)? tag_mem_data_lo[38] : 
                         (N1088)? tag_mem_data_lo[61] : 
                         (N1090)? tag_mem_data_lo[84] : 
                         (N1085)? tag_mem_data_lo[107] : 
                         (N1087)? tag_mem_data_lo[130] : 
                         (N1089)? tag_mem_data_lo[153] : 
                         (N1091)? tag_mem_data_lo[176] : 1'b0;
  assign tag_mem_o[14] = (N1084)? tag_mem_data_lo[14] : 
                         (N1086)? tag_mem_data_lo[37] : 
                         (N1088)? tag_mem_data_lo[60] : 
                         (N1090)? tag_mem_data_lo[83] : 
                         (N1085)? tag_mem_data_lo[106] : 
                         (N1087)? tag_mem_data_lo[129] : 
                         (N1089)? tag_mem_data_lo[152] : 
                         (N1091)? tag_mem_data_lo[175] : 1'b0;
  assign tag_mem_o[13] = (N1084)? tag_mem_data_lo[13] : 
                         (N1086)? tag_mem_data_lo[36] : 
                         (N1088)? tag_mem_data_lo[59] : 
                         (N1090)? tag_mem_data_lo[82] : 
                         (N1085)? tag_mem_data_lo[105] : 
                         (N1087)? tag_mem_data_lo[128] : 
                         (N1089)? tag_mem_data_lo[151] : 
                         (N1091)? tag_mem_data_lo[174] : 1'b0;
  assign tag_mem_o[12] = (N1084)? tag_mem_data_lo[12] : 
                         (N1086)? tag_mem_data_lo[35] : 
                         (N1088)? tag_mem_data_lo[58] : 
                         (N1090)? tag_mem_data_lo[81] : 
                         (N1085)? tag_mem_data_lo[104] : 
                         (N1087)? tag_mem_data_lo[127] : 
                         (N1089)? tag_mem_data_lo[150] : 
                         (N1091)? tag_mem_data_lo[173] : 1'b0;
  assign tag_mem_o[11] = (N1084)? tag_mem_data_lo[11] : 
                         (N1086)? tag_mem_data_lo[34] : 
                         (N1088)? tag_mem_data_lo[57] : 
                         (N1090)? tag_mem_data_lo[80] : 
                         (N1085)? tag_mem_data_lo[103] : 
                         (N1087)? tag_mem_data_lo[126] : 
                         (N1089)? tag_mem_data_lo[149] : 
                         (N1091)? tag_mem_data_lo[172] : 1'b0;
  assign tag_mem_o[10] = (N1084)? tag_mem_data_lo[10] : 
                         (N1086)? tag_mem_data_lo[33] : 
                         (N1088)? tag_mem_data_lo[56] : 
                         (N1090)? tag_mem_data_lo[79] : 
                         (N1085)? tag_mem_data_lo[102] : 
                         (N1087)? tag_mem_data_lo[125] : 
                         (N1089)? tag_mem_data_lo[148] : 
                         (N1091)? tag_mem_data_lo[171] : 1'b0;
  assign tag_mem_o[9] = (N1084)? tag_mem_data_lo[9] : 
                        (N1086)? tag_mem_data_lo[32] : 
                        (N1088)? tag_mem_data_lo[55] : 
                        (N1090)? tag_mem_data_lo[78] : 
                        (N1085)? tag_mem_data_lo[101] : 
                        (N1087)? tag_mem_data_lo[124] : 
                        (N1089)? tag_mem_data_lo[147] : 
                        (N1091)? tag_mem_data_lo[170] : 1'b0;
  assign tag_mem_o[8] = (N1084)? tag_mem_data_lo[8] : 
                        (N1086)? tag_mem_data_lo[31] : 
                        (N1088)? tag_mem_data_lo[54] : 
                        (N1090)? tag_mem_data_lo[77] : 
                        (N1085)? tag_mem_data_lo[100] : 
                        (N1087)? tag_mem_data_lo[123] : 
                        (N1089)? tag_mem_data_lo[146] : 
                        (N1091)? tag_mem_data_lo[169] : 1'b0;
  assign tag_mem_o[7] = (N1084)? tag_mem_data_lo[7] : 
                        (N1086)? tag_mem_data_lo[30] : 
                        (N1088)? tag_mem_data_lo[53] : 
                        (N1090)? tag_mem_data_lo[76] : 
                        (N1085)? tag_mem_data_lo[99] : 
                        (N1087)? tag_mem_data_lo[122] : 
                        (N1089)? tag_mem_data_lo[145] : 
                        (N1091)? tag_mem_data_lo[168] : 1'b0;
  assign tag_mem_o[6] = (N1084)? tag_mem_data_lo[6] : 
                        (N1086)? tag_mem_data_lo[29] : 
                        (N1088)? tag_mem_data_lo[52] : 
                        (N1090)? tag_mem_data_lo[75] : 
                        (N1085)? tag_mem_data_lo[98] : 
                        (N1087)? tag_mem_data_lo[121] : 
                        (N1089)? tag_mem_data_lo[144] : 
                        (N1091)? tag_mem_data_lo[167] : 1'b0;
  assign tag_mem_o[5] = (N1084)? tag_mem_data_lo[5] : 
                        (N1086)? tag_mem_data_lo[28] : 
                        (N1088)? tag_mem_data_lo[51] : 
                        (N1090)? tag_mem_data_lo[74] : 
                        (N1085)? tag_mem_data_lo[97] : 
                        (N1087)? tag_mem_data_lo[120] : 
                        (N1089)? tag_mem_data_lo[143] : 
                        (N1091)? tag_mem_data_lo[166] : 1'b0;
  assign tag_mem_o[4] = (N1084)? tag_mem_data_lo[4] : 
                        (N1086)? tag_mem_data_lo[27] : 
                        (N1088)? tag_mem_data_lo[50] : 
                        (N1090)? tag_mem_data_lo[73] : 
                        (N1085)? tag_mem_data_lo[96] : 
                        (N1087)? tag_mem_data_lo[119] : 
                        (N1089)? tag_mem_data_lo[142] : 
                        (N1091)? tag_mem_data_lo[165] : 1'b0;
  assign tag_mem_o[3] = (N1084)? tag_mem_data_lo[3] : 
                        (N1086)? tag_mem_data_lo[26] : 
                        (N1088)? tag_mem_data_lo[49] : 
                        (N1090)? tag_mem_data_lo[72] : 
                        (N1085)? tag_mem_data_lo[95] : 
                        (N1087)? tag_mem_data_lo[118] : 
                        (N1089)? tag_mem_data_lo[141] : 
                        (N1091)? tag_mem_data_lo[164] : 1'b0;
  assign tag_mem_o[2] = (N1084)? tag_mem_data_lo[2] : 
                        (N1086)? tag_mem_data_lo[25] : 
                        (N1088)? tag_mem_data_lo[48] : 
                        (N1090)? tag_mem_data_lo[71] : 
                        (N1085)? tag_mem_data_lo[94] : 
                        (N1087)? tag_mem_data_lo[117] : 
                        (N1089)? tag_mem_data_lo[140] : 
                        (N1091)? tag_mem_data_lo[163] : 1'b0;
  assign tag_mem_o[1] = (N1084)? tag_mem_data_lo[1] : 
                        (N1086)? tag_mem_data_lo[24] : 
                        (N1088)? tag_mem_data_lo[47] : 
                        (N1090)? tag_mem_data_lo[70] : 
                        (N1085)? tag_mem_data_lo[93] : 
                        (N1087)? tag_mem_data_lo[116] : 
                        (N1089)? tag_mem_data_lo[139] : 
                        (N1091)? tag_mem_data_lo[162] : 1'b0;
  assign tag_mem_o[0] = (N1084)? tag_mem_data_lo[0] : 
                        (N1086)? tag_mem_data_lo[23] : 
                        (N1088)? tag_mem_data_lo[46] : 
                        (N1090)? tag_mem_data_lo[69] : 
                        (N1085)? tag_mem_data_lo[92] : 
                        (N1087)? tag_mem_data_lo[115] : 
                        (N1089)? tag_mem_data_lo[138] : 
                        (N1091)? tag_mem_data_lo[161] : 1'b0;

  bsg_expand_bitmask_in_width_p4_expand_p2
  fill_mask_expand
  (
    .i(data_mem_pkt_i[5:2]),
    .o(data_mem_pkt_fill_mask_expanded)
  );


  bsg_rotate_left_00000008
  write_mask_rotate
  (
    .data_i(data_mem_pkt_fill_mask_expanded),
    .rot_i(data_mem_pkt_i[136:134]),
    .o(data_mem_write_bank_mask)
  );


  bsg_rotate_left_00000080
  write_data_rotate
  (
    .data_i(data_mem_pkt_i[133:6]),
    .rot_i({ data_mem_pkt_i[134:134], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .o(data_mem_pkt_fill_data_li)
  );


  bsg_dff_width_p3
  data_mem_pkt_way_reg
  (
    .clk_i(clk_i),
    .data_i(data_mem_pkt_i[136:134]),
    .data_o(data_mem_pkt_way_r)
  );


  bsg_rotate_right_00000200
  read_data_rotate
  (
    .data_i(data_mem_data_lo),
    .rot_i({ data_mem_pkt_way_r, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .o(data_mem_o)
  );


  bsg_lru_pseudo_tree_decode_00000008
  lru_decode
  (
    .way_id_i(lru_decode_way_li),
    .data_o(lru_decode_data_lo),
    .mask_o(lru_decode_mask_lo)
  );


  bsg_decode_with_v_00000008
  \tdm.dirty_mask_decode 
  (
    .i(\tdm.dirty_mask_way_li ),
    .v_i(\tdm.dirty_mask_v_li ),
    .o(dirty_mask_lo)
  );

  assign N1132 = N1513 & N1131;

  bsg_dff_width_p3
  stat_mem_pkt_way_reg
  (
    .clk_i(clk_i),
    .data_i(stat_mem_pkt_i[4:2]),
    .data_o(stat_mem_pkt_way_r)
  );

  assign N1144 = tag_mem_pkt_i[34:29] == \l1_lrsc.load_reserved_index_r ;
  assign N1145 = tag_mem_pkt_i[22:3] == \l1_lrsc.load_reserved_tag_r ;

  bsg_dff_reset_set_clear_width_p1_clear_over_set_p1
  \l1_lrsc.load_reserved_v_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .set_i(\l1_lrsc.set_reservation ),
    .clear_i(\l1_lrsc.clear_reservation ),
    .data_o(\l1_lrsc.load_reserved_v_r )
  );


  bsg_dff_en_0000001a
  \l1_lrsc.load_reserved_addr 
  (
    .clk_i(clk_i),
    .data_i(cache_req_o[39:14]),
    .en_i(\l1_lrsc.set_reservation ),
    .data_o({ \l1_lrsc.load_reserved_tag_r , \l1_lrsc.load_reserved_index_r  })
  );

  assign N1146 = \l1_lrsc.load_reserved_index_r  == cache_req_o[19:14];
  assign N1147 = \l1_lrsc.load_reserved_tag_r  == cache_req_o[39:20];

  bsg_counter_clear_up_max_val_p15_init_val_p0_disable_overflow_warning_p1
  \l1_lrsc.lrsc_lock_counter 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(sc_success_tv),
    .up_i(\l1_lrsc.lrsc_lock_up ),
    .count_o(\l1_lrsc.lrsc_lock_cnt )
  );


  bsg_dff_en_0000008a
  mshr_reg
  (
    .clk_i(clk_i),
    .data_i({ uncached_tv_r, amo64_reg_in, amo32_reg_in, cache_req_o[47:8], tag_o, decode_tv_r_load_op_, ret_o, decode_tv_r_store_op_, decode_tv_r_signed_op_, float_o, int_o, ptw_o, decode_tv_r_cache_op_, decode_tv_r_block_op_, decode_tv_r_double_op_, decode_tv_r_word_op_, decode_tv_r_half_op_, decode_tv_r_byte_op_, decode_tv_r_uncached_op_, decode_tv_r_lr_op_, decode_tv_r_sc_op_, decode_tv_r_amo_op_, decode_tv_r_clean_op_, decode_tv_r_inval_op_, decode_tv_r_bclean_op_, decode_tv_r_binval_op_, decode_tv_r_bzero_op_, decode_tv_r_amo_subop__3_, decode_tv_r_amo_subop__2_, decode_tv_r_amo_subop__1_, decode_tv_r_amo_subop__0_, rd_addr_o }),
    .en_i(blocking_sent),
    .data_o({ snoop_uncached, snoop_st_data, snoop_paddr, \hum.fill_index , snoop_paddr_5, snoop_paddr_4, snoop_paddr_3, snoop_paddr_2, snoop_paddr_1, snoop_paddr_0, snoop_decode })
  );

  assign { N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << data_mem_pkt_i[136:134];

  bsg_dff_reset_en_00000010
  \hum.fill_reg 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(_25_net_),
    .data_i({ \hum.fill_bank_mask_n , \hum.fill_hit_n  }),
    .data_o({ \hum.fill_bank_mask_r , \hum.fill_hit_r  })
  );

  assign N1178 = \hum.fill_index  == paddr_tl[11:6];
  assign { N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, data_mem_pkt_v_i } << data_mem_pkt_i[136:134];
  assign { N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tag_mem_pkt_v_i } << tag_mem_pkt_i[28:26];

  bsg_decode_00000008
  snoop_offset_decode
  (
    .i({ snoop_paddr_5, snoop_paddr_4, snoop_paddr_3 }),
    .o(snoop_bank_sel_one_hot)
  );

  assign N1195 = tag_mem_data_lo[182] | tag_mem_data_lo[183];
  assign N1196 = tag_mem_data_lo[181] | N1195;
  assign N1197 = tag_mem_data_lo[159] | tag_mem_data_lo[160];
  assign N1198 = tag_mem_data_lo[158] | N1197;
  assign N1199 = tag_mem_data_lo[136] | tag_mem_data_lo[137];
  assign N1200 = tag_mem_data_lo[135] | N1199;
  assign N1201 = tag_mem_data_lo[113] | tag_mem_data_lo[114];
  assign N1202 = tag_mem_data_lo[112] | N1201;
  assign N1203 = tag_mem_data_lo[90] | tag_mem_data_lo[91];
  assign N1204 = tag_mem_data_lo[89] | N1203;
  assign N1205 = tag_mem_data_lo[67] | tag_mem_data_lo[68];
  assign N1206 = tag_mem_data_lo[66] | N1205;
  assign N1207 = tag_mem_data_lo[44] | tag_mem_data_lo[45];
  assign N1208 = tag_mem_data_lo[43] | N1207;
  assign N1209 = tag_mem_data_lo[21] | tag_mem_data_lo[22];
  assign N1210 = tag_mem_data_lo[20] | N1209;
  assign N1211 = load_hit_way_tv[1] & load_hit_way_tv[2];
  assign N1212 = load_hit_way_tv[0] & N1211;
  assign N1213 = ~load_hit_way_tv[2];
  assign N1214 = ~load_hit_way_tv[1];
  assign N1215 = N1214 | N1213;
  assign N1216 = load_hit_way_tv[0] | N1215;
  assign N1217 = ~N1216;
  assign N1218 = ~load_hit_way_tv[2];
  assign N1219 = ~load_hit_way_tv[0];
  assign N1220 = load_hit_way_tv[1] | N1218;
  assign N1221 = N1219 | N1220;
  assign N1222 = ~N1221;
  assign N1223 = ~load_hit_way_tv[2];
  assign N1224 = load_hit_way_tv[1] | N1223;
  assign N1225 = load_hit_way_tv[0] | N1224;
  assign N1226 = ~N1225;
  assign N1227 = ~load_hit_way_tv[1];
  assign N1228 = ~load_hit_way_tv[0];
  assign N1229 = N1227 | load_hit_way_tv[2];
  assign N1230 = N1228 | N1229;
  assign N1231 = ~N1230;
  assign N1232 = ~load_hit_way_tv[1];
  assign N1233 = N1232 | load_hit_way_tv[2];
  assign N1234 = load_hit_way_tv[0] | N1233;
  assign N1235 = ~N1234;
  assign N1236 = ~load_hit_way_tv[0];
  assign N1237 = load_hit_way_tv[1] | load_hit_way_tv[2];
  assign N1238 = N1236 | N1237;
  assign N1239 = ~N1238;
  assign N1240 = load_hit_way_tv[1] | load_hit_way_tv[2];
  assign N1241 = load_hit_way_tv[0] | N1240;
  assign N1242 = ~N1241;
  assign N1243 = ~tag_mem_pkt_i[2];
  assign N1244 = tag_mem_pkt_i[1] | N1243;
  assign N1245 = tag_mem_pkt_i[0] | N1244;
  assign N1246 = ~N1245;
  assign N1247 = ~tag_mem_pkt_i[2];
  assign N1248 = tag_mem_pkt_i[1] | N1247;
  assign N1249 = tag_mem_pkt_i[0] | N1248;
  assign N1250 = ~data_mem_pkt_i[0];
  assign N1251 = N1250 | data_mem_pkt_i[1];
  assign N1252 = ~N1251;
  assign N1253 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1254 = ~N1253;
  assign N1255 = ~data_mem_pkt_i[0];
  assign N1256 = N1255 | data_mem_pkt_i[1];
  assign N1257 = ~N1256;
  assign N1258 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1259 = ~N1258;
  assign N1260 = ~data_mem_pkt_i[0];
  assign N1261 = N1260 | data_mem_pkt_i[1];
  assign N1262 = ~N1261;
  assign N1263 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1264 = ~N1263;
  assign N1265 = ~data_mem_pkt_i[0];
  assign N1266 = N1265 | data_mem_pkt_i[1];
  assign N1267 = ~N1266;
  assign N1268 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1269 = ~N1268;
  assign N1270 = ~data_mem_pkt_i[0];
  assign N1271 = N1270 | data_mem_pkt_i[1];
  assign N1272 = ~N1271;
  assign N1273 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1274 = ~N1273;
  assign N1275 = ~data_mem_pkt_i[0];
  assign N1276 = N1275 | data_mem_pkt_i[1];
  assign N1277 = ~N1276;
  assign N1278 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1279 = ~N1278;
  assign N1280 = ~data_mem_pkt_i[0];
  assign N1281 = N1280 | data_mem_pkt_i[1];
  assign N1282 = ~N1281;
  assign N1283 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1284 = ~N1283;
  assign N1285 = ~data_mem_pkt_i[0];
  assign N1286 = N1285 | data_mem_pkt_i[1];
  assign N1287 = ~N1286;
  assign N1288 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1289 = ~N1288;
  assign N1290 = ~stat_mem_pkt_i[0];
  assign N1291 = N1290 | stat_mem_pkt_i[1];
  assign N1292 = ~N1291;
  assign N1293 = ~stat_mem_pkt_i[0];
  assign N1294 = N1293 | stat_mem_pkt_i[1];
  assign N1295 = tag_mem_data_lo[182] | tag_mem_data_lo[183];
  assign N1296 = tag_mem_data_lo[181] | N1295;
  assign N1297 = tag_mem_data_lo[159] | tag_mem_data_lo[160];
  assign N1298 = tag_mem_data_lo[158] | N1297;
  assign N1299 = tag_mem_data_lo[136] | tag_mem_data_lo[137];
  assign N1300 = tag_mem_data_lo[135] | N1299;
  assign N1301 = tag_mem_data_lo[113] | tag_mem_data_lo[114];
  assign N1302 = tag_mem_data_lo[112] | N1301;
  assign N1303 = tag_mem_data_lo[90] | tag_mem_data_lo[91];
  assign N1304 = tag_mem_data_lo[89] | N1303;
  assign N1305 = tag_mem_data_lo[67] | tag_mem_data_lo[68];
  assign N1306 = tag_mem_data_lo[66] | N1305;
  assign N1307 = tag_mem_data_lo[44] | tag_mem_data_lo[45];
  assign N1308 = tag_mem_data_lo[43] | N1307;
  assign N1309 = tag_mem_data_lo[21] | tag_mem_data_lo[22];
  assign N1310 = tag_mem_data_lo[20] | N1309;
  assign N1311 = data_mem_pkt_i[0] | data_mem_pkt_i[1];
  assign N1312 = ~N1311;
  assign N1313 = ~stat_mem_pkt_i[0];
  assign N1314 = N1313 | stat_mem_pkt_i[1];
  assign N1315 = ~N1314;
  assign N1316 = \l1_lrsc.lrsc_lock_cnt [2] | \l1_lrsc.lrsc_lock_cnt [3];
  assign N1317 = \l1_lrsc.lrsc_lock_cnt [1] | N1316;
  assign N1318 = \l1_lrsc.lrsc_lock_cnt [0] | N1317;
  assign N1319 = ~data_mem_pkt_i[0];
  assign N1320 = N1319 | data_mem_pkt_i[1];
  assign N1321 = ~N1320;
  assign N1322 = ~data_mem_pkt_i[0];
  assign N1323 = N1322 | data_mem_pkt_i[1];
  assign N1324 = ~N1323;
  assign N1325 = state_r[0] | state_r[1];
  assign N1326 = ~N1325;
  assign N1327 = ~state_r[0];
  assign N1328 = N1327 | state_r[1];
  assign N1329 = ~N1328;
  assign \data_mem_lines_0_.data_mem_pkt_offset  = 1'b0 - data_mem_pkt_i[136:134];
  assign \data_mem_lines_1_.data_mem_pkt_offset  = 1'b1 - data_mem_pkt_i[136:134];
  assign \data_mem_lines_2_.data_mem_pkt_offset  = { 1'b1, 1'b0 } - data_mem_pkt_i[136:134];
  assign \data_mem_lines_3_.data_mem_pkt_offset  = { 1'b1, 1'b1 } - data_mem_pkt_i[136:134];
  assign \data_mem_lines_4_.data_mem_pkt_offset  = { 1'b1, 1'b0, 1'b0 } - data_mem_pkt_i[136:134];
  assign \data_mem_lines_5_.data_mem_pkt_offset  = { 1'b1, 1'b0, 1'b1 } - data_mem_pkt_i[136:134];
  assign \data_mem_lines_6_.data_mem_pkt_offset  = { 1'b1, 1'b1, 1'b0 } - data_mem_pkt_i[136:134];
  assign \data_mem_lines_7_.data_mem_pkt_offset  = { 1'b1, 1'b1, 1'b1 } - data_mem_pkt_i[136:134];
  assign { N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374 } = atomic_reg_data + atomic_mem_data;
  assign data_o = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                  (N173)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                  (N171)? final_data_tv : 1'b0;
  assign N0 = N169;
  assign atomic_reg_data = (N1)? { amo64_reg_in, amo32_reg_in } : 
                           (N175)? { amo32_reg_in, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = N174;
  assign atomic_mem_data = (N2)? final_data_tv : 
                           (N177)? { final_data_tv[31:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2 = N176;
  assign { N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440 } = (N3)? atomic_reg_data : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N439)? atomic_mem_data : 1'b0;
  assign N3 = N438;
  assign { N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506 } = (N4)? atomic_reg_data : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N505)? atomic_mem_data : 1'b0;
  assign N4 = N504;
  assign { N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572 } = (N5)? atomic_reg_data : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N571)? atomic_mem_data : 1'b0;
  assign N5 = N570;
  assign { N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638 } = (N6)? atomic_reg_data : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N637)? atomic_mem_data : 1'b0;
  assign N6 = N636;
  assign { N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702 } = (N7)? { N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N8)? { N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N9)? { N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N10)? { N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N11)? { N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N12)? { N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N13)? { N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N14)? { N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N15)? atomic_reg_data : 1'b0;
  assign N7 = N803;
  assign N8 = N805;
  assign N9 = N801;
  assign N10 = N799;
  assign N11 = N809;
  assign N12 = N811;
  assign N13 = N813;
  assign N14 = N815;
  assign N15 = N181;
  assign atomic_alu_result = (N16)? { N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702 } : 
                             (N17)? atomic_reg_data : 1'b0;
  assign N16 = N178;
  assign N17 = N179;
  assign atomic_result = (N18)? atomic_alu_result : 
                         (N845)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, atomic_alu_result[63:32] } : 1'b0;
  assign N18 = N771;
  assign \wbuf_in_2_.slice_data  = (N19)? atomic_result[31:0] : 
                                   (N767)? amo32_reg_in : 1'b0;
  assign N19 = N766;
  assign \wbuf_in_3_.slice_data  = (N20)? atomic_result : 
                                   (N768)? { amo64_reg_in, amo32_reg_in } : 1'b0;
  assign N20 = N782;
  assign cache_req_o[114:51] = (N21)? { wbuf_entry_in_data__63_, wbuf_entry_in_data__62_, wbuf_entry_in_data__61_, wbuf_entry_in_data__60_, wbuf_entry_in_data__59_, wbuf_entry_in_data__58_, wbuf_entry_in_data__57_, wbuf_entry_in_data__56_, wbuf_entry_in_data__55_, wbuf_entry_in_data__54_, wbuf_entry_in_data__53_, wbuf_entry_in_data__52_, wbuf_entry_in_data__51_, wbuf_entry_in_data__50_, wbuf_entry_in_data__49_, wbuf_entry_in_data__48_, wbuf_entry_in_data__47_, wbuf_entry_in_data__46_, wbuf_entry_in_data__45_, wbuf_entry_in_data__44_, wbuf_entry_in_data__43_, wbuf_entry_in_data__42_, wbuf_entry_in_data__41_, wbuf_entry_in_data__40_, wbuf_entry_in_data__39_, wbuf_entry_in_data__38_, wbuf_entry_in_data__37_, wbuf_entry_in_data__36_, wbuf_entry_in_data__35_, wbuf_entry_in_data__34_, wbuf_entry_in_data__33_, wbuf_entry_in_data__32_, wbuf_entry_in_data__31_, wbuf_entry_in_data__30_, wbuf_entry_in_data__29_, wbuf_entry_in_data__28_, wbuf_entry_in_data__27_, wbuf_entry_in_data__26_, wbuf_entry_in_data__25_, wbuf_entry_in_data__24_, wbuf_entry_in_data__23_, wbuf_entry_in_data__22_, wbuf_entry_in_data__21_, wbuf_entry_in_data__20_, wbuf_entry_in_data__19_, wbuf_entry_in_data__18_, wbuf_entry_in_data__17_, wbuf_entry_in_data__16_, wbuf_entry_in_data__15_, wbuf_entry_in_data__14_, wbuf_entry_in_data__13_, wbuf_entry_in_data__12_, wbuf_entry_in_data__11_, wbuf_entry_in_data__10_, wbuf_entry_in_data__9_, wbuf_entry_in_data__8_, wbuf_entry_in_data__7_, wbuf_entry_in_data__6_, wbuf_entry_in_data__5_, wbuf_entry_in_data__4_, wbuf_entry_in_data__3_, wbuf_entry_in_data__2_, wbuf_entry_in_data__1_, wbuf_entry_in_data__0_ } : 
                               (N22)? { amo64_reg_in, amo32_reg_in } : 1'b0;
  assign N21 = nonblocking_req;
  assign N22 = N1439;
  assign cache_req_o[48] = (N23)? 1'b0 : 
                           (N841)? 1'b0 : 
                           (N844)? 1'b1 : 
                           (N847)? 1'b0 : 
                           (N850)? 1'b1 : 
                           (N778)? 1'b0 : 
                           (N24)? 1'b0 : 1'b0;
  assign N23 = N769;
  assign N24 = 1'b0;
  assign cache_req_o[49] = (N23)? 1'b1 : 
                           (N841)? 1'b1 : 
                           (N844)? 1'b1 : 
                           (N847)? 1'b1 : 
                           (N779)? 1'b0 : 
                           (N24)? 1'b0 : 
                           (N24)? 1'b0 : 1'b0;
  assign cache_req_o[50] = (N23)? 1'b1 : 
                           (N841)? 1'b1 : 
                           (N780)? 1'b0 : 
                           (N24)? 1'b0 : 
                           (N24)? 1'b0 : 
                           (N24)? 1'b0 : 
                           (N24)? 1'b0 : 1'b0;
  assign { N824, N823, N822, N821 } = (N25)? { 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                      (N26)? { 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                      (N27)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                      (N10)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                      (N9)? { 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                      (N7)? { 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                      (N8)? { 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                      (N11)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                      (N12)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                                      (N13)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                                      (N14)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                      (N28)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N25 = N787;
  assign N26 = N791;
  assign N27 = N794;
  assign N28 = N820;
  assign cache_req_o[3:0] = (N20)? { N824, N823, N822, N821 } : 
                            (N29)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N29 = N781;
  assign cache_req_o[5:4] = (N30)? { 1'b0, 1'b1 } : 
                            (N852)? { 1'b1, 1'b1 } : 
                            (N855)? { 1'b0, 1'b0 } : 
                            (N858)? { 1'b1, 1'b1 } : 
                            (N861)? { 1'b1, 1'b0 } : 
                            (N864)? { 1'b0, 1'b0 } : 
                            (N867)? { 1'b0, 1'b1 } : 
                            (N870)? { 1'b0, 1'b0 } : 
                            (N873)? { 1'b0, 1'b1 } : 
                            (N876)? { 1'b0, 1'b0 } : 
                            (N879)? { 1'b1, 1'b1 } : 
                            (N837)? { 1'b1, 1'b0 } : 1'b0;
  assign N30 = N825;
  assign cache_req_o[6] = (N30)? 1'b1 : 
                          (N852)? 1'b0 : 
                          (N855)? 1'b1 : 
                          (N858)? 1'b1 : 
                          (N861)? 1'b1 : 
                          (N864)? 1'b0 : 
                          (N867)? 1'b0 : 
                          (N870)? 1'b0 : 
                          (N873)? 1'b1 : 
                          (N876)? 1'b1 : 
                          (N838)? 1'b0 : 
                          (N24)? 1'b0 : 1'b0;
  assign cache_req_o[7] = (N30)? 1'b1 : 
                          (N852)? 1'b1 : 
                          (N855)? 1'b1 : 
                          (N858)? 1'b0 : 
                          (N861)? 1'b0 : 
                          (N864)? 1'b1 : 
                          (N839)? 1'b0 : 
                          (N24)? 1'b0 : 
                          (N24)? 1'b0 : 
                          (N24)? 1'b0 : 
                          (N24)? 1'b0 : 
                          (N24)? 1'b0 : 1'b0;
  assign lru_way_li = (N31)? metadata_invalid_way : 
                      (N32)? lru_encode : 1'b0;
  assign N31 = metadata_invalid_exist;
  assign N32 = N880;
  assign cache_req_metadata_o[3:1] = (N33)? metadata_hit_index_r : 
                                     (N34)? lru_way_li : 1'b0;
  assign N33 = metadata_hit_r;
  assign N34 = N881;
  assign tag_mem_addr_li = (N35)? cache_req_o[19:14] : 
                           (N900)? dcache_pkt_i[11:6] : 
                           (N898)? tag_mem_pkt_i[34:29] : 1'b0;
  assign N35 = tag_mem_fast_write;
  assign tag_mem_data_li[22:0] = (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N36)? tag_mem_pkt_i[25:3] : 
                                 (N37)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N38)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N39)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N36 = N905;
  assign N37 = N910;
  assign N38 = N916;
  assign N39 = N922;
  assign tag_mem_mask_li[22:0] = (N35)? { N1242, N1242, N1242, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N36)? { tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0] } : 
                                 (N37)? { tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], tag_mem_way_one_hot[0:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N38)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N39)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[45:23] = (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N40)? tag_mem_pkt_i[25:3] : 
                                  (N41)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N42)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N43)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N40 = N927;
  assign N41 = N932;
  assign N42 = N938;
  assign N43 = N944;
  assign tag_mem_mask_li[45:23] = (N35)? { N1239, N1239, N1239, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N40)? { tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1] } : 
                                  (N41)? { tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], tag_mem_way_one_hot[1:1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N42)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N43)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[68:46] = (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N44)? tag_mem_pkt_i[25:3] : 
                                  (N45)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N46)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N47)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N44 = N949;
  assign N45 = N954;
  assign N46 = N960;
  assign N47 = N966;
  assign tag_mem_mask_li[68:46] = (N35)? { N1235, N1235, N1235, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N44)? { tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2] } : 
                                  (N45)? { tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], tag_mem_way_one_hot[2:2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N46)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N47)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[91:69] = (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N48)? tag_mem_pkt_i[25:3] : 
                                  (N49)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N50)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N51)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N48 = N971;
  assign N49 = N976;
  assign N50 = N982;
  assign N51 = N988;
  assign tag_mem_mask_li[91:69] = (N35)? { N1231, N1231, N1231, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N48)? { tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3] } : 
                                  (N49)? { tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], tag_mem_way_one_hot[3:3], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N50)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N51)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[114:92] = (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N52)? tag_mem_pkt_i[25:3] : 
                                   (N53)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N54)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N55)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N52 = N993;
  assign N53 = N998;
  assign N54 = N1004;
  assign N55 = N1010;
  assign tag_mem_mask_li[114:92] = (N35)? { N1226, N1226, N1226, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N52)? { tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4] } : 
                                   (N53)? { tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], tag_mem_way_one_hot[4:4], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N54)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N55)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[137:115] = (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N56)? tag_mem_pkt_i[25:3] : 
                                    (N57)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N58)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N59)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N56 = N1015;
  assign N57 = N1020;
  assign N58 = N1026;
  assign N59 = N1032;
  assign tag_mem_mask_li[137:115] = (N35)? { N1222, N1222, N1222, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N56)? { tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5] } : 
                                    (N57)? { tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], tag_mem_way_one_hot[5:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N58)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N59)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[160:138] = (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N60)? tag_mem_pkt_i[25:3] : 
                                    (N61)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N62)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N63)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N60 = N1037;
  assign N61 = N1042;
  assign N62 = N1048;
  assign N63 = N1054;
  assign tag_mem_mask_li[160:138] = (N35)? { N1217, N1217, N1217, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N60)? { tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6] } : 
                                    (N61)? { tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], tag_mem_way_one_hot[6:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N62)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N63)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tag_mem_data_li[183:161] = (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N64)? tag_mem_pkt_i[25:3] : 
                                    (N65)? { tag_mem_pkt_i[25:23], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N66)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N67)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N64 = N1059;
  assign N65 = N1064;
  assign N66 = N1070;
  assign N67 = N1076;
  assign tag_mem_mask_li[183:161] = (N35)? { N1212, N1212, N1212, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N64)? { tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7] } : 
                                    (N65)? { tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], tag_mem_way_one_hot[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N66)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N67)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign data_mem_mask_li[7:0] = (N68)? wbuf_data_mem_mask : 
                                 (N1092)? { data_mem_write_bank_mask[0:0], data_mem_write_bank_mask[0:0], data_mem_write_bank_mask[0:0], data_mem_write_bank_mask[0:0], data_mem_write_bank_mask[0:0], data_mem_write_bank_mask[0:0], data_mem_write_bank_mask[0:0], data_mem_write_bank_mask[0:0] } : 1'b0;
  assign N68 = data_mem_fast_write[0];
  assign data_mem_addr_li[8:0] = (N68)? { wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_ } : 
                                 (N1095)? dcache_pkt_i[11:3] : 
                                 (N1094)? { data_mem_pkt_i[142:137], \data_mem_lines_0_.data_mem_pkt_offset  } : 1'b0;
  assign data_mem_data_li[63:0] = (N68)? { wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_ } : 
                                  (N1092)? data_mem_pkt_fill_data_li[63:0] : 1'b0;
  assign data_mem_mask_li[15:8] = (N69)? wbuf_data_mem_mask : 
                                  (N1096)? { data_mem_write_bank_mask[1:1], data_mem_write_bank_mask[1:1], data_mem_write_bank_mask[1:1], data_mem_write_bank_mask[1:1], data_mem_write_bank_mask[1:1], data_mem_write_bank_mask[1:1], data_mem_write_bank_mask[1:1], data_mem_write_bank_mask[1:1] } : 1'b0;
  assign N69 = data_mem_fast_write[1];
  assign data_mem_addr_li[17:9] = (N69)? { wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_ } : 
                                  (N1099)? dcache_pkt_i[11:3] : 
                                  (N1098)? { data_mem_pkt_i[142:137], \data_mem_lines_1_.data_mem_pkt_offset  } : 1'b0;
  assign data_mem_data_li[127:64] = (N69)? { wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_ } : 
                                    (N1096)? data_mem_pkt_fill_data_li[127:64] : 1'b0;
  assign data_mem_mask_li[23:16] = (N70)? wbuf_data_mem_mask : 
                                   (N1100)? { data_mem_write_bank_mask[2:2], data_mem_write_bank_mask[2:2], data_mem_write_bank_mask[2:2], data_mem_write_bank_mask[2:2], data_mem_write_bank_mask[2:2], data_mem_write_bank_mask[2:2], data_mem_write_bank_mask[2:2], data_mem_write_bank_mask[2:2] } : 1'b0;
  assign N70 = data_mem_fast_write[2];
  assign data_mem_addr_li[26:18] = (N70)? { wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_ } : 
                                   (N1103)? dcache_pkt_i[11:3] : 
                                   (N1102)? { data_mem_pkt_i[142:137], \data_mem_lines_2_.data_mem_pkt_offset  } : 1'b0;
  assign data_mem_data_li[191:128] = (N70)? { wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_ } : 
                                     (N1100)? data_mem_pkt_fill_data_li[63:0] : 1'b0;
  assign data_mem_mask_li[31:24] = (N71)? wbuf_data_mem_mask : 
                                   (N1104)? { data_mem_write_bank_mask[3:3], data_mem_write_bank_mask[3:3], data_mem_write_bank_mask[3:3], data_mem_write_bank_mask[3:3], data_mem_write_bank_mask[3:3], data_mem_write_bank_mask[3:3], data_mem_write_bank_mask[3:3], data_mem_write_bank_mask[3:3] } : 1'b0;
  assign N71 = data_mem_fast_write[3];
  assign data_mem_addr_li[35:27] = (N71)? { wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_ } : 
                                   (N1107)? dcache_pkt_i[11:3] : 
                                   (N1106)? { data_mem_pkt_i[142:137], \data_mem_lines_3_.data_mem_pkt_offset  } : 1'b0;
  assign data_mem_data_li[255:192] = (N71)? { wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_ } : 
                                     (N1104)? data_mem_pkt_fill_data_li[127:64] : 1'b0;
  assign data_mem_mask_li[39:32] = (N72)? wbuf_data_mem_mask : 
                                   (N1108)? { data_mem_write_bank_mask[4:4], data_mem_write_bank_mask[4:4], data_mem_write_bank_mask[4:4], data_mem_write_bank_mask[4:4], data_mem_write_bank_mask[4:4], data_mem_write_bank_mask[4:4], data_mem_write_bank_mask[4:4], data_mem_write_bank_mask[4:4] } : 1'b0;
  assign N72 = data_mem_fast_write[4];
  assign data_mem_addr_li[44:36] = (N72)? { wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_ } : 
                                   (N1111)? dcache_pkt_i[11:3] : 
                                   (N1110)? { data_mem_pkt_i[142:137], \data_mem_lines_4_.data_mem_pkt_offset  } : 1'b0;
  assign data_mem_data_li[319:256] = (N72)? { wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_ } : 
                                     (N1108)? data_mem_pkt_fill_data_li[63:0] : 1'b0;
  assign data_mem_mask_li[47:40] = (N73)? wbuf_data_mem_mask : 
                                   (N1112)? { data_mem_write_bank_mask[5:5], data_mem_write_bank_mask[5:5], data_mem_write_bank_mask[5:5], data_mem_write_bank_mask[5:5], data_mem_write_bank_mask[5:5], data_mem_write_bank_mask[5:5], data_mem_write_bank_mask[5:5], data_mem_write_bank_mask[5:5] } : 1'b0;
  assign N73 = data_mem_fast_write[5];
  assign data_mem_addr_li[53:45] = (N73)? { wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_ } : 
                                   (N1115)? dcache_pkt_i[11:3] : 
                                   (N1114)? { data_mem_pkt_i[142:137], \data_mem_lines_5_.data_mem_pkt_offset  } : 1'b0;
  assign data_mem_data_li[383:320] = (N73)? { wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_ } : 
                                     (N1112)? data_mem_pkt_fill_data_li[127:64] : 1'b0;
  assign data_mem_mask_li[55:48] = (N74)? wbuf_data_mem_mask : 
                                   (N1116)? { data_mem_write_bank_mask[6:6], data_mem_write_bank_mask[6:6], data_mem_write_bank_mask[6:6], data_mem_write_bank_mask[6:6], data_mem_write_bank_mask[6:6], data_mem_write_bank_mask[6:6], data_mem_write_bank_mask[6:6], data_mem_write_bank_mask[6:6] } : 1'b0;
  assign N74 = data_mem_fast_write[6];
  assign data_mem_addr_li[62:54] = (N74)? { wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_ } : 
                                   (N1119)? dcache_pkt_i[11:3] : 
                                   (N1118)? { data_mem_pkt_i[142:137], \data_mem_lines_6_.data_mem_pkt_offset  } : 1'b0;
  assign data_mem_data_li[447:384] = (N74)? { wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_ } : 
                                     (N1116)? data_mem_pkt_fill_data_li[63:0] : 1'b0;
  assign data_mem_mask_li[63:56] = (N75)? wbuf_data_mem_mask : 
                                   (N1120)? { data_mem_write_bank_mask[7:7], data_mem_write_bank_mask[7:7], data_mem_write_bank_mask[7:7], data_mem_write_bank_mask[7:7], data_mem_write_bank_mask[7:7], data_mem_write_bank_mask[7:7], data_mem_write_bank_mask[7:7], data_mem_write_bank_mask[7:7] } : 1'b0;
  assign N75 = data_mem_fast_write[7];
  assign data_mem_addr_li[71:63] = (N75)? { wbuf_entry_out_caddr__11_, wbuf_entry_out_caddr__10_, wbuf_entry_out_caddr__9_, wbuf_entry_out_caddr__8_, wbuf_entry_out_caddr__7_, wbuf_entry_out_caddr__6_, wbuf_entry_out_caddr__5_, wbuf_entry_out_caddr__4_, wbuf_entry_out_caddr__3_ } : 
                                   (N1123)? dcache_pkt_i[11:3] : 
                                   (N1122)? { data_mem_pkt_i[142:137], \data_mem_lines_7_.data_mem_pkt_offset  } : 1'b0;
  assign data_mem_data_li[511:448] = (N75)? { wbuf_entry_out_data__63_, wbuf_entry_out_data__62_, wbuf_entry_out_data__61_, wbuf_entry_out_data__60_, wbuf_entry_out_data__59_, wbuf_entry_out_data__58_, wbuf_entry_out_data__57_, wbuf_entry_out_data__56_, wbuf_entry_out_data__55_, wbuf_entry_out_data__54_, wbuf_entry_out_data__53_, wbuf_entry_out_data__52_, wbuf_entry_out_data__51_, wbuf_entry_out_data__50_, wbuf_entry_out_data__49_, wbuf_entry_out_data__48_, wbuf_entry_out_data__47_, wbuf_entry_out_data__46_, wbuf_entry_out_data__45_, wbuf_entry_out_data__44_, wbuf_entry_out_data__43_, wbuf_entry_out_data__42_, wbuf_entry_out_data__41_, wbuf_entry_out_data__40_, wbuf_entry_out_data__39_, wbuf_entry_out_data__38_, wbuf_entry_out_data__37_, wbuf_entry_out_data__36_, wbuf_entry_out_data__35_, wbuf_entry_out_data__34_, wbuf_entry_out_data__33_, wbuf_entry_out_data__32_, wbuf_entry_out_data__31_, wbuf_entry_out_data__30_, wbuf_entry_out_data__29_, wbuf_entry_out_data__28_, wbuf_entry_out_data__27_, wbuf_entry_out_data__26_, wbuf_entry_out_data__25_, wbuf_entry_out_data__24_, wbuf_entry_out_data__23_, wbuf_entry_out_data__22_, wbuf_entry_out_data__21_, wbuf_entry_out_data__20_, wbuf_entry_out_data__19_, wbuf_entry_out_data__18_, wbuf_entry_out_data__17_, wbuf_entry_out_data__16_, wbuf_entry_out_data__15_, wbuf_entry_out_data__14_, wbuf_entry_out_data__13_, wbuf_entry_out_data__12_, wbuf_entry_out_data__11_, wbuf_entry_out_data__10_, wbuf_entry_out_data__9_, wbuf_entry_out_data__8_, wbuf_entry_out_data__7_, wbuf_entry_out_data__6_, wbuf_entry_out_data__5_, wbuf_entry_out_data__4_, wbuf_entry_out_data__3_, wbuf_entry_out_data__2_, wbuf_entry_out_data__1_, wbuf_entry_out_data__0_ } : 
                                     (N1120)? data_mem_pkt_fill_data_li[127:64] : 1'b0;
  assign stat_mem_addr_li = (N76)? cache_req_o[19:14] : 
                            (N1125)? stat_mem_pkt_i[10:5] : 1'b0;
  assign N76 = N1124;
  assign { N1130, N1129, N1128 } = (N77)? store_hit_way_tv : 
                                   (N1127)? load_hit_way_tv : 1'b0;
  assign N77 = N1126;
  assign lru_decode_way_li = (N78)? { N1130, N1129, N1128 } : 
                             (N79)? stat_mem_pkt_i[4:2] : 1'b0;
  assign N78 = v_tv_r;
  assign N79 = N1513;
  assign \tdm.dirty_mask_way_li  = (N78)? store_hit_way_tv : 
                                   (N79)? stat_mem_pkt_i[4:2] : 1'b0;
  assign { N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136 } = (N80)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                      (N81)? dirty_mask_lo : 1'b0;
  assign N80 = N1134;
  assign N81 = N1135;
  assign stat_mem_data_li[0] = ~N1132;
  assign stat_mem_data_li[1] = ~N1132;
  assign stat_mem_data_li[2] = ~N1132;
  assign stat_mem_data_li[3] = ~N1132;
  assign stat_mem_data_li[4] = ~N1132;
  assign stat_mem_data_li[5] = ~N1132;
  assign stat_mem_data_li[6] = ~N1132;
  assign stat_mem_data_li[7] = ~N1132;
  assign stat_mem_data_li[14:8] = (N82)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N1133)? lru_decode_data_lo : 1'b0;
  assign N82 = N1132;
  assign stat_mem_mask_li = (N82)? { N1134, N1134, N1134, N1134, N1134, N1134, N1134, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136 } : 
                            (N1133)? { lru_decode_mask_lo, dirty_mask_lo } : 1'b0;
  assign N1154 = ~N1155;
  assign state_n = (N83)? { 1'b0, 1'b0 } : 
                   (N1157)? { N1155, N1154 } : 
                   (N1160)? { 1'b1, 1'b0 } : 
                   (N1153)? state_r : 1'b0;
  assign N83 = N1148;
  assign \hum.fill_bank_mask_n  = (N84)? { N1162, N1163, N1164, N1165, N1166, N1167, N1168, N1169 } : 
                                  (N85)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N84 = \hum.fill_v ;
  assign N85 = N1161;
  assign \hum.fill_hit_n  = (N84)? { N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170 } : 
                            (N85)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N1330 = N86 & decode_tv_r_amo_subop__0_;
  assign N86 = ~decode_tv_r_amo_subop__1_;
  assign N1331 = N1330 | decode_tv_r_amo_subop__1_;
  assign N1332 = N87 & N1331;
  assign N87 = ~decode_tv_r_amo_subop__2_;
  assign N1333 = N1332 | decode_tv_r_amo_subop__2_;
  assign N1334 = ~decode_tv_r_amo_subop__2_;
  assign N1335 = N88 & N1333;
  assign N88 = ~decode_tv_r_amo_subop__3_;
  assign N1336 = decode_tv_r_amo_subop__3_ & N1334;
  assign N178 = N1335 | N1336;
  assign flush_tv = N1339 | fill_hazard;
  assign N1339 = N1338 | nonblocking_hazard;
  assign N1338 = N1337 | blocking_hazard;
  assign N1337 = flush_i | tag_mem_fast_write;
  assign flush_tl = flush_tv | data_mem_write_hazard;
  assign critical_recv = N1345 & N1347;
  assign N1345 = N1342 & N1344;
  assign N1342 = cache_req_critical_i & N1341;
  assign N1341 = N1340 | stat_mem_pkt_yumi_o;
  assign N1340 = ~stat_mem_pkt_v_i;
  assign N1344 = N1343 | tag_mem_pkt_yumi_o;
  assign N1343 = ~tag_mem_pkt_v_i;
  assign N1347 = N1346 | data_mem_pkt_yumi_o;
  assign N1346 = ~data_mem_pkt_v_i;
  assign complete_recv = N1353 & N1355;
  assign N1353 = N1350 & N1352;
  assign N1350 = cache_req_last_i & N1349;
  assign N1349 = N1348 | stat_mem_pkt_yumi_o;
  assign N1348 = ~stat_mem_pkt_v_i;
  assign N1352 = N1351 | tag_mem_pkt_yumi_o;
  assign N1351 = ~tag_mem_pkt_v_i;
  assign N1355 = N1354 | data_mem_pkt_yumi_o;
  assign N1354 = ~data_mem_pkt_v_i;
  assign safe_tl_we = v_i & N1356;
  assign N1356 = ~busy_o;
  assign tl_we = safe_tl_we & N1357;
  assign N1357 = ~flush_tl;
  assign \tag_comp_tl_0_.tag_match_tl  = N1366 & N89;
  assign N1366 = ptag_v_i & N1365;
  assign N1365 = ~N1364;
  assign N1364 = N1363 | ptag_i[20];
  assign N1363 = N1362 | ptag_i[21];
  assign N1362 = N1361 | ptag_i[22];
  assign N1361 = N1360 | ptag_i[23];
  assign N1360 = N1359 | ptag_i[24];
  assign N1359 = N1358 | ptag_i[25];
  assign N1358 = ptag_i[27] | ptag_i[26];
  assign load_hit_tl[0] = \tag_comp_tl_0_.tag_match_tl  & N1310;
  assign store_hit_tl[0] = \tag_comp_tl_0_.tag_match_tl  & N98;
  assign \tag_comp_tl_1_.tag_match_tl  = N1375 & N99;
  assign N1375 = ptag_v_i & N1374;
  assign N1374 = ~N1373;
  assign N1373 = N1372 | ptag_i[20];
  assign N1372 = N1371 | ptag_i[21];
  assign N1371 = N1370 | ptag_i[22];
  assign N1370 = N1369 | ptag_i[23];
  assign N1369 = N1368 | ptag_i[24];
  assign N1368 = N1367 | ptag_i[25];
  assign N1367 = ptag_i[27] | ptag_i[26];
  assign load_hit_tl[1] = \tag_comp_tl_1_.tag_match_tl  & N1308;
  assign store_hit_tl[1] = \tag_comp_tl_1_.tag_match_tl  & N108;
  assign \tag_comp_tl_2_.tag_match_tl  = N1384 & N109;
  assign N1384 = ptag_v_i & N1383;
  assign N1383 = ~N1382;
  assign N1382 = N1381 | ptag_i[20];
  assign N1381 = N1380 | ptag_i[21];
  assign N1380 = N1379 | ptag_i[22];
  assign N1379 = N1378 | ptag_i[23];
  assign N1378 = N1377 | ptag_i[24];
  assign N1377 = N1376 | ptag_i[25];
  assign N1376 = ptag_i[27] | ptag_i[26];
  assign load_hit_tl[2] = \tag_comp_tl_2_.tag_match_tl  & N1306;
  assign store_hit_tl[2] = \tag_comp_tl_2_.tag_match_tl  & N118;
  assign \tag_comp_tl_3_.tag_match_tl  = N1393 & N119;
  assign N1393 = ptag_v_i & N1392;
  assign N1392 = ~N1391;
  assign N1391 = N1390 | ptag_i[20];
  assign N1390 = N1389 | ptag_i[21];
  assign N1389 = N1388 | ptag_i[22];
  assign N1388 = N1387 | ptag_i[23];
  assign N1387 = N1386 | ptag_i[24];
  assign N1386 = N1385 | ptag_i[25];
  assign N1385 = ptag_i[27] | ptag_i[26];
  assign load_hit_tl[3] = \tag_comp_tl_3_.tag_match_tl  & N1304;
  assign store_hit_tl[3] = \tag_comp_tl_3_.tag_match_tl  & N128;
  assign \tag_comp_tl_4_.tag_match_tl  = N1402 & N129;
  assign N1402 = ptag_v_i & N1401;
  assign N1401 = ~N1400;
  assign N1400 = N1399 | ptag_i[20];
  assign N1399 = N1398 | ptag_i[21];
  assign N1398 = N1397 | ptag_i[22];
  assign N1397 = N1396 | ptag_i[23];
  assign N1396 = N1395 | ptag_i[24];
  assign N1395 = N1394 | ptag_i[25];
  assign N1394 = ptag_i[27] | ptag_i[26];
  assign load_hit_tl[4] = \tag_comp_tl_4_.tag_match_tl  & N1302;
  assign store_hit_tl[4] = \tag_comp_tl_4_.tag_match_tl  & N138;
  assign \tag_comp_tl_5_.tag_match_tl  = N1411 & N139;
  assign N1411 = ptag_v_i & N1410;
  assign N1410 = ~N1409;
  assign N1409 = N1408 | ptag_i[20];
  assign N1408 = N1407 | ptag_i[21];
  assign N1407 = N1406 | ptag_i[22];
  assign N1406 = N1405 | ptag_i[23];
  assign N1405 = N1404 | ptag_i[24];
  assign N1404 = N1403 | ptag_i[25];
  assign N1403 = ptag_i[27] | ptag_i[26];
  assign load_hit_tl[5] = \tag_comp_tl_5_.tag_match_tl  & N1300;
  assign store_hit_tl[5] = \tag_comp_tl_5_.tag_match_tl  & N148;
  assign \tag_comp_tl_6_.tag_match_tl  = N1420 & N149;
  assign N1420 = ptag_v_i & N1419;
  assign N1419 = ~N1418;
  assign N1418 = N1417 | ptag_i[20];
  assign N1417 = N1416 | ptag_i[21];
  assign N1416 = N1415 | ptag_i[22];
  assign N1415 = N1414 | ptag_i[23];
  assign N1414 = N1413 | ptag_i[24];
  assign N1413 = N1412 | ptag_i[25];
  assign N1412 = ptag_i[27] | ptag_i[26];
  assign load_hit_tl[6] = \tag_comp_tl_6_.tag_match_tl  & N1298;
  assign store_hit_tl[6] = \tag_comp_tl_6_.tag_match_tl  & N158;
  assign \tag_comp_tl_7_.tag_match_tl  = N1429 & N159;
  assign N1429 = ptag_v_i & N1428;
  assign N1428 = ~N1427;
  assign N1427 = N1426 | ptag_i[20];
  assign N1426 = N1425 | ptag_i[21];
  assign N1425 = N1424 | ptag_i[22];
  assign N1424 = N1423 | ptag_i[23];
  assign N1423 = N1422 | ptag_i[24];
  assign N1422 = N1421 | ptag_i[25];
  assign N1421 = ptag_i[27] | ptag_i[26];
  assign load_hit_tl[7] = \tag_comp_tl_7_.tag_match_tl  & N1296;
  assign store_hit_tl[7] = \tag_comp_tl_7_.tag_match_tl  & N168;
  assign uncached_tl = N1430 & N1431;
  assign N1430 = ~decode_tl_r[23];
  assign N1431 = decode_tl_r[17] | ptag_uncached_i;
  assign safe_tv_we = v_tl_r & N1432;
  assign N1432 = ptag_v_i | decode_tl_r[23];
  assign tv_we = safe_tv_we & N1433;
  assign N1433 = ~flush_tv;
  assign _2_net_ = tv_we | critical_recv;
  assign store_miss_tv = N1438 & N1439;
  assign N1438 = N1436 & N1437;
  assign N1436 = N1434 & N1435;
  assign N1434 = decode_tv_r_store_op_ | decode_tv_r_lr_op_;
  assign N1435 = ~store_hit_tv;
  assign N1437 = ~sc_fail_tv;
  assign N1439 = ~nonblocking_req;
  assign load_miss_tv = N1442 & N1439;
  assign N1442 = N1441 & N1437;
  assign N1441 = decode_tv_r_load_op_ & N1440;
  assign N1440 = ~cache_req_o[115];
  assign nonblocking_miss_tv = nonblocking_req & N1443;
  assign N1443 = ~cache_req_yumi_i;
  assign engine_miss_tv = cache_req_v_o & N1444;
  assign N1444 = ~cache_req_yumi_i;
  assign any_miss_tv = N1445 | engine_miss_tv;
  assign N1445 = blocking_miss_tv | nonblocking_miss_tv;
  assign v_o = v_tv_r & N1446;
  assign N1446 = ~any_miss_tv;
  assign N169 = sc_success_tv;
  assign N170 = sc_fail_tv | N169;
  assign N171 = ~N170;
  assign N172 = ~N169;
  assign N173 = sc_fail_tv & N172;
  assign unsigned_o = ~decode_tv_r_signed_op_;
  assign wbuf_v_li = N1451 & N1446;
  assign N1451 = N1449 & N1450;
  assign N1449 = N1448 & N1437;
  assign N1448 = N1447 & store_hit_tv;
  assign N1447 = v_tv_r & decode_tv_r_store_op_;
  assign N1450 = ~uncached_tv_r;
  assign N174 = decode_tv_r_double_op_;
  assign N175 = ~N174;
  assign N176 = decode_tv_r_double_op_;
  assign N177 = ~N176;
  assign N179 = ~N178;
  assign N180 = N178;
  assign N181 = N816 | N817;
  assign N182 = atomic_reg_data[63] & atomic_mem_data[63];
  assign N183 = atomic_reg_data[62] & atomic_mem_data[62];
  assign N184 = atomic_reg_data[61] & atomic_mem_data[61];
  assign N185 = atomic_reg_data[60] & atomic_mem_data[60];
  assign N186 = atomic_reg_data[59] & atomic_mem_data[59];
  assign N187 = atomic_reg_data[58] & atomic_mem_data[58];
  assign N188 = atomic_reg_data[57] & atomic_mem_data[57];
  assign N189 = atomic_reg_data[56] & atomic_mem_data[56];
  assign N190 = atomic_reg_data[55] & atomic_mem_data[55];
  assign N191 = atomic_reg_data[54] & atomic_mem_data[54];
  assign N192 = atomic_reg_data[53] & atomic_mem_data[53];
  assign N193 = atomic_reg_data[52] & atomic_mem_data[52];
  assign N194 = atomic_reg_data[51] & atomic_mem_data[51];
  assign N195 = atomic_reg_data[50] & atomic_mem_data[50];
  assign N196 = atomic_reg_data[49] & atomic_mem_data[49];
  assign N197 = atomic_reg_data[48] & atomic_mem_data[48];
  assign N198 = atomic_reg_data[47] & atomic_mem_data[47];
  assign N199 = atomic_reg_data[46] & atomic_mem_data[46];
  assign N200 = atomic_reg_data[45] & atomic_mem_data[45];
  assign N201 = atomic_reg_data[44] & atomic_mem_data[44];
  assign N202 = atomic_reg_data[43] & atomic_mem_data[43];
  assign N203 = atomic_reg_data[42] & atomic_mem_data[42];
  assign N204 = atomic_reg_data[41] & atomic_mem_data[41];
  assign N205 = atomic_reg_data[40] & atomic_mem_data[40];
  assign N206 = atomic_reg_data[39] & atomic_mem_data[39];
  assign N207 = atomic_reg_data[38] & atomic_mem_data[38];
  assign N208 = atomic_reg_data[37] & atomic_mem_data[37];
  assign N209 = atomic_reg_data[36] & atomic_mem_data[36];
  assign N210 = atomic_reg_data[35] & atomic_mem_data[35];
  assign N211 = atomic_reg_data[34] & atomic_mem_data[34];
  assign N212 = atomic_reg_data[33] & atomic_mem_data[33];
  assign N213 = atomic_reg_data[32] & atomic_mem_data[32];
  assign N214 = atomic_reg_data[31] & atomic_mem_data[31];
  assign N215 = atomic_reg_data[30] & atomic_mem_data[30];
  assign N216 = atomic_reg_data[29] & atomic_mem_data[29];
  assign N217 = atomic_reg_data[28] & atomic_mem_data[28];
  assign N218 = atomic_reg_data[27] & atomic_mem_data[27];
  assign N219 = atomic_reg_data[26] & atomic_mem_data[26];
  assign N220 = atomic_reg_data[25] & atomic_mem_data[25];
  assign N221 = atomic_reg_data[24] & atomic_mem_data[24];
  assign N222 = atomic_reg_data[23] & atomic_mem_data[23];
  assign N223 = atomic_reg_data[22] & atomic_mem_data[22];
  assign N224 = atomic_reg_data[21] & atomic_mem_data[21];
  assign N225 = atomic_reg_data[20] & atomic_mem_data[20];
  assign N226 = atomic_reg_data[19] & atomic_mem_data[19];
  assign N227 = atomic_reg_data[18] & atomic_mem_data[18];
  assign N228 = atomic_reg_data[17] & atomic_mem_data[17];
  assign N229 = atomic_reg_data[16] & atomic_mem_data[16];
  assign N230 = atomic_reg_data[15] & atomic_mem_data[15];
  assign N231 = atomic_reg_data[14] & atomic_mem_data[14];
  assign N232 = atomic_reg_data[13] & atomic_mem_data[13];
  assign N233 = atomic_reg_data[12] & atomic_mem_data[12];
  assign N234 = atomic_reg_data[11] & atomic_mem_data[11];
  assign N235 = atomic_reg_data[10] & atomic_mem_data[10];
  assign N236 = atomic_reg_data[9] & atomic_mem_data[9];
  assign N237 = atomic_reg_data[8] & atomic_mem_data[8];
  assign N238 = atomic_reg_data[7] & atomic_mem_data[7];
  assign N239 = atomic_reg_data[6] & atomic_mem_data[6];
  assign N240 = atomic_reg_data[5] & atomic_mem_data[5];
  assign N241 = atomic_reg_data[4] & atomic_mem_data[4];
  assign N242 = atomic_reg_data[3] & atomic_mem_data[3];
  assign N243 = atomic_reg_data[2] & atomic_mem_data[2];
  assign N244 = atomic_reg_data[1] & atomic_mem_data[1];
  assign N245 = atomic_reg_data[0] & atomic_mem_data[0];
  assign N246 = atomic_reg_data[63] | atomic_mem_data[63];
  assign N247 = atomic_reg_data[62] | atomic_mem_data[62];
  assign N248 = atomic_reg_data[61] | atomic_mem_data[61];
  assign N249 = atomic_reg_data[60] | atomic_mem_data[60];
  assign N250 = atomic_reg_data[59] | atomic_mem_data[59];
  assign N251 = atomic_reg_data[58] | atomic_mem_data[58];
  assign N252 = atomic_reg_data[57] | atomic_mem_data[57];
  assign N253 = atomic_reg_data[56] | atomic_mem_data[56];
  assign N254 = atomic_reg_data[55] | atomic_mem_data[55];
  assign N255 = atomic_reg_data[54] | atomic_mem_data[54];
  assign N256 = atomic_reg_data[53] | atomic_mem_data[53];
  assign N257 = atomic_reg_data[52] | atomic_mem_data[52];
  assign N258 = atomic_reg_data[51] | atomic_mem_data[51];
  assign N259 = atomic_reg_data[50] | atomic_mem_data[50];
  assign N260 = atomic_reg_data[49] | atomic_mem_data[49];
  assign N261 = atomic_reg_data[48] | atomic_mem_data[48];
  assign N262 = atomic_reg_data[47] | atomic_mem_data[47];
  assign N263 = atomic_reg_data[46] | atomic_mem_data[46];
  assign N264 = atomic_reg_data[45] | atomic_mem_data[45];
  assign N265 = atomic_reg_data[44] | atomic_mem_data[44];
  assign N266 = atomic_reg_data[43] | atomic_mem_data[43];
  assign N267 = atomic_reg_data[42] | atomic_mem_data[42];
  assign N268 = atomic_reg_data[41] | atomic_mem_data[41];
  assign N269 = atomic_reg_data[40] | atomic_mem_data[40];
  assign N270 = atomic_reg_data[39] | atomic_mem_data[39];
  assign N271 = atomic_reg_data[38] | atomic_mem_data[38];
  assign N272 = atomic_reg_data[37] | atomic_mem_data[37];
  assign N273 = atomic_reg_data[36] | atomic_mem_data[36];
  assign N274 = atomic_reg_data[35] | atomic_mem_data[35];
  assign N275 = atomic_reg_data[34] | atomic_mem_data[34];
  assign N276 = atomic_reg_data[33] | atomic_mem_data[33];
  assign N277 = atomic_reg_data[32] | atomic_mem_data[32];
  assign N278 = atomic_reg_data[31] | atomic_mem_data[31];
  assign N279 = atomic_reg_data[30] | atomic_mem_data[30];
  assign N280 = atomic_reg_data[29] | atomic_mem_data[29];
  assign N281 = atomic_reg_data[28] | atomic_mem_data[28];
  assign N282 = atomic_reg_data[27] | atomic_mem_data[27];
  assign N283 = atomic_reg_data[26] | atomic_mem_data[26];
  assign N284 = atomic_reg_data[25] | atomic_mem_data[25];
  assign N285 = atomic_reg_data[24] | atomic_mem_data[24];
  assign N286 = atomic_reg_data[23] | atomic_mem_data[23];
  assign N287 = atomic_reg_data[22] | atomic_mem_data[22];
  assign N288 = atomic_reg_data[21] | atomic_mem_data[21];
  assign N289 = atomic_reg_data[20] | atomic_mem_data[20];
  assign N290 = atomic_reg_data[19] | atomic_mem_data[19];
  assign N291 = atomic_reg_data[18] | atomic_mem_data[18];
  assign N292 = atomic_reg_data[17] | atomic_mem_data[17];
  assign N293 = atomic_reg_data[16] | atomic_mem_data[16];
  assign N294 = atomic_reg_data[15] | atomic_mem_data[15];
  assign N295 = atomic_reg_data[14] | atomic_mem_data[14];
  assign N296 = atomic_reg_data[13] | atomic_mem_data[13];
  assign N297 = atomic_reg_data[12] | atomic_mem_data[12];
  assign N298 = atomic_reg_data[11] | atomic_mem_data[11];
  assign N299 = atomic_reg_data[10] | atomic_mem_data[10];
  assign N300 = atomic_reg_data[9] | atomic_mem_data[9];
  assign N301 = atomic_reg_data[8] | atomic_mem_data[8];
  assign N302 = atomic_reg_data[7] | atomic_mem_data[7];
  assign N303 = atomic_reg_data[6] | atomic_mem_data[6];
  assign N304 = atomic_reg_data[5] | atomic_mem_data[5];
  assign N305 = atomic_reg_data[4] | atomic_mem_data[4];
  assign N306 = atomic_reg_data[3] | atomic_mem_data[3];
  assign N307 = atomic_reg_data[2] | atomic_mem_data[2];
  assign N308 = atomic_reg_data[1] | atomic_mem_data[1];
  assign N309 = atomic_reg_data[0] | atomic_mem_data[0];
  assign N310 = atomic_reg_data[63] ^ atomic_mem_data[63];
  assign N311 = atomic_reg_data[62] ^ atomic_mem_data[62];
  assign N312 = atomic_reg_data[61] ^ atomic_mem_data[61];
  assign N313 = atomic_reg_data[60] ^ atomic_mem_data[60];
  assign N314 = atomic_reg_data[59] ^ atomic_mem_data[59];
  assign N315 = atomic_reg_data[58] ^ atomic_mem_data[58];
  assign N316 = atomic_reg_data[57] ^ atomic_mem_data[57];
  assign N317 = atomic_reg_data[56] ^ atomic_mem_data[56];
  assign N318 = atomic_reg_data[55] ^ atomic_mem_data[55];
  assign N319 = atomic_reg_data[54] ^ atomic_mem_data[54];
  assign N320 = atomic_reg_data[53] ^ atomic_mem_data[53];
  assign N321 = atomic_reg_data[52] ^ atomic_mem_data[52];
  assign N322 = atomic_reg_data[51] ^ atomic_mem_data[51];
  assign N323 = atomic_reg_data[50] ^ atomic_mem_data[50];
  assign N324 = atomic_reg_data[49] ^ atomic_mem_data[49];
  assign N325 = atomic_reg_data[48] ^ atomic_mem_data[48];
  assign N326 = atomic_reg_data[47] ^ atomic_mem_data[47];
  assign N327 = atomic_reg_data[46] ^ atomic_mem_data[46];
  assign N328 = atomic_reg_data[45] ^ atomic_mem_data[45];
  assign N329 = atomic_reg_data[44] ^ atomic_mem_data[44];
  assign N330 = atomic_reg_data[43] ^ atomic_mem_data[43];
  assign N331 = atomic_reg_data[42] ^ atomic_mem_data[42];
  assign N332 = atomic_reg_data[41] ^ atomic_mem_data[41];
  assign N333 = atomic_reg_data[40] ^ atomic_mem_data[40];
  assign N334 = atomic_reg_data[39] ^ atomic_mem_data[39];
  assign N335 = atomic_reg_data[38] ^ atomic_mem_data[38];
  assign N336 = atomic_reg_data[37] ^ atomic_mem_data[37];
  assign N337 = atomic_reg_data[36] ^ atomic_mem_data[36];
  assign N338 = atomic_reg_data[35] ^ atomic_mem_data[35];
  assign N339 = atomic_reg_data[34] ^ atomic_mem_data[34];
  assign N340 = atomic_reg_data[33] ^ atomic_mem_data[33];
  assign N341 = atomic_reg_data[32] ^ atomic_mem_data[32];
  assign N342 = atomic_reg_data[31] ^ atomic_mem_data[31];
  assign N343 = atomic_reg_data[30] ^ atomic_mem_data[30];
  assign N344 = atomic_reg_data[29] ^ atomic_mem_data[29];
  assign N345 = atomic_reg_data[28] ^ atomic_mem_data[28];
  assign N346 = atomic_reg_data[27] ^ atomic_mem_data[27];
  assign N347 = atomic_reg_data[26] ^ atomic_mem_data[26];
  assign N348 = atomic_reg_data[25] ^ atomic_mem_data[25];
  assign N349 = atomic_reg_data[24] ^ atomic_mem_data[24];
  assign N350 = atomic_reg_data[23] ^ atomic_mem_data[23];
  assign N351 = atomic_reg_data[22] ^ atomic_mem_data[22];
  assign N352 = atomic_reg_data[21] ^ atomic_mem_data[21];
  assign N353 = atomic_reg_data[20] ^ atomic_mem_data[20];
  assign N354 = atomic_reg_data[19] ^ atomic_mem_data[19];
  assign N355 = atomic_reg_data[18] ^ atomic_mem_data[18];
  assign N356 = atomic_reg_data[17] ^ atomic_mem_data[17];
  assign N357 = atomic_reg_data[16] ^ atomic_mem_data[16];
  assign N358 = atomic_reg_data[15] ^ atomic_mem_data[15];
  assign N359 = atomic_reg_data[14] ^ atomic_mem_data[14];
  assign N360 = atomic_reg_data[13] ^ atomic_mem_data[13];
  assign N361 = atomic_reg_data[12] ^ atomic_mem_data[12];
  assign N362 = atomic_reg_data[11] ^ atomic_mem_data[11];
  assign N363 = atomic_reg_data[10] ^ atomic_mem_data[10];
  assign N364 = atomic_reg_data[9] ^ atomic_mem_data[9];
  assign N365 = atomic_reg_data[8] ^ atomic_mem_data[8];
  assign N366 = atomic_reg_data[7] ^ atomic_mem_data[7];
  assign N367 = atomic_reg_data[6] ^ atomic_mem_data[6];
  assign N368 = atomic_reg_data[5] ^ atomic_mem_data[5];
  assign N369 = atomic_reg_data[4] ^ atomic_mem_data[4];
  assign N370 = atomic_reg_data[3] ^ atomic_mem_data[3];
  assign N371 = atomic_reg_data[2] ^ atomic_mem_data[2];
  assign N372 = atomic_reg_data[1] ^ atomic_mem_data[1];
  assign N373 = atomic_reg_data[0] ^ atomic_mem_data[0];
  assign N439 = ~N438;
  assign N505 = ~N504;
  assign N571 = ~N570;
  assign N637 = ~N636;
  assign N766 = decode_tv_r_amo_op_;
  assign N767 = ~N766;
  assign N768 = ~N782;
  assign wbuf_entry_in_bank_sel__7_ = ld_data_way_select_tv[7] | decode_tv_r_block_op_;
  assign wbuf_entry_in_bank_sel__6_ = ld_data_way_select_tv[6] | decode_tv_r_block_op_;
  assign wbuf_entry_in_bank_sel__5_ = ld_data_way_select_tv[5] | decode_tv_r_block_op_;
  assign wbuf_entry_in_bank_sel__4_ = ld_data_way_select_tv[4] | decode_tv_r_block_op_;
  assign wbuf_entry_in_bank_sel__3_ = ld_data_way_select_tv[3] | decode_tv_r_block_op_;
  assign wbuf_entry_in_bank_sel__2_ = ld_data_way_select_tv[2] | decode_tv_r_block_op_;
  assign wbuf_entry_in_bank_sel__1_ = ld_data_way_select_tv[1] | decode_tv_r_block_op_;
  assign wbuf_entry_in_bank_sel__0_ = ld_data_way_select_tv[0] | decode_tv_r_block_op_;
  assign load_req = N1454 & N1455;
  assign N1454 = N1453 & load_miss_tv;
  assign N1453 = v_tv_r & N1452;
  assign N1452 = ~uncached_tv_r;
  assign N1455 = ~late_o;
  assign store_req = N1458 & N1459;
  assign N1458 = N1457 & store_miss_tv;
  assign N1457 = v_tv_r & N1456;
  assign N1456 = ~uncached_tv_r;
  assign N1459 = ~late_o;
  assign uncached_amo_req = N1462 & N1463;
  assign N1462 = N1461 & ret_o;
  assign N1461 = N1460 & decode_tv_r_amo_op_;
  assign N1460 = v_tv_r & uncached_tv_r;
  assign N1463 = ~late_o;
  assign uncached_load_req = N1467 & N1468;
  assign N1467 = N1466 & decode_tv_r_load_op_;
  assign N1466 = N1464 & N1465;
  assign N1464 = v_tv_r & uncached_tv_r;
  assign N1465 = ~decode_tv_r_amo_op_;
  assign N1468 = ~late_o;
  assign uncached_store_req = N1472 & N1473;
  assign N1472 = N1470 & N1471;
  assign N1470 = N1469 & decode_tv_r_store_op_;
  assign N1469 = v_tv_r & uncached_tv_r;
  assign N1471 = ~ret_o;
  assign N1473 = ~late_o;
  assign bclean_req = N1477 & N1478;
  assign N1477 = N1476 & store_hit_tv;
  assign N1476 = N1475 & decode_tv_r_bclean_op_;
  assign N1475 = v_tv_r & N1474;
  assign N1474 = ~uncached_tv_r;
  assign N1478 = ~late_o;
  assign inval_req = N1483 & N1484;
  assign N1483 = N1481 & N1482;
  assign N1481 = N1480 & decode_tv_r_inval_op_;
  assign N1480 = v_tv_r & N1479;
  assign N1479 = ~uncached_tv_r;
  assign N1482 = ~decode_tv_r_clean_op_;
  assign N1484 = ~late_o;
  assign clean_req = N1489 & N1490;
  assign N1489 = N1487 & N1488;
  assign N1487 = N1486 & decode_tv_r_clean_op_;
  assign N1486 = v_tv_r & N1485;
  assign N1485 = ~uncached_tv_r;
  assign N1488 = ~decode_tv_r_inval_op_;
  assign N1490 = ~late_o;
  assign flush_req = N1494 & N1495;
  assign N1494 = N1493 & decode_tv_r_clean_op_;
  assign N1493 = N1492 & decode_tv_r_inval_op_;
  assign N1492 = v_tv_r & N1491;
  assign N1491 = ~uncached_tv_r;
  assign N1495 = ~late_o;
  assign nonblocking_req = N1496 | N1498;
  assign N1496 = uncached_store_req | 1'b0;
  assign N1498 = N1497 | 1'b0;
  assign N1497 = 1'b0 | bclean_req;
  assign blocking_miss_tv = N1501 | N1503;
  assign N1501 = N1500 | uncached_load_req;
  assign N1500 = N1499 | uncached_amo_req;
  assign N1499 = load_req | store_req;
  assign N1503 = N1502 | flush_req;
  assign N1502 = inval_req | clean_req;
  assign blocking_sent = blocking_miss_tv & cache_req_yumi_i;
  assign cache_req_v_o = N1326 & N1504;
  assign N1504 = blocking_miss_tv | nonblocking_req;
  assign blocking_hazard = cache_req_v_o & blocking_miss_tv;
  assign nonblocking_hazard = nonblocking_req & N1505;
  assign N1505 = ~cache_req_yumi_i;
  assign N769 = N1509 | clean_req;
  assign N1509 = N1508 | inval_req;
  assign N1508 = N1507 | 1'b0;
  assign N1507 = N1506 | bclean_req;
  assign N1506 = load_req | store_req;
  assign N770 = decode_tv_r_block_op_;
  assign N771 = decode_tv_r_double_op_;
  assign N772 = decode_tv_r_word_op_;
  assign N773 = decode_tv_r_half_op_;
  assign N774 = N770 | N769;
  assign N775 = N771 | N774;
  assign N776 = N772 | N775;
  assign N777 = N773 | N776;
  assign N778 = ~N777;
  assign N779 = ~N776;
  assign N780 = ~N774;
  assign N781 = ~decode_tv_r_amo_op_;
  assign N782 = decode_tv_r_amo_op_;
  assign N783 = ~decode_tv_r_amo_subop__0_;
  assign N787 = ~N786;
  assign N788 = ~decode_tv_r_amo_subop__1_;
  assign N791 = ~N790;
  assign N794 = ~N793;
  assign N795 = ~decode_tv_r_amo_subop__2_;
  assign N799 = ~N798;
  assign N801 = ~N800;
  assign N803 = ~N802;
  assign N805 = ~N804;
  assign N806 = ~decode_tv_r_amo_subop__3_;
  assign N809 = ~N808;
  assign N811 = ~N810;
  assign N813 = ~N812;
  assign N815 = ~N814;
  assign N820 = N816 | N819;
  assign N825 = 1'b0;
  assign N826 = 1'b0;
  assign N827 = bclean_req | N825;
  assign N828 = N826 | N827;
  assign N829 = inval_req | N828;
  assign N830 = clean_req | N829;
  assign N831 = flush_req | N830;
  assign N832 = store_req | N831;
  assign N833 = load_req | N832;
  assign N834 = uncached_amo_req | N833;
  assign N835 = uncached_store_req | N834;
  assign N836 = uncached_load_req | N835;
  assign N837 = ~N836;
  assign N838 = ~N835;
  assign N839 = ~N831;
  assign N840 = ~N769;
  assign N841 = N770 & N840;
  assign N842 = ~N770;
  assign N843 = N840 & N842;
  assign N844 = N771 & N843;
  assign N845 = ~N771;
  assign N846 = N843 & N845;
  assign N847 = N772 & N846;
  assign N848 = ~N772;
  assign N849 = N846 & N848;
  assign N850 = N773 & N849;
  assign N851 = ~N825;
  assign N852 = bclean_req & N851;
  assign N853 = ~bclean_req;
  assign N854 = N851 & N853;
  assign N855 = N826 & N854;
  assign N856 = ~N826;
  assign N857 = N854 & N856;
  assign N858 = inval_req & N857;
  assign N859 = ~inval_req;
  assign N860 = N857 & N859;
  assign N861 = clean_req & N860;
  assign N862 = ~clean_req;
  assign N863 = N860 & N862;
  assign N864 = flush_req & N863;
  assign N865 = ~flush_req;
  assign N866 = N863 & N865;
  assign N867 = store_req & N866;
  assign N868 = ~store_req;
  assign N869 = N866 & N868;
  assign N870 = load_req & N869;
  assign N871 = ~load_req;
  assign N872 = N869 & N871;
  assign N873 = uncached_amo_req & N872;
  assign N874 = ~uncached_amo_req;
  assign N875 = N872 & N874;
  assign N876 = uncached_store_req & N875;
  assign N877 = ~uncached_store_req;
  assign N878 = N875 & N877;
  assign N879 = uncached_load_req & N878;
  assign _14_net__7_ = ~metadata_way_v_r[7];
  assign _14_net__6_ = ~metadata_way_v_r[6];
  assign _14_net__5_ = ~metadata_way_v_r[5];
  assign _14_net__4_ = ~metadata_way_v_r[4];
  assign _14_net__3_ = ~metadata_way_v_r[3];
  assign _14_net__2_ = ~metadata_way_v_r[2];
  assign _14_net__1_ = ~metadata_way_v_r[1];
  assign _14_net__0_ = ~metadata_way_v_r[0];
  assign N880 = ~metadata_invalid_exist;
  assign N881 = ~metadata_hit_r;
  assign N882 = ~cache_req_metadata_o[1];
  assign N883 = ~cache_req_metadata_o[2];
  assign N884 = N882 & N883;
  assign N885 = N882 & cache_req_metadata_o[2];
  assign N886 = cache_req_metadata_o[1] & N883;
  assign N887 = cache_req_metadata_o[1] & cache_req_metadata_o[2];
  assign N888 = ~cache_req_metadata_o[3];
  assign N889 = N884 & N888;
  assign N890 = N884 & cache_req_metadata_o[3];
  assign N891 = N886 & N888;
  assign N892 = N886 & cache_req_metadata_o[3];
  assign N893 = N885 & N888;
  assign N894 = N885 & cache_req_metadata_o[3];
  assign N895 = N887 & N888;
  assign N896 = N887 & cache_req_metadata_o[3];
  assign busy_o = cache_req_lock_i | N1511;
  assign N1511 = ~N1510;
  assign N1510 = N1326 | N1329;
  assign ordered_o = N1514 & cache_req_credits_empty_i;
  assign N1514 = N1512 & N1513;
  assign N1512 = ~v_tl_r;
  assign N1513 = ~v_tv_r;
  assign tag_mem_fast_read = safe_tl_we & N1515;
  assign N1515 = ~decode_lo[23];
  assign tag_mem_slow_read = tag_mem_pkt_yumi_o & N1246;
  assign tag_mem_slow_write = tag_mem_pkt_yumi_o & N1249;
  assign tag_mem_fast_write = N1519 | N1522;
  assign N1519 = N1517 & N1518;
  assign N1517 = N1516 & cache_req_o[115];
  assign N1516 = v_tv_r & uncached_tv_r;
  assign N1518 = ~late_o;
  assign N1522 = N1521 & N1518;
  assign N1521 = N1520 & cache_req_o[115];
  assign N1520 = v_tv_r & decode_tv_r_binval_op_;
  assign tag_mem_v_li = N1524 | tag_mem_fast_write;
  assign N1524 = N1523 | tag_mem_slow_write;
  assign N1523 = tag_mem_fast_read | tag_mem_slow_read;
  assign tag_mem_w_li = tag_mem_slow_write | tag_mem_fast_write;
  assign N897 = tag_mem_fast_read | tag_mem_fast_write;
  assign N898 = ~N897;
  assign N899 = ~tag_mem_fast_write;
  assign N900 = tag_mem_fast_read & N899;
  assign tag_mem_pkt_yumi_o = N1530 & N1531;
  assign N1530 = N1528 & N1529;
  assign N1528 = N1526 & N1527;
  assign N1526 = tag_mem_pkt_v_i & N1525;
  assign N1525 = ~N1318;
  assign N1527 = ~tag_mem_fast_read;
  assign N1529 = ~tag_mem_fast_write;
  assign N1531 = ~wbuf_snoop_match_lo;
  assign N901 = ~tag_mem_pkt_i[0];
  assign N905 = ~N904;
  assign N906 = ~tag_mem_pkt_i[1];
  assign N910 = ~N909;
  assign N911 = ~tag_mem_pkt_i[1];
  assign N912 = ~tag_mem_pkt_i[0];
  assign N916 = ~N915;
  assign N918 = ~tag_mem_pkt_i[1];
  assign N919 = ~tag_mem_pkt_i[0];
  assign N922 = N917 | N921;
  assign N923 = ~tag_mem_pkt_i[0];
  assign N927 = ~N926;
  assign N928 = ~tag_mem_pkt_i[1];
  assign N932 = ~N931;
  assign N933 = ~tag_mem_pkt_i[1];
  assign N934 = ~tag_mem_pkt_i[0];
  assign N938 = ~N937;
  assign N940 = ~tag_mem_pkt_i[1];
  assign N941 = ~tag_mem_pkt_i[0];
  assign N944 = N939 | N943;
  assign N945 = ~tag_mem_pkt_i[0];
  assign N949 = ~N948;
  assign N950 = ~tag_mem_pkt_i[1];
  assign N954 = ~N953;
  assign N955 = ~tag_mem_pkt_i[1];
  assign N956 = ~tag_mem_pkt_i[0];
  assign N960 = ~N959;
  assign N962 = ~tag_mem_pkt_i[1];
  assign N963 = ~tag_mem_pkt_i[0];
  assign N966 = N961 | N965;
  assign N967 = ~tag_mem_pkt_i[0];
  assign N971 = ~N970;
  assign N972 = ~tag_mem_pkt_i[1];
  assign N976 = ~N975;
  assign N977 = ~tag_mem_pkt_i[1];
  assign N978 = ~tag_mem_pkt_i[0];
  assign N982 = ~N981;
  assign N984 = ~tag_mem_pkt_i[1];
  assign N985 = ~tag_mem_pkt_i[0];
  assign N988 = N983 | N987;
  assign N989 = ~tag_mem_pkt_i[0];
  assign N993 = ~N992;
  assign N994 = ~tag_mem_pkt_i[1];
  assign N998 = ~N997;
  assign N999 = ~tag_mem_pkt_i[1];
  assign N1000 = ~tag_mem_pkt_i[0];
  assign N1004 = ~N1003;
  assign N1006 = ~tag_mem_pkt_i[1];
  assign N1007 = ~tag_mem_pkt_i[0];
  assign N1010 = N1005 | N1009;
  assign N1011 = ~tag_mem_pkt_i[0];
  assign N1015 = ~N1014;
  assign N1016 = ~tag_mem_pkt_i[1];
  assign N1020 = ~N1019;
  assign N1021 = ~tag_mem_pkt_i[1];
  assign N1022 = ~tag_mem_pkt_i[0];
  assign N1026 = ~N1025;
  assign N1028 = ~tag_mem_pkt_i[1];
  assign N1029 = ~tag_mem_pkt_i[0];
  assign N1032 = N1027 | N1031;
  assign N1033 = ~tag_mem_pkt_i[0];
  assign N1037 = ~N1036;
  assign N1038 = ~tag_mem_pkt_i[1];
  assign N1042 = ~N1041;
  assign N1043 = ~tag_mem_pkt_i[1];
  assign N1044 = ~tag_mem_pkt_i[0];
  assign N1048 = ~N1047;
  assign N1050 = ~tag_mem_pkt_i[1];
  assign N1051 = ~tag_mem_pkt_i[0];
  assign N1054 = N1049 | N1053;
  assign N1055 = ~tag_mem_pkt_i[0];
  assign N1059 = ~N1058;
  assign N1060 = ~tag_mem_pkt_i[1];
  assign N1064 = ~N1063;
  assign N1065 = ~tag_mem_pkt_i[1];
  assign N1066 = ~tag_mem_pkt_i[0];
  assign N1070 = ~N1069;
  assign N1072 = ~tag_mem_pkt_i[1];
  assign N1073 = ~tag_mem_pkt_i[0];
  assign N1076 = N1071 | N1075;
  assign N1077 = ~tag_mem_pkt_way_r[0];
  assign N1078 = ~tag_mem_pkt_way_r[1];
  assign N1079 = N1077 & N1078;
  assign N1080 = N1077 & tag_mem_pkt_way_r[1];
  assign N1081 = tag_mem_pkt_way_r[0] & N1078;
  assign N1082 = tag_mem_pkt_way_r[0] & tag_mem_pkt_way_r[1];
  assign N1083 = ~tag_mem_pkt_way_r[2];
  assign N1084 = N1079 & N1083;
  assign N1085 = N1079 & tag_mem_pkt_way_r[2];
  assign N1086 = N1081 & N1083;
  assign N1087 = N1081 & tag_mem_pkt_way_r[2];
  assign N1088 = N1080 & N1083;
  assign N1089 = N1080 & tag_mem_pkt_way_r[2];
  assign N1090 = N1082 & N1083;
  assign N1091 = N1082 & tag_mem_pkt_way_r[2];
  assign data_mem_fast_read[0] = safe_tl_we & decode_lo[30];
  assign data_mem_force_write[0] = N1532 & wbuf_entry_out_bank_sel__0_;
  assign N1532 = wbuf_v_lo & wbuf_force_lo;
  assign data_mem_slow_write[0] = N1533 & data_mem_write_bank_mask[0];
  assign N1533 = data_mem_pkt_yumi_o & N1254;
  assign data_mem_slow_read[0] = data_mem_pkt_yumi_o & N1252;
  assign data_mem_fast_write[0] = wbuf_yumi_li & wbuf_entry_out_bank_sel__0_;
  assign data_mem_v_li[0] = N1535 | data_mem_slow_write[0];
  assign N1535 = N1534 | data_mem_slow_read[0];
  assign N1534 = data_mem_fast_read[0] | data_mem_fast_write[0];
  assign data_mem_w_li[0] = data_mem_fast_write[0] | data_mem_slow_write[0];
  assign N1092 = ~data_mem_fast_write[0];
  assign N1093 = data_mem_fast_read[0] | data_mem_fast_write[0];
  assign N1094 = ~N1093;
  assign N1095 = data_mem_fast_read[0] & N1092;
  assign data_mem_force_write[1] = N1536 & wbuf_entry_out_bank_sel__1_;
  assign N1536 = wbuf_v_lo & wbuf_force_lo;
  assign data_mem_slow_write[1] = N1537 & data_mem_write_bank_mask[1];
  assign N1537 = data_mem_pkt_yumi_o & N1259;
  assign data_mem_slow_read[1] = data_mem_pkt_yumi_o & N1257;
  assign data_mem_fast_write[1] = wbuf_yumi_li & wbuf_entry_out_bank_sel__1_;
  assign data_mem_v_li[1] = N1539 | data_mem_slow_write[1];
  assign N1539 = N1538 | data_mem_slow_read[1];
  assign N1538 = data_mem_fast_read[0] | data_mem_fast_write[1];
  assign data_mem_w_li[1] = data_mem_fast_write[1] | data_mem_slow_write[1];
  assign N1096 = ~data_mem_fast_write[1];
  assign N1097 = data_mem_fast_read[0] | data_mem_fast_write[1];
  assign N1098 = ~N1097;
  assign N1099 = data_mem_fast_read[0] & N1096;
  assign data_mem_force_write[2] = N1540 & wbuf_entry_out_bank_sel__2_;
  assign N1540 = wbuf_v_lo & wbuf_force_lo;
  assign data_mem_slow_write[2] = N1541 & data_mem_write_bank_mask[2];
  assign N1541 = data_mem_pkt_yumi_o & N1264;
  assign data_mem_slow_read[2] = data_mem_pkt_yumi_o & N1262;
  assign data_mem_fast_write[2] = wbuf_yumi_li & wbuf_entry_out_bank_sel__2_;
  assign data_mem_v_li[2] = N1543 | data_mem_slow_write[2];
  assign N1543 = N1542 | data_mem_slow_read[2];
  assign N1542 = data_mem_fast_read[0] | data_mem_fast_write[2];
  assign data_mem_w_li[2] = data_mem_fast_write[2] | data_mem_slow_write[2];
  assign N1100 = ~data_mem_fast_write[2];
  assign N1101 = data_mem_fast_read[0] | data_mem_fast_write[2];
  assign N1102 = ~N1101;
  assign N1103 = data_mem_fast_read[0] & N1100;
  assign data_mem_force_write[3] = N1544 & wbuf_entry_out_bank_sel__3_;
  assign N1544 = wbuf_v_lo & wbuf_force_lo;
  assign data_mem_slow_write[3] = N1545 & data_mem_write_bank_mask[3];
  assign N1545 = data_mem_pkt_yumi_o & N1269;
  assign data_mem_slow_read[3] = data_mem_pkt_yumi_o & N1267;
  assign data_mem_fast_write[3] = wbuf_yumi_li & wbuf_entry_out_bank_sel__3_;
  assign data_mem_v_li[3] = N1547 | data_mem_slow_write[3];
  assign N1547 = N1546 | data_mem_slow_read[3];
  assign N1546 = data_mem_fast_read[0] | data_mem_fast_write[3];
  assign data_mem_w_li[3] = data_mem_fast_write[3] | data_mem_slow_write[3];
  assign N1104 = ~data_mem_fast_write[3];
  assign N1105 = data_mem_fast_read[0] | data_mem_fast_write[3];
  assign N1106 = ~N1105;
  assign N1107 = data_mem_fast_read[0] & N1104;
  assign data_mem_force_write[4] = N1548 & wbuf_entry_out_bank_sel__4_;
  assign N1548 = wbuf_v_lo & wbuf_force_lo;
  assign data_mem_slow_write[4] = N1549 & data_mem_write_bank_mask[4];
  assign N1549 = data_mem_pkt_yumi_o & N1274;
  assign data_mem_slow_read[4] = data_mem_pkt_yumi_o & N1272;
  assign data_mem_fast_write[4] = wbuf_yumi_li & wbuf_entry_out_bank_sel__4_;
  assign data_mem_v_li[4] = N1551 | data_mem_slow_write[4];
  assign N1551 = N1550 | data_mem_slow_read[4];
  assign N1550 = data_mem_fast_read[0] | data_mem_fast_write[4];
  assign data_mem_w_li[4] = data_mem_fast_write[4] | data_mem_slow_write[4];
  assign N1108 = ~data_mem_fast_write[4];
  assign N1109 = data_mem_fast_read[0] | data_mem_fast_write[4];
  assign N1110 = ~N1109;
  assign N1111 = data_mem_fast_read[0] & N1108;
  assign data_mem_force_write[5] = N1552 & wbuf_entry_out_bank_sel__5_;
  assign N1552 = wbuf_v_lo & wbuf_force_lo;
  assign data_mem_slow_write[5] = N1553 & data_mem_write_bank_mask[5];
  assign N1553 = data_mem_pkt_yumi_o & N1279;
  assign data_mem_slow_read[5] = data_mem_pkt_yumi_o & N1277;
  assign data_mem_fast_write[5] = wbuf_yumi_li & wbuf_entry_out_bank_sel__5_;
  assign data_mem_v_li[5] = N1555 | data_mem_slow_write[5];
  assign N1555 = N1554 | data_mem_slow_read[5];
  assign N1554 = data_mem_fast_read[0] | data_mem_fast_write[5];
  assign data_mem_w_li[5] = data_mem_fast_write[5] | data_mem_slow_write[5];
  assign N1112 = ~data_mem_fast_write[5];
  assign N1113 = data_mem_fast_read[0] | data_mem_fast_write[5];
  assign N1114 = ~N1113;
  assign N1115 = data_mem_fast_read[0] & N1112;
  assign data_mem_force_write[6] = N1556 & wbuf_entry_out_bank_sel__6_;
  assign N1556 = wbuf_v_lo & wbuf_force_lo;
  assign data_mem_slow_write[6] = N1557 & data_mem_write_bank_mask[6];
  assign N1557 = data_mem_pkt_yumi_o & N1284;
  assign data_mem_slow_read[6] = data_mem_pkt_yumi_o & N1282;
  assign data_mem_fast_write[6] = wbuf_yumi_li & wbuf_entry_out_bank_sel__6_;
  assign data_mem_v_li[6] = N1559 | data_mem_slow_write[6];
  assign N1559 = N1558 | data_mem_slow_read[6];
  assign N1558 = data_mem_fast_read[0] | data_mem_fast_write[6];
  assign data_mem_w_li[6] = data_mem_fast_write[6] | data_mem_slow_write[6];
  assign N1116 = ~data_mem_fast_write[6];
  assign N1117 = data_mem_fast_read[0] | data_mem_fast_write[6];
  assign N1118 = ~N1117;
  assign N1119 = data_mem_fast_read[0] & N1116;
  assign data_mem_force_write[7] = N1560 & wbuf_entry_out_bank_sel__7_;
  assign N1560 = wbuf_v_lo & wbuf_force_lo;
  assign data_mem_slow_write[7] = N1561 & data_mem_write_bank_mask[7];
  assign N1561 = data_mem_pkt_yumi_o & N1289;
  assign data_mem_slow_read[7] = data_mem_pkt_yumi_o & N1287;
  assign data_mem_fast_write[7] = wbuf_yumi_li & wbuf_entry_out_bank_sel__7_;
  assign data_mem_v_li[7] = N1563 | data_mem_slow_write[7];
  assign N1563 = N1562 | data_mem_slow_read[7];
  assign N1562 = data_mem_fast_read[0] | data_mem_fast_write[7];
  assign data_mem_w_li[7] = data_mem_fast_write[7] | data_mem_slow_write[7];
  assign N1120 = ~data_mem_fast_write[7];
  assign N1121 = data_mem_fast_read[0] | data_mem_fast_write[7];
  assign N1122 = ~N1121;
  assign N1123 = data_mem_fast_read[0] & N1120;
  assign wbuf_yumi_li = wbuf_v_lo & N1580;
  assign N1580 = N1579 | wbuf_force_lo;
  assign N1579 = ~N1578;
  assign N1578 = N1576 | N1577;
  assign N1576 = N1574 | N1575;
  assign N1574 = N1572 | N1573;
  assign N1572 = N1570 | N1571;
  assign N1570 = N1568 | N1569;
  assign N1568 = N1566 | N1567;
  assign N1566 = N1564 | N1565;
  assign N1564 = data_mem_fast_read[0] & wbuf_entry_out_bank_sel__7_;
  assign N1565 = data_mem_fast_read[0] & wbuf_entry_out_bank_sel__6_;
  assign N1567 = data_mem_fast_read[0] & wbuf_entry_out_bank_sel__5_;
  assign N1569 = data_mem_fast_read[0] & wbuf_entry_out_bank_sel__4_;
  assign N1571 = data_mem_fast_read[0] & wbuf_entry_out_bank_sel__3_;
  assign N1573 = data_mem_fast_read[0] & wbuf_entry_out_bank_sel__2_;
  assign N1575 = data_mem_fast_read[0] & wbuf_entry_out_bank_sel__1_;
  assign N1577 = data_mem_fast_read[0] & wbuf_entry_out_bank_sel__0_;
  assign data_mem_write_hazard = N1593 | N1594;
  assign N1593 = N1591 | N1592;
  assign N1591 = N1589 | N1590;
  assign N1589 = N1587 | N1588;
  assign N1587 = N1585 | N1586;
  assign N1585 = N1583 | N1584;
  assign N1583 = N1581 | N1582;
  assign N1581 = data_mem_fast_read[0] & data_mem_force_write[7];
  assign N1582 = data_mem_fast_read[0] & data_mem_force_write[6];
  assign N1584 = data_mem_fast_read[0] & data_mem_force_write[5];
  assign N1586 = data_mem_fast_read[0] & data_mem_force_write[4];
  assign N1588 = data_mem_fast_read[0] & data_mem_force_write[3];
  assign N1590 = data_mem_fast_read[0] & data_mem_force_write[2];
  assign N1592 = data_mem_fast_read[0] & data_mem_force_write[1];
  assign N1594 = data_mem_fast_read[0] & data_mem_force_write[0];
  assign data_mem_pkt_yumi_o = N1652 & N1531;
  assign N1652 = N1649 & N1651;
  assign N1649 = N1632 & N1648;
  assign N1632 = N1615 & N1631;
  assign N1615 = N1605 & N1614;
  assign N1605 = N1595 & N1604;
  assign N1595 = data_mem_pkt_v_i & N1525;
  assign N1604 = ~N1603;
  assign N1603 = N1602 & N1321;
  assign N1602 = N1601 | data_mem_fast_read[0];
  assign N1601 = N1600 | data_mem_fast_read[0];
  assign N1600 = N1599 | data_mem_fast_read[0];
  assign N1599 = N1598 | data_mem_fast_read[0];
  assign N1598 = N1597 | data_mem_fast_read[0];
  assign N1597 = N1596 | data_mem_fast_read[0];
  assign N1596 = data_mem_fast_read[0] | data_mem_fast_read[0];
  assign N1614 = ~N1613;
  assign N1613 = N1612 & N1324;
  assign N1612 = N1611 | data_mem_fast_write[0];
  assign N1611 = N1610 | data_mem_fast_write[1];
  assign N1610 = N1609 | data_mem_fast_write[2];
  assign N1609 = N1608 | data_mem_fast_write[3];
  assign N1608 = N1607 | data_mem_fast_write[4];
  assign N1607 = N1606 | data_mem_fast_write[5];
  assign N1606 = data_mem_fast_write[7] | data_mem_fast_write[6];
  assign N1631 = ~N1630;
  assign N1630 = N1628 | N1629;
  assign N1628 = N1626 | N1627;
  assign N1626 = N1624 | N1625;
  assign N1624 = N1622 | N1623;
  assign N1622 = N1620 | N1621;
  assign N1620 = N1618 | N1619;
  assign N1618 = N1616 | N1617;
  assign N1616 = data_mem_fast_read[0] & data_mem_write_bank_mask[7];
  assign N1617 = data_mem_fast_read[0] & data_mem_write_bank_mask[6];
  assign N1619 = data_mem_fast_read[0] & data_mem_write_bank_mask[5];
  assign N1621 = data_mem_fast_read[0] & data_mem_write_bank_mask[4];
  assign N1623 = data_mem_fast_read[0] & data_mem_write_bank_mask[3];
  assign N1625 = data_mem_fast_read[0] & data_mem_write_bank_mask[2];
  assign N1627 = data_mem_fast_read[0] & data_mem_write_bank_mask[1];
  assign N1629 = data_mem_fast_read[0] & data_mem_write_bank_mask[0];
  assign N1648 = ~N1647;
  assign N1647 = N1645 | N1646;
  assign N1645 = N1643 | N1644;
  assign N1643 = N1641 | N1642;
  assign N1641 = N1639 | N1640;
  assign N1639 = N1637 | N1638;
  assign N1637 = N1635 | N1636;
  assign N1635 = N1633 | N1634;
  assign N1633 = data_mem_fast_write[7] & data_mem_write_bank_mask[7];
  assign N1634 = data_mem_fast_write[6] & data_mem_write_bank_mask[6];
  assign N1636 = data_mem_fast_write[5] & data_mem_write_bank_mask[5];
  assign N1638 = data_mem_fast_write[4] & data_mem_write_bank_mask[4];
  assign N1640 = data_mem_fast_write[3] & data_mem_write_bank_mask[3];
  assign N1642 = data_mem_fast_write[2] & data_mem_write_bank_mask[2];
  assign N1644 = data_mem_fast_write[1] & data_mem_write_bank_mask[1];
  assign N1646 = data_mem_fast_write[0] & data_mem_write_bank_mask[0];
  assign N1651 = ~N1650;
  assign N1650 = v_tl_r & cache_req_critical_i;
  assign stat_mem_fast_read = N1653 & N1654;
  assign N1653 = v_tv_r & cache_req_yumi_i;
  assign N1654 = ~decode_tv_r_cache_op_;
  assign stat_mem_fast_write = N1659 & N1660;
  assign N1659 = N1657 & N1658;
  assign N1657 = N1655 & N1656;
  assign N1655 = v_tv_r & cache_req_o[115];
  assign N1656 = ~decode_tv_r_cache_op_;
  assign N1658 = ~uncached_tv_r;
  assign N1660 = ~cache_req_yumi_i;
  assign stat_mem_slow_write = stat_mem_pkt_yumi_o & N1294;
  assign stat_mem_slow_read = stat_mem_pkt_yumi_o & N1292;
  assign stat_mem_v_li = N1661 | N1662;
  assign N1661 = stat_mem_fast_read | stat_mem_fast_write;
  assign N1662 = stat_mem_slow_write | stat_mem_slow_read;
  assign stat_mem_w_li = stat_mem_fast_write | stat_mem_slow_write;
  assign N1124 = stat_mem_fast_write | stat_mem_fast_read;
  assign N1125 = ~N1124;
  assign stat_mem_pkt_yumi_o = N1667 & N1669;
  assign N1667 = N1665 & N1666;
  assign N1665 = N1663 & N1664;
  assign N1663 = stat_mem_pkt_v_i & N1525;
  assign N1664 = ~stat_mem_fast_read;
  assign N1666 = ~stat_mem_fast_write;
  assign N1669 = ~N1668;
  assign N1668 = wbuf_snoop_match_lo & N1315;
  assign N1126 = decode_tv_r_store_op_;
  assign N1127 = ~N1126;
  assign \tdm.dirty_mask_v_li  = stat_mem_slow_write | N1670;
  assign N1670 = v_tv_r & decode_tv_r_store_op_;
  assign N1131 = ~stat_mem_pkt_i[0];
  assign N1133 = ~N1132;
  assign N1134 = ~stat_mem_pkt_i[1];
  assign N1135 = stat_mem_pkt_i[1];
  assign \l1_lrsc.set_reservation  = N1671 & store_hit_tv;
  assign N1671 = v_tv_r & decode_tv_r_lr_op_;
  assign \l1_lrsc.clear_reservation  = N1672 | N1675;
  assign N1672 = v_tv_r & decode_tv_r_sc_op_;
  assign N1675 = N1674 & N1145;
  assign N1674 = N1673 & N1144;
  assign N1673 = tag_mem_pkt_yumi_o & \l1_lrsc.load_reserved_v_r ;
  assign \l1_lrsc.load_reservation_match_tv  = N1676 & N1147;
  assign N1676 = \l1_lrsc.load_reserved_v_r  & N1146;
  assign sc_success_tv = N1678 & \l1_lrsc.load_reservation_match_tv ;
  assign N1678 = N1677 & store_hit_tv;
  assign N1677 = v_tv_r & decode_tv_r_sc_op_;
  assign sc_fail_tv = N1679 & N1680;
  assign N1679 = v_tv_r & decode_tv_r_sc_op_;
  assign N1680 = ~sc_success_tv;
  assign \l1_lrsc.lrsc_lock_up  = sc_fail_tv | N1318;
  assign N1148 = N1325 & complete_recv;
  assign N1149 = N1326 & blocking_sent;
  assign N1150 = N1681 & any_miss_tv;
  assign N1681 = N1329 & v_tv_r;
  assign N1151 = N1149 | N1148;
  assign N1152 = N1150 | N1151;
  assign N1153 = ~N1152;
  assign N1155 = decode_tv_r_cache_op_;
  assign N1156 = ~N1148;
  assign N1157 = N1149 & N1156;
  assign N1158 = ~N1149;
  assign N1159 = N1156 & N1158;
  assign N1160 = N1150 & N1159;
  assign \hum.fill_v  = data_mem_pkt_v_i & N1312;
  assign \hum.fill_recv  = N1687 & N1689;
  assign N1687 = N1684 & N1686;
  assign N1684 = \hum.fill_v  & N1683;
  assign N1683 = N1682 | stat_mem_pkt_yumi_o;
  assign N1682 = ~stat_mem_pkt_v_i;
  assign N1686 = N1685 | tag_mem_pkt_yumi_o;
  assign N1685 = ~tag_mem_pkt_v_i;
  assign N1689 = N1688 | data_mem_pkt_yumi_o;
  assign N1688 = ~data_mem_pkt_v_i;
  assign N1161 = ~\hum.fill_v ;
  assign N1162 = \hum.fill_bank_mask_r [7] & N1690;
  assign N1690 = ~data_mem_pkt_fill_mask_expanded[7];
  assign N1163 = \hum.fill_bank_mask_r [6] & N1691;
  assign N1691 = ~data_mem_pkt_fill_mask_expanded[6];
  assign N1164 = \hum.fill_bank_mask_r [5] & N1692;
  assign N1692 = ~data_mem_pkt_fill_mask_expanded[5];
  assign N1165 = \hum.fill_bank_mask_r [4] & N1693;
  assign N1693 = ~data_mem_pkt_fill_mask_expanded[4];
  assign N1166 = \hum.fill_bank_mask_r [3] & N1694;
  assign N1694 = ~data_mem_pkt_fill_mask_expanded[3];
  assign N1167 = \hum.fill_bank_mask_r [2] & N1695;
  assign N1695 = ~data_mem_pkt_fill_mask_expanded[2];
  assign N1168 = \hum.fill_bank_mask_r [1] & N1696;
  assign N1696 = ~data_mem_pkt_fill_mask_expanded[1];
  assign N1169 = \hum.fill_bank_mask_r [0] & N1697;
  assign N1697 = ~data_mem_pkt_fill_mask_expanded[0];
  assign _25_net_ = \hum.fill_recv  | blocking_sent;
  assign fill_hazard = N1715 & N1730;
  assign N1715 = N1699 & N1714;
  assign N1699 = N1698 & N1178;
  assign N1698 = N1325 & v_tl_r;
  assign N1714 = N1712 | N1713;
  assign N1712 = N1710 | N1711;
  assign N1710 = N1708 | N1709;
  assign N1708 = N1706 | N1707;
  assign N1706 = N1704 | N1705;
  assign N1704 = N1702 | N1703;
  assign N1702 = N1700 | N1701;
  assign N1700 = \hum.fill_hit_r [7] & load_hit_tl[7];
  assign N1701 = \hum.fill_hit_r [6] & load_hit_tl[6];
  assign N1703 = \hum.fill_hit_r [5] & load_hit_tl[5];
  assign N1705 = \hum.fill_hit_r [4] & load_hit_tl[4];
  assign N1707 = \hum.fill_hit_r [3] & load_hit_tl[3];
  assign N1709 = \hum.fill_hit_r [2] & load_hit_tl[2];
  assign N1711 = \hum.fill_hit_r [1] & load_hit_tl[1];
  assign N1713 = \hum.fill_hit_r [0] & load_hit_tl[0];
  assign N1730 = N1728 | N1729;
  assign N1728 = N1726 | N1727;
  assign N1726 = N1724 | N1725;
  assign N1724 = N1722 | N1723;
  assign N1722 = N1720 | N1721;
  assign N1720 = N1718 | N1719;
  assign N1718 = N1716 | N1717;
  assign N1716 = \hum.fill_bank_mask_r [7] & bank_sel_one_hot_tl[7];
  assign N1717 = \hum.fill_bank_mask_r [6] & bank_sel_one_hot_tl[6];
  assign N1719 = \hum.fill_bank_mask_r [5] & bank_sel_one_hot_tl[5];
  assign N1721 = \hum.fill_bank_mask_r [4] & bank_sel_one_hot_tl[4];
  assign N1723 = \hum.fill_bank_mask_r [3] & bank_sel_one_hot_tl[3];
  assign N1725 = \hum.fill_bank_mask_r [2] & bank_sel_one_hot_tl[2];
  assign N1727 = \hum.fill_bank_mask_r [1] & bank_sel_one_hot_tl[1];
  assign N1729 = \hum.fill_bank_mask_r [0] & bank_sel_one_hot_tl[0];
  assign pseudo_hit[7] = N1186 | N1194;
  assign pseudo_hit[6] = N1185 | N1193;
  assign pseudo_hit[5] = N1184 | N1192;
  assign pseudo_hit[4] = N1183 | N1191;
  assign pseudo_hit[3] = N1182 | N1190;
  assign pseudo_hit[2] = N1181 | N1189;
  assign pseudo_hit[1] = N1180 | N1188;
  assign pseudo_hit[0] = N1179 | N1187;

  always @(posedge clk_i) begin
    if(reset_i) begin
      state_r_1_sv2v_reg <= 1'b0;
      state_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      state_r_1_sv2v_reg <= state_n[1];
      state_r_0_sv2v_reg <= state_n[0];
    end 
  end


endmodule



module bsg_dff_chain_width_p1_num_stages_p1
(
  clk_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  wire [0:0] data_o;

  bsg_dff_width_p1
  \chained.genblk1_1_.ch_reg 
  (
    .clk_i(clk_i),
    .data_i(data_i[0]),
    .data_o(data_o[0])
  );


endmodule



module bsg_dff_width_p71
(
  clk_i,
  data_i,
  data_o
);

  input [70:0] data_i;
  output [70:0] data_o;
  input clk_i;
  wire [70:0] data_o;
  reg data_o_70_sv2v_reg,data_o_69_sv2v_reg,data_o_68_sv2v_reg,data_o_67_sv2v_reg,
  data_o_66_sv2v_reg,data_o_65_sv2v_reg,data_o_64_sv2v_reg,data_o_63_sv2v_reg,
  data_o_62_sv2v_reg,data_o_61_sv2v_reg,data_o_60_sv2v_reg,data_o_59_sv2v_reg,
  data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,data_o_55_sv2v_reg,
  data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,data_o_51_sv2v_reg,data_o_50_sv2v_reg,
  data_o_49_sv2v_reg,data_o_48_sv2v_reg,data_o_47_sv2v_reg,data_o_46_sv2v_reg,
  data_o_45_sv2v_reg,data_o_44_sv2v_reg,data_o_43_sv2v_reg,data_o_42_sv2v_reg,
  data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,
  data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,
  data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,
  data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,
  data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,
  data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,
  data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,
  data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,
  data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_width_p6
(
  clk_i,
  data_i,
  data_o
);

  input [5:0] data_i;
  output [5:0] data_o;
  input clk_i;
  wire [5:0] data_o;
  reg data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_width_p2
(
  clk_i,
  data_i,
  data_o
);

  input [1:0] data_i;
  output [1:0] data_o;
  input clk_i;
  wire [1:0] data_o;
  reg data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bp_be_pipe_mem_00
(
  clk_i,
  reset_i,
  cfg_bus_i,
  flush_i,
  sfence_i,
  busy_o,
  ordered_o,
  reservation_i,
  rs2_val_i,
  commit_pkt_i,
  tlb_load_miss_v_o,
  tlb_store_miss_v_o,
  cache_miss_v_o,
  cache_replay_v_o,
  load_misaligned_v_o,
  load_access_fault_v_o,
  load_page_fault_v_o,
  store_misaligned_v_o,
  store_access_fault_v_o,
  store_page_fault_v_o,
  early_data_o,
  early_v_o,
  final_data_o,
  final_v_o,
  late_wb_pkt_o,
  late_wb_v_o,
  trans_info_i,
  cache_req_o,
  cache_req_v_o,
  cache_req_yumi_i,
  cache_req_lock_i,
  cache_req_metadata_o,
  cache_req_metadata_v_o,
  cache_req_id_i,
  cache_req_critical_i,
  cache_req_last_i,
  cache_req_credits_full_i,
  cache_req_credits_empty_i,
  data_mem_pkt_v_i,
  data_mem_pkt_i,
  data_mem_pkt_yumi_o,
  data_mem_o,
  tag_mem_pkt_v_i,
  tag_mem_pkt_i,
  tag_mem_pkt_yumi_o,
  tag_mem_o,
  stat_mem_pkt_v_i,
  stat_mem_pkt_i,
  stat_mem_pkt_yumi_o,
  stat_mem_o
);

  input [60:0] cfg_bus_i;
  input [520:0] reservation_i;
  input [63:0] rs2_val_i;
  input [213:0] commit_pkt_i;
  output [65:0] early_data_o;
  output [65:0] final_data_o;
  output [78:0] late_wb_pkt_o;
  input [32:0] trans_info_i;
  output [116:0] cache_req_o;
  output [3:0] cache_req_metadata_o;
  input [0:0] cache_req_id_i;
  input [142:0] data_mem_pkt_i;
  output [511:0] data_mem_o;
  input [34:0] tag_mem_pkt_i;
  output [22:0] tag_mem_o;
  input [10:0] stat_mem_pkt_i;
  output [14:0] stat_mem_o;
  input clk_i;
  input reset_i;
  input flush_i;
  input sfence_i;
  input cache_req_yumi_i;
  input cache_req_lock_i;
  input cache_req_critical_i;
  input cache_req_last_i;
  input cache_req_credits_full_i;
  input cache_req_credits_empty_i;
  input data_mem_pkt_v_i;
  input tag_mem_pkt_v_i;
  input stat_mem_pkt_v_i;
  output busy_o;
  output ordered_o;
  output tlb_load_miss_v_o;
  output tlb_store_miss_v_o;
  output cache_miss_v_o;
  output cache_replay_v_o;
  output load_misaligned_v_o;
  output load_access_fault_v_o;
  output load_page_fault_v_o;
  output store_misaligned_v_o;
  output store_access_fault_v_o;
  output store_page_fault_v_o;
  output early_v_o;
  output final_v_o;
  output late_wb_v_o;
  output cache_req_v_o;
  output cache_req_metadata_v_o;
  output data_mem_pkt_yumi_o;
  output tag_mem_pkt_yumi_o;
  output stat_mem_pkt_yumi_o;
  wire [65:0] early_data_o,final_data_o,dcache_fdata,dcache_data_n;
  wire [78:0] late_wb_pkt_o;
  wire [116:0] cache_req_o;
  wire [3:0] cache_req_metadata_o;
  wire [511:0] data_mem_o;
  wire [22:0] tag_mem_o;
  wire [14:0] stat_mem_o;
  wire busy_o,ordered_o,tlb_load_miss_v_o,tlb_store_miss_v_o,cache_miss_v_o,
  cache_replay_v_o,load_misaligned_v_o,load_access_fault_v_o,load_page_fault_v_o,
  store_misaligned_v_o,store_access_fault_v_o,store_page_fault_v_o,early_v_o,final_v_o,
  late_wb_v_o,cache_req_v_o,cache_req_metadata_v_o,data_mem_pkt_yumi_o,
  tag_mem_pkt_yumi_o,stat_mem_pkt_yumi_o,N0,N1,N2,N3,N4,N5,negedge_clk,is_req,early_v_r,
  dtlb_r_store,dtlb_r_load,dtlb_r_cbo,dtlb_r_ptw,dtlb_r_v,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,
  N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,
  N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,
  N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,
  N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,
  N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,
  N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,
  N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,
  N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,
  N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,
  N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,
  N192,N193,dtlb_v_lo,dtlb_ptag_uncached_lo,dtlb_ptag_dram_lo,frs2_r_v_r,
  dcache_ptag_v,dcache_busy_lo,dcache_ordered_lo,dcache_v,dcache_unsigned,dcache_int,
  dcache_float,dcache_ptw,dcache_ret,dcache_late,early_v_li,N194,N195,dcache_v_r,
  dcache_late_r,dcache_ret_r,final_v_li,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,
  N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,
  N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,
  N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,
  N254,N255,N256,N257,N258,N259,N260,N261,N262,N263;
  wire [63:0] eaddr,dcache_data;
  wire [1:0] dtlb_r_size,dcache_tag;
  wire [27:0] dtlb_ptag_lo;
  wire [4:0] dcache_rd_addr;
  assign late_wb_pkt_o[0] = 1'b0;
  assign late_wb_pkt_o[1] = 1'b0;
  assign late_wb_pkt_o[2] = 1'b0;
  assign late_wb_pkt_o[3] = 1'b0;
  assign late_wb_pkt_o[4] = 1'b0;
  assign late_wb_pkt_o[70] = final_data_o[65];
  assign late_wb_pkt_o[69] = final_data_o[64];
  assign late_wb_pkt_o[68] = final_data_o[63];
  assign late_wb_pkt_o[67] = final_data_o[62];
  assign late_wb_pkt_o[66] = final_data_o[61];
  assign late_wb_pkt_o[65] = final_data_o[60];
  assign late_wb_pkt_o[64] = final_data_o[59];
  assign late_wb_pkt_o[63] = final_data_o[58];
  assign late_wb_pkt_o[62] = final_data_o[57];
  assign late_wb_pkt_o[61] = final_data_o[56];
  assign late_wb_pkt_o[60] = final_data_o[55];
  assign late_wb_pkt_o[59] = final_data_o[54];
  assign late_wb_pkt_o[58] = final_data_o[53];
  assign late_wb_pkt_o[57] = final_data_o[52];
  assign late_wb_pkt_o[56] = final_data_o[51];
  assign late_wb_pkt_o[55] = final_data_o[50];
  assign late_wb_pkt_o[54] = final_data_o[49];
  assign late_wb_pkt_o[53] = final_data_o[48];
  assign late_wb_pkt_o[52] = final_data_o[47];
  assign late_wb_pkt_o[51] = final_data_o[46];
  assign late_wb_pkt_o[50] = final_data_o[45];
  assign late_wb_pkt_o[49] = final_data_o[44];
  assign late_wb_pkt_o[48] = final_data_o[43];
  assign late_wb_pkt_o[47] = final_data_o[42];
  assign late_wb_pkt_o[46] = final_data_o[41];
  assign late_wb_pkt_o[45] = final_data_o[40];
  assign late_wb_pkt_o[44] = final_data_o[39];
  assign late_wb_pkt_o[43] = final_data_o[38];
  assign late_wb_pkt_o[42] = final_data_o[37];
  assign late_wb_pkt_o[41] = final_data_o[36];
  assign late_wb_pkt_o[40] = final_data_o[35];
  assign late_wb_pkt_o[39] = final_data_o[34];
  assign late_wb_pkt_o[38] = final_data_o[33];
  assign late_wb_pkt_o[37] = final_data_o[32];
  assign late_wb_pkt_o[36] = final_data_o[31];
  assign late_wb_pkt_o[35] = final_data_o[30];
  assign late_wb_pkt_o[34] = final_data_o[29];
  assign late_wb_pkt_o[33] = final_data_o[28];
  assign late_wb_pkt_o[32] = final_data_o[27];
  assign late_wb_pkt_o[31] = final_data_o[26];
  assign late_wb_pkt_o[30] = final_data_o[25];
  assign late_wb_pkt_o[29] = final_data_o[24];
  assign late_wb_pkt_o[28] = final_data_o[23];
  assign late_wb_pkt_o[27] = final_data_o[22];
  assign late_wb_pkt_o[26] = final_data_o[21];
  assign late_wb_pkt_o[25] = final_data_o[20];
  assign late_wb_pkt_o[24] = final_data_o[19];
  assign late_wb_pkt_o[23] = final_data_o[18];
  assign late_wb_pkt_o[22] = final_data_o[17];
  assign late_wb_pkt_o[21] = final_data_o[16];
  assign late_wb_pkt_o[20] = final_data_o[15];
  assign late_wb_pkt_o[19] = final_data_o[14];
  assign late_wb_pkt_o[18] = final_data_o[13];
  assign late_wb_pkt_o[17] = final_data_o[12];
  assign late_wb_pkt_o[16] = final_data_o[11];
  assign late_wb_pkt_o[15] = final_data_o[10];
  assign late_wb_pkt_o[14] = final_data_o[9];
  assign late_wb_pkt_o[13] = final_data_o[8];
  assign late_wb_pkt_o[12] = final_data_o[7];
  assign late_wb_pkt_o[11] = final_data_o[6];
  assign late_wb_pkt_o[10] = final_data_o[5];
  assign late_wb_pkt_o[9] = final_data_o[4];
  assign late_wb_pkt_o[8] = final_data_o[3];
  assign late_wb_pkt_o[7] = final_data_o[2];
  assign late_wb_pkt_o[6] = final_data_o[1];
  assign late_wb_pkt_o[5] = final_data_o[0];

  bsg_dff_chain_width_p1_num_stages_p2
  req_chain
  (
    .clk_i(negedge_clk),
    .data_i(is_req),
    .data_o(early_v_r)
  );

  assign N12 = N6 & N7;
  assign N13 = N8 & N9;
  assign N14 = N10 & N11;
  assign N15 = N12 & N13;
  assign N16 = N15 & N14;
  assign N18 = reservation_i[409] | reservation_i[408];
  assign N19 = reservation_i[407] | N17;
  assign N20 = reservation_i[405] | reservation_i[404];
  assign N21 = N18 | N19;
  assign N22 = N21 | N20;
  assign N24 = reservation_i[409] | reservation_i[408];
  assign N25 = N23 | reservation_i[406];
  assign N26 = reservation_i[405] | reservation_i[404];
  assign N27 = N24 | N25;
  assign N28 = N27 | N26;
  assign N31 = reservation_i[409] | reservation_i[408];
  assign N32 = reservation_i[407] | reservation_i[406];
  assign N33 = reservation_i[405] | N30;
  assign N34 = N31 | N32;
  assign N35 = N34 | N33;
  assign N38 = reservation_i[409] | reservation_i[408];
  assign N39 = reservation_i[407] | N36;
  assign N40 = reservation_i[405] | N37;
  assign N41 = N38 | N39;
  assign N42 = N41 | N40;
  assign N45 = reservation_i[409] | reservation_i[408];
  assign N46 = N43 | reservation_i[406];
  assign N47 = reservation_i[405] | N44;
  assign N48 = N45 | N46;
  assign N49 = N48 | N47;
  assign N52 = reservation_i[409] | N51;
  assign N53 = reservation_i[407] | reservation_i[406];
  assign N54 = reservation_i[405] | reservation_i[404];
  assign N55 = N52 | N53;
  assign N56 = N55 | N54;
  assign N59 = reservation_i[409] | N57;
  assign N60 = reservation_i[407] | reservation_i[406];
  assign N61 = reservation_i[405] | N58;
  assign N62 = N59 | N60;
  assign N63 = N62 | N61;
  assign N66 = reservation_i[409] | N64;
  assign N67 = reservation_i[407] | reservation_i[406];
  assign N68 = N65 | reservation_i[404];
  assign N69 = N66 | N67;
  assign N70 = N69 | N68;
  assign N74 = reservation_i[409] | N71;
  assign N75 = reservation_i[407] | reservation_i[406];
  assign N76 = N72 | N73;
  assign N77 = N74 | N75;
  assign N78 = N77 | N76;
  assign N81 = reservation_i[409] | N79;
  assign N82 = reservation_i[407] | N80;
  assign N83 = reservation_i[405] | reservation_i[404];
  assign N84 = N81 | N82;
  assign N85 = N84 | N83;
  assign N89 = reservation_i[409] | N86;
  assign N90 = reservation_i[407] | N87;
  assign N91 = reservation_i[405] | N88;
  assign N92 = N89 | N90;
  assign N93 = N92 | N91;
  assign N97 = reservation_i[409] | N94;
  assign N98 = reservation_i[407] | N95;
  assign N99 = N96 | reservation_i[404];
  assign N100 = N97 | N98;
  assign N101 = N100 | N99;
  assign N106 = reservation_i[409] | N102;
  assign N107 = reservation_i[407] | N103;
  assign N108 = N104 | N105;
  assign N109 = N106 | N107;
  assign N110 = N109 | N108;
  assign N113 = reservation_i[409] | N111;
  assign N114 = N112 | reservation_i[406];
  assign N115 = reservation_i[405] | reservation_i[404];
  assign N116 = N113 | N114;
  assign N117 = N116 | N115;
  assign N119 = reservation_i[409] | reservation_i[408];
  assign N120 = reservation_i[407] | reservation_i[406];
  assign N121 = N118 | reservation_i[404];
  assign N122 = N119 | N120;
  assign N123 = N122 | N121;
  assign N126 = reservation_i[409] | reservation_i[408];
  assign N127 = reservation_i[407] | N124;
  assign N128 = N125 | reservation_i[404];
  assign N129 = N126 | N127;
  assign N130 = N129 | N128;
  assign N133 = reservation_i[409] | reservation_i[408];
  assign N134 = N131 | reservation_i[406];
  assign N135 = N132 | reservation_i[404];
  assign N136 = N133 | N134;
  assign N137 = N136 | N135;
  assign N140 = N138 | reservation_i[408];
  assign N141 = reservation_i[407] | reservation_i[406];
  assign N142 = N139 | reservation_i[404];
  assign N143 = N140 | N141;
  assign N144 = N143 | N142;
  assign N147 = N145 | reservation_i[408];
  assign N148 = reservation_i[407] | N146;
  assign N149 = reservation_i[405] | reservation_i[404];
  assign N150 = N147 | N148;
  assign N151 = N150 | N149;
  assign N155 = reservation_i[409] | reservation_i[408];
  assign N156 = reservation_i[407] | N152;
  assign N157 = N153 | N154;
  assign N158 = N155 | N156;
  assign N159 = N158 | N157;
  assign N162 = reservation_i[409] | reservation_i[408];
  assign N163 = N160 | N161;
  assign N164 = reservation_i[405] | reservation_i[404];
  assign N165 = N162 | N163;
  assign N166 = N165 | N164;
  assign N168 = reservation_i[409] & reservation_i[406];
  assign N169 = N168 & reservation_i[404];
  assign N170 = reservation_i[407] & reservation_i[406];
  assign N171 = N170 & reservation_i[404];
  assign N172 = reservation_i[409] & reservation_i[406];
  assign N173 = N172 & reservation_i[405];
  assign N174 = reservation_i[407] & reservation_i[406];
  assign N175 = N174 & reservation_i[405];
  assign N176 = reservation_i[408] & reservation_i[407];
  assign N177 = N176 & reservation_i[406];
  assign N178 = reservation_i[409] & reservation_i[408];
  assign N179 = reservation_i[408] & reservation_i[407];
  assign N180 = N179 & reservation_i[405];
  assign N183 = N181 & N182;
  assign N184 = reservation_i[405] & reservation_i[404];
  assign N185 = N183 & N184;
  assign N186 = reservation_i[409] & reservation_i[407];
  assign N189 = reservation_i[409] & N187;
  assign N190 = N189 & N188;
  assign N191 = reservation_i[408] & reservation_i[407];
  assign N192 = N191 & reservation_i[404];

  bp_mmu_00_00000008_00000002_00000001_0
  dmmu
  (
    .clk_i(negedge_clk),
    .reset_i(reset_i),
    .flush_i(flush_i),
    .fence_i(sfence_i),
    .priv_mode_i(trans_info_i[32:31]),
    .trans_en_i(trans_info_i[2]),
    .sum_i(trans_info_i[1]),
    .mxr_i(trans_info_i[0]),
    .uncached_mode_i(N197),
    .nonspec_mode_i(N200),
    .hio_mask_i(cfg_bus_i[9:3]),
    .w_v_i(commit_pkt_i[2]),
    .w_vtag_i(commit_pkt_i[127:101]),
    .w_entry_i(commit_pkt_i[56:21]),
    .r_v_i(dtlb_r_v),
    .r_instr_i(1'b0),
    .r_load_i(dtlb_r_load),
    .r_store_i(dtlb_r_store),
    .r_eaddr_i(eaddr),
    .r_size_i(dtlb_r_size),
    .r_cbo_i(dtlb_r_cbo),
    .r_ptw_i(dtlb_r_ptw),
    .r_v_o(dtlb_v_lo),
    .r_ptag_o(dtlb_ptag_lo),
    .r_load_miss_o(tlb_load_miss_v_o),
    .r_store_miss_o(tlb_store_miss_v_o),
    .r_uncached_o(dtlb_ptag_uncached_lo),
    .r_dram_o(dtlb_ptag_dram_lo),
    .r_load_access_fault_o(load_access_fault_v_o),
    .r_store_access_fault_o(store_access_fault_v_o),
    .r_load_misaligned_o(load_misaligned_v_o),
    .r_store_misaligned_o(store_misaligned_v_o),
    .r_load_page_fault_o(load_page_fault_v_o),
    .r_store_page_fault_o(store_page_fault_v_o)
  );


  bsg_dff_width_p1
  freg
  (
    .clk_i(clk_i),
    .data_i(reservation_i[437]),
    .data_o(frs2_r_v_r)
  );


  bp_be_dcache_00
  dcache
  (
    .clk_i(negedge_clk),
    .reset_i(reset_i),
    .cfg_bus_i(cfg_bus_i),
    .busy_o(dcache_busy_lo),
    .ordered_o(dcache_ordered_lo),
    .dcache_pkt_i({ reservation_i[460:456], reservation_i[409:404], eaddr[11:0] }),
    .v_i(is_req),
    .ptag_i(dtlb_ptag_lo),
    .ptag_v_i(dcache_ptag_v),
    .ptag_uncached_i(dtlb_ptag_uncached_lo),
    .ptag_dram_i(dtlb_ptag_dram_lo),
    .st_data_i(rs2_val_i),
    .flush_i(flush_i),
    .v_o(dcache_v),
    .data_o(dcache_data),
    .rd_addr_o(dcache_rd_addr),
    .tag_o(dcache_tag),
    .unsigned_o(dcache_unsigned),
    .int_o(dcache_int),
    .float_o(dcache_float),
    .ptw_o(dcache_ptw),
    .ret_o(dcache_ret),
    .late_o(dcache_late),
    .cache_req_o(cache_req_o),
    .cache_req_v_o(cache_req_v_o),
    .cache_req_yumi_i(cache_req_yumi_i),
    .cache_req_lock_i(cache_req_lock_i),
    .cache_req_metadata_o(cache_req_metadata_o),
    .cache_req_metadata_v_o(cache_req_metadata_v_o),
    .cache_req_id_i(cache_req_id_i[0]),
    .cache_req_critical_i(cache_req_critical_i),
    .cache_req_last_i(cache_req_last_i),
    .cache_req_credits_full_i(cache_req_credits_full_i),
    .cache_req_credits_empty_i(cache_req_credits_empty_i),
    .data_mem_pkt_v_i(data_mem_pkt_v_i),
    .data_mem_pkt_i(data_mem_pkt_i),
    .data_mem_pkt_yumi_o(data_mem_pkt_yumi_o),
    .data_mem_o(data_mem_o),
    .tag_mem_pkt_v_i(tag_mem_pkt_v_i),
    .tag_mem_pkt_i(tag_mem_pkt_i),
    .tag_mem_pkt_yumi_o(tag_mem_pkt_yumi_o),
    .tag_mem_o(tag_mem_o),
    .stat_mem_pkt_v_i(stat_mem_pkt_v_i),
    .stat_mem_pkt_i(stat_mem_pkt_i),
    .stat_mem_pkt_yumi_o(stat_mem_pkt_yumi_o),
    .stat_mem_o(stat_mem_o)
  );


  bsg_dff_chain_width_p1_num_stages_p1
  early_chain
  (
    .clk_i(clk_i),
    .data_i(early_v_li),
    .data_o(early_v_o)
  );


  bp_be_int_box_00
  int_box
  (
    .raw_i(dcache_data),
    .tag_i(dcache_tag),
    .unsigned_i(dcache_unsigned),
    .reg_o(early_data_o)
  );


  bp_be_fp_box_00
  fp_box
  (
    .ieee_i(dcache_data),
    .tag_i(dcache_tag[0]),
    .reg_o(dcache_fdata)
  );


  bsg_dff_width_p71
  data_reg
  (
    .clk_i(negedge_clk),
    .data_i({ dcache_data_n, dcache_rd_addr }),
    .data_o({ final_data_o, late_wb_pkt_o[75:71] })
  );


  bsg_dff_width_p6
  final_reg
  (
    .clk_i(clk_i),
    .data_i({ dcache_v, dcache_int, dcache_float, dcache_ptw, dcache_late, dcache_ret }),
    .data_o({ dcache_v_r, late_wb_pkt_o[78:76], dcache_late_r, dcache_ret_r })
  );


  bsg_dff_chain_width_p1_num_stages_p2
  final_chain
  (
    .clk_i(clk_i),
    .data_i(final_v_li),
    .data_o(final_v_o)
  );


  bsg_dff_width_p2
  sync_reg
  (
    .clk_i(clk_i),
    .data_i({ dcache_ordered_lo, dcache_busy_lo }),
    .data_o({ ordered_o, busy_o })
  );

  assign N196 = cfg_bus_i[12] | cfg_bus_i[13];
  assign N197 = ~N196;
  assign N198 = ~cfg_bus_i[13];
  assign N199 = cfg_bus_i[12] | N198;
  assign N200 = ~N199;
  assign eaddr = reservation_i[388:325] + reservation_i[258:195];
  assign dtlb_r_size = (N0)? { 1'b0, 1'b0 } : 
                       (N1)? { 1'b0, 1'b1 } : 
                       (N2)? { 1'b1, 1'b0 } : 
                       (N3)? { 1'b1, 1'b1 } : 1'b0;
  assign N0 = N29;
  assign N1 = N50;
  assign N2 = N167;
  assign N3 = N193;
  assign dcache_data_n = (N4)? dcache_fdata : 
                         (N5)? early_data_o : 1'b0;
  assign N4 = N195;
  assign N5 = N194;
  assign negedge_clk = ~clk_i;
  assign is_req = reservation_i[520] & N201;
  assign N201 = reservation_i[447] | reservation_i[445];
  assign dtlb_r_store = is_req & N202;
  assign N202 = reservation_i[428] | reservation_i[427];
  assign dtlb_r_load = is_req & reservation_i[429];
  assign dtlb_r_cbo = is_req & reservation_i[427];
  assign dtlb_r_ptw = is_req & reservation_i[426];
  assign dtlb_r_v = N204 | dtlb_r_ptw;
  assign N204 = N203 | dtlb_r_cbo;
  assign N203 = dtlb_r_store | dtlb_r_load;
  assign N6 = ~reservation_i[409];
  assign N7 = ~reservation_i[408];
  assign N8 = ~reservation_i[407];
  assign N9 = ~reservation_i[406];
  assign N10 = ~reservation_i[405];
  assign N11 = ~reservation_i[404];
  assign N17 = ~reservation_i[406];
  assign N23 = ~reservation_i[407];
  assign N29 = N206 | N207;
  assign N206 = N16 | N205;
  assign N205 = ~N22;
  assign N207 = ~N28;
  assign N30 = ~reservation_i[404];
  assign N36 = ~reservation_i[406];
  assign N37 = ~reservation_i[404];
  assign N43 = ~reservation_i[407];
  assign N44 = ~reservation_i[404];
  assign N50 = N210 | N211;
  assign N210 = N208 | N209;
  assign N208 = ~N35;
  assign N209 = ~N42;
  assign N211 = ~N49;
  assign N51 = ~reservation_i[408];
  assign N57 = ~reservation_i[408];
  assign N58 = ~reservation_i[404];
  assign N64 = ~reservation_i[408];
  assign N65 = ~reservation_i[405];
  assign N71 = ~reservation_i[408];
  assign N72 = ~reservation_i[405];
  assign N73 = ~reservation_i[404];
  assign N79 = ~reservation_i[408];
  assign N80 = ~reservation_i[406];
  assign N86 = ~reservation_i[408];
  assign N87 = ~reservation_i[406];
  assign N88 = ~reservation_i[404];
  assign N94 = ~reservation_i[408];
  assign N95 = ~reservation_i[406];
  assign N96 = ~reservation_i[405];
  assign N102 = ~reservation_i[408];
  assign N103 = ~reservation_i[406];
  assign N104 = ~reservation_i[405];
  assign N105 = ~reservation_i[404];
  assign N111 = ~reservation_i[408];
  assign N112 = ~reservation_i[407];
  assign N118 = ~reservation_i[405];
  assign N124 = ~reservation_i[406];
  assign N125 = ~reservation_i[405];
  assign N131 = ~reservation_i[407];
  assign N132 = ~reservation_i[405];
  assign N138 = ~reservation_i[409];
  assign N139 = ~reservation_i[405];
  assign N145 = ~reservation_i[409];
  assign N146 = ~reservation_i[406];
  assign N152 = ~reservation_i[406];
  assign N153 = ~reservation_i[405];
  assign N154 = ~reservation_i[404];
  assign N160 = ~reservation_i[407];
  assign N161 = ~reservation_i[406];
  assign N167 = N240 | N241;
  assign N240 = N238 | N239;
  assign N238 = N236 | N237;
  assign N236 = N234 | N235;
  assign N234 = N232 | N233;
  assign N232 = N230 | N231;
  assign N230 = N228 | N229;
  assign N228 = N226 | N227;
  assign N226 = N224 | N225;
  assign N224 = N222 | N223;
  assign N222 = N220 | N221;
  assign N220 = N218 | N219;
  assign N218 = N216 | N217;
  assign N216 = N214 | N215;
  assign N214 = N212 | N213;
  assign N212 = ~N56;
  assign N213 = ~N63;
  assign N215 = ~N70;
  assign N217 = ~N78;
  assign N219 = ~N85;
  assign N221 = ~N93;
  assign N223 = ~N101;
  assign N225 = ~N110;
  assign N227 = ~N117;
  assign N229 = ~N123;
  assign N231 = ~N130;
  assign N233 = ~N137;
  assign N235 = ~N144;
  assign N237 = ~N151;
  assign N239 = ~N159;
  assign N241 = ~N166;
  assign N181 = ~reservation_i[408];
  assign N182 = ~reservation_i[406];
  assign N187 = ~reservation_i[406];
  assign N188 = ~reservation_i[405];
  assign N193 = N169 | N250;
  assign N250 = N171 | N249;
  assign N249 = N173 | N248;
  assign N248 = N175 | N247;
  assign N247 = N177 | N246;
  assign N246 = N178 | N245;
  assign N245 = N180 | N244;
  assign N244 = N185 | N243;
  assign N243 = N186 | N242;
  assign N242 = N190 | N192;
  assign dcache_ptag_v = N252 & N253;
  assign N252 = dtlb_v_lo & N251;
  assign N251 = ~load_misaligned_v_o;
  assign N253 = ~store_misaligned_v_o;
  assign early_v_li = reservation_i[520] & reservation_i[447];
  assign cache_miss_v_o = N256 & cache_req_yumi_i;
  assign N256 = early_v_r & N255;
  assign N255 = ~N254;
  assign N254 = dcache_v | dcache_late;
  assign cache_replay_v_o = N260 & N261;
  assign N260 = early_v_r & N259;
  assign N259 = ~N258;
  assign N258 = dcache_v & N257;
  assign N257 = ~dcache_late;
  assign N261 = ~cache_req_yumi_i;
  assign N194 = ~dcache_float;
  assign N195 = dcache_float;
  assign final_v_li = reservation_i[520] & reservation_i[445];
  assign late_wb_v_o = N262 & N263;
  assign N262 = dcache_v_r & dcache_ret_r;
  assign N263 = dcache_late_r | late_wb_pkt_o[76];

endmodule



module bsg_dff_chain_width_p4_num_stages_p0
(
  clk_i,
  data_i,
  data_o
);

  input [3:0] data_i;
  output [3:0] data_o;
  input clk_i;
  wire [3:0] data_o;
  assign data_o[3] = data_i[3];
  assign data_o[2] = data_i[2];
  assign data_o[1] = data_i[1];
  assign data_o[0] = data_i[0];

endmodule



module bsg_dff_chain_width_p2_num_stages_p0
(
  clk_i,
  data_i,
  data_o
);

  input [1:0] data_i;
  output [1:0] data_o;
  input clk_i;
  wire [1:0] data_o;
  assign data_o[1] = data_i[1];
  assign data_o[0] = data_i[0];

endmodule



module compressBy4_inWidth54
(
  in,
  out
);

  input [53:0] in;
  output [13:0] out;
  wire [13:0] out;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25;
  assign out[0] = N1 | in[0];
  assign N1 = N0 | in[1];
  assign N0 = in[3] | in[2];
  assign out[1] = N3 | in[4];
  assign N3 = N2 | in[5];
  assign N2 = in[7] | in[6];
  assign out[2] = N5 | in[8];
  assign N5 = N4 | in[9];
  assign N4 = in[11] | in[10];
  assign out[3] = N7 | in[12];
  assign N7 = N6 | in[13];
  assign N6 = in[15] | in[14];
  assign out[4] = N9 | in[16];
  assign N9 = N8 | in[17];
  assign N8 = in[19] | in[18];
  assign out[5] = N11 | in[20];
  assign N11 = N10 | in[21];
  assign N10 = in[23] | in[22];
  assign out[6] = N13 | in[24];
  assign N13 = N12 | in[25];
  assign N12 = in[27] | in[26];
  assign out[7] = N15 | in[28];
  assign N15 = N14 | in[29];
  assign N14 = in[31] | in[30];
  assign out[8] = N17 | in[32];
  assign N17 = N16 | in[33];
  assign N16 = in[35] | in[34];
  assign out[9] = N19 | in[36];
  assign N19 = N18 | in[37];
  assign N18 = in[39] | in[38];
  assign out[10] = N21 | in[40];
  assign N21 = N20 | in[41];
  assign N20 = in[43] | in[42];
  assign out[11] = N23 | in[44];
  assign N23 = N22 | in[45];
  assign N22 = in[47] | in[46];
  assign out[12] = N25 | in[48];
  assign N25 = N24 | in[49];
  assign N24 = in[51] | in[50];
  assign out[13] = in[53] | in[52];

endmodule



module reverse_width13
(
  in,
  out
);

  input [12:0] in;
  output [12:0] out;
  wire [12:0] out;
  assign out[12] = in[0];
  assign out[11] = in[1];
  assign out[10] = in[2];
  assign out[9] = in[3];
  assign out[8] = in[4];
  assign out[7] = in[5];
  assign out[6] = in[6];
  assign out[5] = in[7];
  assign out[4] = in[8];
  assign out[3] = in[9];
  assign out[2] = in[10];
  assign out[1] = in[11];
  assign out[0] = in[12];

endmodule



module lowMaskHiLo_inWidth6_topBound40_bottomBound27
(
  in,
  out
);

  input [5:0] in;
  output [12:0] out;
  wire [12:0] out,reverseOut;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,
  sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,
  sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,sv2v_dc_21,sv2v_dc_22,
  sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,sv2v_dc_27,sv2v_dc_28;

  reverse_width13
  reverse
  (
    .in(reverseOut),
    .out(out)
  );

  assign { sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, reverseOut } = $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) >>> in;

endmodule



module mulAddRecFNToRaw_preMul_expWidth11_sigWidth53_imulEn1
(
  control,
  op,
  a,
  b,
  c,
  roundingMode,
  mulAddA,
  mulAddB,
  mulAddC,
  intermed_compactState,
  intermed_sExp,
  intermed_CDom_CAlignDist,
  intermed_highAlignedSigC
);

  input [0:0] control;
  input [2:0] op;
  input [64:0] a;
  input [64:0] b;
  input [64:0] c;
  input [2:0] roundingMode;
  output [52:0] mulAddA;
  output [52:0] mulAddB;
  output [105:0] mulAddC;
  output [5:0] intermed_compactState;
  output [12:0] intermed_sExp;
  output [5:0] intermed_CDom_CAlignDist;
  output [54:0] intermed_highAlignedSigC;
  wire [52:0] mulAddA,mulAddB;
  wire [105:0] mulAddC;
  wire [5:0] intermed_compactState,intermed_CDom_CAlignDist;
  wire [12:0] intermed_sExp,sExpA,sExpB,sExpC,CExtraMask;
  wire [54:0] intermed_highAlignedSigC;
  wire N0,N1,N2,N3,N4,N5,isNaNA,isInfA,isZeroA,signA,isSigNaNA,isNaNB,isInfB,isZeroB,
  signB,isSigNaNB,isNaNC,isInfC,isZeroC,signC,isSigNaNC,signProd,N6,N7,N8,N9,N10,
  N11,N12,N13,N14,N15,N16,N17,N18,N19,opSignC,N20,isMinCAlign,N21,CIsDominant,N22,
  N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,
  N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,
  N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,
  N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,reduced4CExtra,N96,N97,
  isNaNAOrB,isNaNAny,isInfAOrB,invalidProd,notSigNaN_invalidExc,invalidExc,
  notNaN_addZeros,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,
  N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,
  N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,
  N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,
  N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,
  N178,N179,N180,N181,N182,N183,N184,N185,sv2v_dc_1;
  wire [53:0] sigA,sigB,sigC;
  wire [13:0] sExpAlignedProd,sNatCAlignDist,reduced4SigC;
  wire [7:6] CAlignDist;
  wire [164:110] extComplSigC;
  wire [108:0] mainAlignedSigC;
  wire [0:0] alignedSigC;
  wire [10:0] \fi1.aux_part ;

  recFNToRawFN_expWidth11_sigWidth53
  recFNToRawFN_a
  (
    .in(a),
    .isNaN(isNaNA),
    .isInf(isInfA),
    .isZero(isZeroA),
    .sign(signA),
    .sExp(sExpA),
    .sig(sigA)
  );


  isSigNaNRecFN_expWidth11_sigWidth53
  isSigNaN_a
  (
    .in(a),
    .isSigNaN(isSigNaNA)
  );


  recFNToRawFN_expWidth11_sigWidth53
  recFNToRawFN_b
  (
    .in(b),
    .isNaN(isNaNB),
    .isInf(isInfB),
    .isZero(isZeroB),
    .sign(signB),
    .sExp(sExpB),
    .sig(sigB)
  );


  isSigNaNRecFN_expWidth11_sigWidth53
  isSigNaN_b
  (
    .in(b),
    .isSigNaN(isSigNaNB)
  );


  recFNToRawFN_expWidth11_sigWidth53
  recFNToRawFN_c
  (
    .in(c),
    .isNaN(isNaNC),
    .isInf(isInfC),
    .isZero(isZeroC),
    .sign(signC),
    .sExp(sExpC),
    .sig(sigC)
  );


  isSigNaNRecFN_expWidth11_sigWidth53
  isSigNaN_c
  (
    .in(c),
    .isSigNaN(isSigNaNC)
  );

  assign N20 = $signed(sNatCAlignDist) < $signed(1'b0);
  assign N21 = sNatCAlignDist[12:0] <= { 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1 };
  assign N36 = sNatCAlignDist[12:0] < { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 };
  assign { sv2v_dc_1, intermed_highAlignedSigC, mainAlignedSigC } = $signed({ extComplSigC, extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110], extComplSigC[110:110] }) >>> { CAlignDist, intermed_CDom_CAlignDist };

  compressBy4_inWidth54
  compressBy4_sigC
  (
    .in(sigC),
    .out(reduced4SigC)
  );


  lowMaskHiLo_inWidth6_topBound40_bottomBound27
  lowMask_CExtraMask
  (
    .in({ CAlignDist, intermed_CDom_CAlignDist[5:2] }),
    .out(CExtraMask)
  );

  assign N121 = ~roundingMode[1];
  assign N122 = N121 | roundingMode[2];
  assign N123 = roundingMode[0] | N122;
  assign N124 = ~N123;
  assign { N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99 } = a[10:0] * b[63:53];
  assign { N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110 } = a[63:53] * b[10:0];
  assign { N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6 } = $signed(sExpA) + $signed(sExpB);
  assign \fi1.aux_part  = { N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99 } + { N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110 };
  assign sExpAlignedProd = $signed({ N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6 }) + $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 });
  assign sNatCAlignDist = $signed(sExpAlignedProd) - $signed(sExpC);
  assign { N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23 } = $signed(sExpAlignedProd[12:0]) - $signed({ 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1 });
  assign intermed_sExp = (N0)? sExpC : 
                         (N1)? { N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23 } : 1'b0;
  assign N0 = CIsDominant;
  assign N1 = N22;
  assign { CAlignDist, intermed_CDom_CAlignDist } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                    (N40)? sNatCAlignDist[7:0] : 
                                                    (N38)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 1'b0;
  assign N2 = isMinCAlign;
  assign extComplSigC[164:111] = (N3)? { N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95 } : 
                                 (N4)? sigC : 1'b0;
  assign N3 = extComplSigC[110];
  assign N4 = N41;
  assign alignedSigC[0] = (N3)? N96 : 
                          (N4)? N97 : 1'b0;
  assign mulAddA = (N5)? a[52:0] : 
                   (N98)? sigA[52:0] : 1'b0;
  assign N5 = op[2];
  assign mulAddB = (N5)? b[52:0] : 
                   (N98)? sigB[52:0] : 1'b0;
  assign mulAddC = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \fi1.aux_part , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                   (N98)? mainAlignedSigC[108:3] : 1'b0;
  assign signProd = N125 ^ op[1];
  assign N125 = signA ^ signB;
  assign extComplSigC[110] = N126 ^ op[0];
  assign N126 = signProd ^ signC;
  assign opSignC = signProd ^ extComplSigC[110];
  assign isMinCAlign = N127 | N20;
  assign N127 = isZeroA | isZeroB;
  assign CIsDominant = N128 & N129;
  assign N128 = ~isZeroC;
  assign N129 = isMinCAlign | N21;
  assign N22 = ~CIsDominant;
  assign N37 = N36 | isMinCAlign;
  assign N38 = ~N37;
  assign N39 = ~isMinCAlign;
  assign N40 = N36 & N39;
  assign N41 = ~extComplSigC[110];
  assign N42 = ~sigC[53];
  assign N43 = ~sigC[52];
  assign N44 = ~sigC[51];
  assign N45 = ~sigC[50];
  assign N46 = ~sigC[49];
  assign N47 = ~sigC[48];
  assign N48 = ~sigC[47];
  assign N49 = ~sigC[46];
  assign N50 = ~sigC[45];
  assign N51 = ~sigC[44];
  assign N52 = ~sigC[43];
  assign N53 = ~sigC[42];
  assign N54 = ~sigC[41];
  assign N55 = ~sigC[40];
  assign N56 = ~sigC[39];
  assign N57 = ~sigC[38];
  assign N58 = ~sigC[37];
  assign N59 = ~sigC[36];
  assign N60 = ~sigC[35];
  assign N61 = ~sigC[34];
  assign N62 = ~sigC[33];
  assign N63 = ~sigC[32];
  assign N64 = ~sigC[31];
  assign N65 = ~sigC[30];
  assign N66 = ~sigC[29];
  assign N67 = ~sigC[28];
  assign N68 = ~sigC[27];
  assign N69 = ~sigC[26];
  assign N70 = ~sigC[25];
  assign N71 = ~sigC[24];
  assign N72 = ~sigC[23];
  assign N73 = ~sigC[22];
  assign N74 = ~sigC[21];
  assign N75 = ~sigC[20];
  assign N76 = ~sigC[19];
  assign N77 = ~sigC[18];
  assign N78 = ~sigC[17];
  assign N79 = ~sigC[16];
  assign N80 = ~sigC[15];
  assign N81 = ~sigC[14];
  assign N82 = ~sigC[13];
  assign N83 = ~sigC[12];
  assign N84 = ~sigC[11];
  assign N85 = ~sigC[10];
  assign N86 = ~sigC[9];
  assign N87 = ~sigC[8];
  assign N88 = ~sigC[7];
  assign N89 = ~sigC[6];
  assign N90 = ~sigC[5];
  assign N91 = ~sigC[4];
  assign N92 = ~sigC[3];
  assign N93 = ~sigC[2];
  assign N94 = ~sigC[1];
  assign N95 = ~sigC[0];
  assign reduced4CExtra = N152 | N153;
  assign N152 = N150 | N151;
  assign N150 = N148 | N149;
  assign N148 = N146 | N147;
  assign N146 = N144 | N145;
  assign N144 = N142 | N143;
  assign N142 = N140 | N141;
  assign N140 = N138 | N139;
  assign N138 = N136 | N137;
  assign N136 = N134 | N135;
  assign N134 = N132 | N133;
  assign N132 = N130 | N131;
  assign N130 = reduced4SigC[12] & CExtraMask[12];
  assign N131 = reduced4SigC[11] & CExtraMask[11];
  assign N133 = reduced4SigC[10] & CExtraMask[10];
  assign N135 = reduced4SigC[9] & CExtraMask[9];
  assign N137 = reduced4SigC[8] & CExtraMask[8];
  assign N139 = reduced4SigC[7] & CExtraMask[7];
  assign N141 = reduced4SigC[6] & CExtraMask[6];
  assign N143 = reduced4SigC[5] & CExtraMask[5];
  assign N145 = reduced4SigC[4] & CExtraMask[4];
  assign N147 = reduced4SigC[3] & CExtraMask[3];
  assign N149 = reduced4SigC[2] & CExtraMask[2];
  assign N151 = reduced4SigC[1] & CExtraMask[1];
  assign N153 = reduced4SigC[0] & CExtraMask[0];
  assign N96 = N155 & N156;
  assign N155 = N154 & mainAlignedSigC[0];
  assign N154 = mainAlignedSigC[2] & mainAlignedSigC[1];
  assign N156 = ~reduced4CExtra;
  assign N97 = N158 | reduced4CExtra;
  assign N158 = N157 | mainAlignedSigC[0];
  assign N157 = mainAlignedSigC[2] | mainAlignedSigC[1];
  assign isNaNAOrB = isNaNA | isNaNB;
  assign isNaNAny = isNaNAOrB | isNaNC;
  assign isInfAOrB = isInfA | isInfB;
  assign invalidProd = N159 | N160;
  assign N159 = isInfA & isZeroB;
  assign N160 = isZeroA & isInfB;
  assign notSigNaN_invalidExc = invalidProd | N164;
  assign N164 = N163 & extComplSigC[110];
  assign N163 = N162 & isInfC;
  assign N162 = N161 & isInfAOrB;
  assign N161 = ~isNaNAOrB;
  assign invalidExc = N166 | notSigNaN_invalidExc;
  assign N166 = N165 | isSigNaNC;
  assign N165 = isSigNaNA | isSigNaNB;
  assign notNaN_addZeros = N167 & isZeroC;
  assign N167 = isZeroA | isZeroB;
  assign intermed_compactState[5] = N169 | notNaN_addZeros;
  assign N169 = N168 | isInfC;
  assign N168 = isNaNAny | isInfAOrB;
  assign intermed_compactState[0] = N176 | N179;
  assign N176 = N172 | N175;
  assign N172 = N170 | N171;
  assign N170 = isInfAOrB & signProd;
  assign N171 = isInfC & opSignC;
  assign N175 = N174 & opSignC;
  assign N174 = N173 & signProd;
  assign N173 = notNaN_addZeros & N123;
  assign N179 = N177 & N178;
  assign N177 = notNaN_addZeros & N124;
  assign N178 = signProd | opSignC;
  assign N98 = ~op[2];
  assign intermed_compactState[4] = invalidExc | N181;
  assign N181 = N180 & signProd;
  assign N180 = ~intermed_compactState[5];
  assign intermed_compactState[3] = isNaNAny | N182;
  assign N182 = N180 & extComplSigC[110];
  assign intermed_compactState[2] = N183 | N184;
  assign N183 = isInfAOrB | isInfC;
  assign N184 = N180 & CIsDominant;
  assign intermed_compactState[1] = notNaN_addZeros | N185;
  assign N185 = N180 & alignedSigC[0];

endmodule



module bsg_dff_chain_width_p212_num_stages_p0
(
  clk_i,
  data_i,
  data_o
);

  input [211:0] data_i;
  output [211:0] data_o;
  input clk_i;
  wire [211:0] data_o;
  assign data_o[211] = data_i[211];
  assign data_o[210] = data_i[210];
  assign data_o[209] = data_i[209];
  assign data_o[208] = data_i[208];
  assign data_o[207] = data_i[207];
  assign data_o[206] = data_i[206];
  assign data_o[205] = data_i[205];
  assign data_o[204] = data_i[204];
  assign data_o[203] = data_i[203];
  assign data_o[202] = data_i[202];
  assign data_o[201] = data_i[201];
  assign data_o[200] = data_i[200];
  assign data_o[199] = data_i[199];
  assign data_o[198] = data_i[198];
  assign data_o[197] = data_i[197];
  assign data_o[196] = data_i[196];
  assign data_o[195] = data_i[195];
  assign data_o[194] = data_i[194];
  assign data_o[193] = data_i[193];
  assign data_o[192] = data_i[192];
  assign data_o[191] = data_i[191];
  assign data_o[190] = data_i[190];
  assign data_o[189] = data_i[189];
  assign data_o[188] = data_i[188];
  assign data_o[187] = data_i[187];
  assign data_o[186] = data_i[186];
  assign data_o[185] = data_i[185];
  assign data_o[184] = data_i[184];
  assign data_o[183] = data_i[183];
  assign data_o[182] = data_i[182];
  assign data_o[181] = data_i[181];
  assign data_o[180] = data_i[180];
  assign data_o[179] = data_i[179];
  assign data_o[178] = data_i[178];
  assign data_o[177] = data_i[177];
  assign data_o[176] = data_i[176];
  assign data_o[175] = data_i[175];
  assign data_o[174] = data_i[174];
  assign data_o[173] = data_i[173];
  assign data_o[172] = data_i[172];
  assign data_o[171] = data_i[171];
  assign data_o[170] = data_i[170];
  assign data_o[169] = data_i[169];
  assign data_o[168] = data_i[168];
  assign data_o[167] = data_i[167];
  assign data_o[166] = data_i[166];
  assign data_o[165] = data_i[165];
  assign data_o[164] = data_i[164];
  assign data_o[163] = data_i[163];
  assign data_o[162] = data_i[162];
  assign data_o[161] = data_i[161];
  assign data_o[160] = data_i[160];
  assign data_o[159] = data_i[159];
  assign data_o[158] = data_i[158];
  assign data_o[157] = data_i[157];
  assign data_o[156] = data_i[156];
  assign data_o[155] = data_i[155];
  assign data_o[154] = data_i[154];
  assign data_o[153] = data_i[153];
  assign data_o[152] = data_i[152];
  assign data_o[151] = data_i[151];
  assign data_o[150] = data_i[150];
  assign data_o[149] = data_i[149];
  assign data_o[148] = data_i[148];
  assign data_o[147] = data_i[147];
  assign data_o[146] = data_i[146];
  assign data_o[145] = data_i[145];
  assign data_o[144] = data_i[144];
  assign data_o[143] = data_i[143];
  assign data_o[142] = data_i[142];
  assign data_o[141] = data_i[141];
  assign data_o[140] = data_i[140];
  assign data_o[139] = data_i[139];
  assign data_o[138] = data_i[138];
  assign data_o[137] = data_i[137];
  assign data_o[136] = data_i[136];
  assign data_o[135] = data_i[135];
  assign data_o[134] = data_i[134];
  assign data_o[133] = data_i[133];
  assign data_o[132] = data_i[132];
  assign data_o[131] = data_i[131];
  assign data_o[130] = data_i[130];
  assign data_o[129] = data_i[129];
  assign data_o[128] = data_i[128];
  assign data_o[127] = data_i[127];
  assign data_o[126] = data_i[126];
  assign data_o[125] = data_i[125];
  assign data_o[124] = data_i[124];
  assign data_o[123] = data_i[123];
  assign data_o[122] = data_i[122];
  assign data_o[121] = data_i[121];
  assign data_o[120] = data_i[120];
  assign data_o[119] = data_i[119];
  assign data_o[118] = data_i[118];
  assign data_o[117] = data_i[117];
  assign data_o[116] = data_i[116];
  assign data_o[115] = data_i[115];
  assign data_o[114] = data_i[114];
  assign data_o[113] = data_i[113];
  assign data_o[112] = data_i[112];
  assign data_o[111] = data_i[111];
  assign data_o[110] = data_i[110];
  assign data_o[109] = data_i[109];
  assign data_o[108] = data_i[108];
  assign data_o[107] = data_i[107];
  assign data_o[106] = data_i[106];
  assign data_o[105] = data_i[105];
  assign data_o[104] = data_i[104];
  assign data_o[103] = data_i[103];
  assign data_o[102] = data_i[102];
  assign data_o[101] = data_i[101];
  assign data_o[100] = data_i[100];
  assign data_o[99] = data_i[99];
  assign data_o[98] = data_i[98];
  assign data_o[97] = data_i[97];
  assign data_o[96] = data_i[96];
  assign data_o[95] = data_i[95];
  assign data_o[94] = data_i[94];
  assign data_o[93] = data_i[93];
  assign data_o[92] = data_i[92];
  assign data_o[91] = data_i[91];
  assign data_o[90] = data_i[90];
  assign data_o[89] = data_i[89];
  assign data_o[88] = data_i[88];
  assign data_o[87] = data_i[87];
  assign data_o[86] = data_i[86];
  assign data_o[85] = data_i[85];
  assign data_o[84] = data_i[84];
  assign data_o[83] = data_i[83];
  assign data_o[82] = data_i[82];
  assign data_o[81] = data_i[81];
  assign data_o[80] = data_i[80];
  assign data_o[79] = data_i[79];
  assign data_o[78] = data_i[78];
  assign data_o[77] = data_i[77];
  assign data_o[76] = data_i[76];
  assign data_o[75] = data_i[75];
  assign data_o[74] = data_i[74];
  assign data_o[73] = data_i[73];
  assign data_o[72] = data_i[72];
  assign data_o[71] = data_i[71];
  assign data_o[70] = data_i[70];
  assign data_o[69] = data_i[69];
  assign data_o[68] = data_i[68];
  assign data_o[67] = data_i[67];
  assign data_o[66] = data_i[66];
  assign data_o[65] = data_i[65];
  assign data_o[64] = data_i[64];
  assign data_o[63] = data_i[63];
  assign data_o[62] = data_i[62];
  assign data_o[61] = data_i[61];
  assign data_o[60] = data_i[60];
  assign data_o[59] = data_i[59];
  assign data_o[58] = data_i[58];
  assign data_o[57] = data_i[57];
  assign data_o[56] = data_i[56];
  assign data_o[55] = data_i[55];
  assign data_o[54] = data_i[54];
  assign data_o[53] = data_i[53];
  assign data_o[52] = data_i[52];
  assign data_o[51] = data_i[51];
  assign data_o[50] = data_i[50];
  assign data_o[49] = data_i[49];
  assign data_o[48] = data_i[48];
  assign data_o[47] = data_i[47];
  assign data_o[46] = data_i[46];
  assign data_o[45] = data_i[45];
  assign data_o[44] = data_i[44];
  assign data_o[43] = data_i[43];
  assign data_o[42] = data_i[42];
  assign data_o[41] = data_i[41];
  assign data_o[40] = data_i[40];
  assign data_o[39] = data_i[39];
  assign data_o[38] = data_i[38];
  assign data_o[37] = data_i[37];
  assign data_o[36] = data_i[36];
  assign data_o[35] = data_i[35];
  assign data_o[34] = data_i[34];
  assign data_o[33] = data_i[33];
  assign data_o[32] = data_i[32];
  assign data_o[31] = data_i[31];
  assign data_o[30] = data_i[30];
  assign data_o[29] = data_i[29];
  assign data_o[28] = data_i[28];
  assign data_o[27] = data_i[27];
  assign data_o[26] = data_i[26];
  assign data_o[25] = data_i[25];
  assign data_o[24] = data_i[24];
  assign data_o[23] = data_i[23];
  assign data_o[22] = data_i[22];
  assign data_o[21] = data_i[21];
  assign data_o[20] = data_i[20];
  assign data_o[19] = data_i[19];
  assign data_o[18] = data_i[18];
  assign data_o[17] = data_i[17];
  assign data_o[16] = data_i[16];
  assign data_o[15] = data_i[15];
  assign data_o[14] = data_i[14];
  assign data_o[13] = data_i[13];
  assign data_o[12] = data_i[12];
  assign data_o[11] = data_i[11];
  assign data_o[10] = data_i[10];
  assign data_o[9] = data_i[9];
  assign data_o[8] = data_i[8];
  assign data_o[7] = data_i[7];
  assign data_o[6] = data_i[6];
  assign data_o[5] = data_i[5];
  assign data_o[4] = data_i[4];
  assign data_o[3] = data_i[3];
  assign data_o[2] = data_i[2];
  assign data_o[1] = data_i[1];
  assign data_o[0] = data_i[0];

endmodule



module bsg_dff_chain_width_p107_num_stages_p0
(
  clk_i,
  data_i,
  data_o
);

  input [106:0] data_i;
  output [106:0] data_o;
  input clk_i;
  wire [106:0] data_o;
  assign data_o[106] = data_i[106];
  assign data_o[105] = data_i[105];
  assign data_o[104] = data_i[104];
  assign data_o[103] = data_i[103];
  assign data_o[102] = data_i[102];
  assign data_o[101] = data_i[101];
  assign data_o[100] = data_i[100];
  assign data_o[99] = data_i[99];
  assign data_o[98] = data_i[98];
  assign data_o[97] = data_i[97];
  assign data_o[96] = data_i[96];
  assign data_o[95] = data_i[95];
  assign data_o[94] = data_i[94];
  assign data_o[93] = data_i[93];
  assign data_o[92] = data_i[92];
  assign data_o[91] = data_i[91];
  assign data_o[90] = data_i[90];
  assign data_o[89] = data_i[89];
  assign data_o[88] = data_i[88];
  assign data_o[87] = data_i[87];
  assign data_o[86] = data_i[86];
  assign data_o[85] = data_i[85];
  assign data_o[84] = data_i[84];
  assign data_o[83] = data_i[83];
  assign data_o[82] = data_i[82];
  assign data_o[81] = data_i[81];
  assign data_o[80] = data_i[80];
  assign data_o[79] = data_i[79];
  assign data_o[78] = data_i[78];
  assign data_o[77] = data_i[77];
  assign data_o[76] = data_i[76];
  assign data_o[75] = data_i[75];
  assign data_o[74] = data_i[74];
  assign data_o[73] = data_i[73];
  assign data_o[72] = data_i[72];
  assign data_o[71] = data_i[71];
  assign data_o[70] = data_i[70];
  assign data_o[69] = data_i[69];
  assign data_o[68] = data_i[68];
  assign data_o[67] = data_i[67];
  assign data_o[66] = data_i[66];
  assign data_o[65] = data_i[65];
  assign data_o[64] = data_i[64];
  assign data_o[63] = data_i[63];
  assign data_o[62] = data_i[62];
  assign data_o[61] = data_i[61];
  assign data_o[60] = data_i[60];
  assign data_o[59] = data_i[59];
  assign data_o[58] = data_i[58];
  assign data_o[57] = data_i[57];
  assign data_o[56] = data_i[56];
  assign data_o[55] = data_i[55];
  assign data_o[54] = data_i[54];
  assign data_o[53] = data_i[53];
  assign data_o[52] = data_i[52];
  assign data_o[51] = data_i[51];
  assign data_o[50] = data_i[50];
  assign data_o[49] = data_i[49];
  assign data_o[48] = data_i[48];
  assign data_o[47] = data_i[47];
  assign data_o[46] = data_i[46];
  assign data_o[45] = data_i[45];
  assign data_o[44] = data_i[44];
  assign data_o[43] = data_i[43];
  assign data_o[42] = data_i[42];
  assign data_o[41] = data_i[41];
  assign data_o[40] = data_i[40];
  assign data_o[39] = data_i[39];
  assign data_o[38] = data_i[38];
  assign data_o[37] = data_i[37];
  assign data_o[36] = data_i[36];
  assign data_o[35] = data_i[35];
  assign data_o[34] = data_i[34];
  assign data_o[33] = data_i[33];
  assign data_o[32] = data_i[32];
  assign data_o[31] = data_i[31];
  assign data_o[30] = data_i[30];
  assign data_o[29] = data_i[29];
  assign data_o[28] = data_i[28];
  assign data_o[27] = data_i[27];
  assign data_o[26] = data_i[26];
  assign data_o[25] = data_i[25];
  assign data_o[24] = data_i[24];
  assign data_o[23] = data_i[23];
  assign data_o[22] = data_i[22];
  assign data_o[21] = data_i[21];
  assign data_o[20] = data_i[20];
  assign data_o[19] = data_i[19];
  assign data_o[18] = data_i[18];
  assign data_o[17] = data_i[17];
  assign data_o[16] = data_i[16];
  assign data_o[15] = data_i[15];
  assign data_o[14] = data_i[14];
  assign data_o[13] = data_i[13];
  assign data_o[12] = data_i[12];
  assign data_o[11] = data_i[11];
  assign data_o[10] = data_i[10];
  assign data_o[9] = data_i[9];
  assign data_o[8] = data_i[8];
  assign data_o[7] = data_i[7];
  assign data_o[6] = data_i[6];
  assign data_o[5] = data_i[5];
  assign data_o[4] = data_i[4];
  assign data_o[3] = data_i[3];
  assign data_o[2] = data_i[2];
  assign data_o[1] = data_i[1];
  assign data_o[0] = data_i[0];

endmodule



module bsg_mul_add_unsigned_width_a_p53_width_b_p53_width_c_p106_width_o_p107_pipeline_p0
(
  clk_i,
  a_i,
  b_i,
  c_i,
  o
);

  input [52:0] a_i;
  input [52:0] b_i;
  input [105:0] c_i;
  output [106:0] o;
  input clk_i;
  wire [106:0] o,o_r;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105;
  wire [52:0] a_r,b_r;
  wire [105:0] c_r;

  bsg_dff_chain_width_p212_num_stages_p0
  pre_mul_add
  (
    .clk_i(clk_i),
    .data_i({ a_i, b_i, c_i }),
    .data_o({ a_r, b_r, c_r })
  );


  bsg_dff_chain_width_p107_num_stages_p0
  post_mul_add
  (
    .clk_i(clk_i),
    .data_i(o_r),
    .data_o(o)
  );

  assign { N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0 } = a_r * b_r;
  assign o_r = { N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0 } + c_r;

endmodule



module bsg_dff_chain_width_p83_num_stages_p0
(
  clk_i,
  data_i,
  data_o
);

  input [82:0] data_i;
  output [82:0] data_o;
  input clk_i;
  wire [82:0] data_o;
  assign data_o[82] = data_i[82];
  assign data_o[81] = data_i[81];
  assign data_o[80] = data_i[80];
  assign data_o[79] = data_i[79];
  assign data_o[78] = data_i[78];
  assign data_o[77] = data_i[77];
  assign data_o[76] = data_i[76];
  assign data_o[75] = data_i[75];
  assign data_o[74] = data_i[74];
  assign data_o[73] = data_i[73];
  assign data_o[72] = data_i[72];
  assign data_o[71] = data_i[71];
  assign data_o[70] = data_i[70];
  assign data_o[69] = data_i[69];
  assign data_o[68] = data_i[68];
  assign data_o[67] = data_i[67];
  assign data_o[66] = data_i[66];
  assign data_o[65] = data_i[65];
  assign data_o[64] = data_i[64];
  assign data_o[63] = data_i[63];
  assign data_o[62] = data_i[62];
  assign data_o[61] = data_i[61];
  assign data_o[60] = data_i[60];
  assign data_o[59] = data_i[59];
  assign data_o[58] = data_i[58];
  assign data_o[57] = data_i[57];
  assign data_o[56] = data_i[56];
  assign data_o[55] = data_i[55];
  assign data_o[54] = data_i[54];
  assign data_o[53] = data_i[53];
  assign data_o[52] = data_i[52];
  assign data_o[51] = data_i[51];
  assign data_o[50] = data_i[50];
  assign data_o[49] = data_i[49];
  assign data_o[48] = data_i[48];
  assign data_o[47] = data_i[47];
  assign data_o[46] = data_i[46];
  assign data_o[45] = data_i[45];
  assign data_o[44] = data_i[44];
  assign data_o[43] = data_i[43];
  assign data_o[42] = data_i[42];
  assign data_o[41] = data_i[41];
  assign data_o[40] = data_i[40];
  assign data_o[39] = data_i[39];
  assign data_o[38] = data_i[38];
  assign data_o[37] = data_i[37];
  assign data_o[36] = data_i[36];
  assign data_o[35] = data_i[35];
  assign data_o[34] = data_i[34];
  assign data_o[33] = data_i[33];
  assign data_o[32] = data_i[32];
  assign data_o[31] = data_i[31];
  assign data_o[30] = data_i[30];
  assign data_o[29] = data_i[29];
  assign data_o[28] = data_i[28];
  assign data_o[27] = data_i[27];
  assign data_o[26] = data_i[26];
  assign data_o[25] = data_i[25];
  assign data_o[24] = data_i[24];
  assign data_o[23] = data_i[23];
  assign data_o[22] = data_i[22];
  assign data_o[21] = data_i[21];
  assign data_o[20] = data_i[20];
  assign data_o[19] = data_i[19];
  assign data_o[18] = data_i[18];
  assign data_o[17] = data_i[17];
  assign data_o[16] = data_i[16];
  assign data_o[15] = data_i[15];
  assign data_o[14] = data_i[14];
  assign data_o[13] = data_i[13];
  assign data_o[12] = data_i[12];
  assign data_o[11] = data_i[11];
  assign data_o[10] = data_i[10];
  assign data_o[9] = data_i[9];
  assign data_o[8] = data_i[8];
  assign data_o[7] = data_i[7];
  assign data_o[6] = data_i[6];
  assign data_o[5] = data_i[5];
  assign data_o[4] = data_i[4];
  assign data_o[3] = data_i[3];
  assign data_o[2] = data_i[2];
  assign data_o[1] = data_i[1];
  assign data_o[0] = data_i[0];

endmodule



module compressBy4_inWidth55
(
  in,
  out
);

  input [54:0] in;
  output [13:0] out;
  wire [13:0] out;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26;
  assign out[0] = N1 | in[0];
  assign N1 = N0 | in[1];
  assign N0 = in[3] | in[2];
  assign out[1] = N3 | in[4];
  assign N3 = N2 | in[5];
  assign N2 = in[7] | in[6];
  assign out[2] = N5 | in[8];
  assign N5 = N4 | in[9];
  assign N4 = in[11] | in[10];
  assign out[3] = N7 | in[12];
  assign N7 = N6 | in[13];
  assign N6 = in[15] | in[14];
  assign out[4] = N9 | in[16];
  assign N9 = N8 | in[17];
  assign N8 = in[19] | in[18];
  assign out[5] = N11 | in[20];
  assign N11 = N10 | in[21];
  assign N10 = in[23] | in[22];
  assign out[6] = N13 | in[24];
  assign N13 = N12 | in[25];
  assign N12 = in[27] | in[26];
  assign out[7] = N15 | in[28];
  assign N15 = N14 | in[29];
  assign N14 = in[31] | in[30];
  assign out[8] = N17 | in[32];
  assign N17 = N16 | in[33];
  assign N16 = in[35] | in[34];
  assign out[9] = N19 | in[36];
  assign N19 = N18 | in[37];
  assign N18 = in[39] | in[38];
  assign out[10] = N21 | in[40];
  assign N21 = N20 | in[41];
  assign N20 = in[43] | in[42];
  assign out[11] = N23 | in[44];
  assign N23 = N22 | in[45];
  assign N22 = in[47] | in[46];
  assign out[12] = N25 | in[48];
  assign N25 = N24 | in[49];
  assign N24 = in[51] | in[50];
  assign out[13] = N26 | in[52];
  assign N26 = in[54] | in[53];

endmodule



module lowMaskLoHi_inWidth4_topBound0_bottomBound13
(
  in,
  out
);

  input [3:0] in;
  output [12:0] out;
  wire [12:0] out,reverseOut;
  wire N0,N1,N2,N3,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3;

  reverse_width13
  reverse
  (
    .in(reverseOut),
    .out(out)
  );

  assign { sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, reverseOut } = $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) >>> { N0, N1, N2, N3 };
  assign N0 = ~in[3];
  assign N1 = ~in[2];
  assign N2 = ~in[1];
  assign N3 = ~in[0];

endmodule



module compressBy2_inWidth109
(
  in,
  out
);

  input [108:0] in;
  output [54:0] out;
  wire [54:0] out;
  wire out_54_;
  assign out_54_ = in[108];
  assign out[54] = out_54_;
  assign out[0] = in[1] | in[0];
  assign out[1] = in[3] | in[2];
  assign out[2] = in[5] | in[4];
  assign out[3] = in[7] | in[6];
  assign out[4] = in[9] | in[8];
  assign out[5] = in[11] | in[10];
  assign out[6] = in[13] | in[12];
  assign out[7] = in[15] | in[14];
  assign out[8] = in[17] | in[16];
  assign out[9] = in[19] | in[18];
  assign out[10] = in[21] | in[20];
  assign out[11] = in[23] | in[22];
  assign out[12] = in[25] | in[24];
  assign out[13] = in[27] | in[26];
  assign out[14] = in[29] | in[28];
  assign out[15] = in[31] | in[30];
  assign out[16] = in[33] | in[32];
  assign out[17] = in[35] | in[34];
  assign out[18] = in[37] | in[36];
  assign out[19] = in[39] | in[38];
  assign out[20] = in[41] | in[40];
  assign out[21] = in[43] | in[42];
  assign out[22] = in[45] | in[44];
  assign out[23] = in[47] | in[46];
  assign out[24] = in[49] | in[48];
  assign out[25] = in[51] | in[50];
  assign out[26] = in[53] | in[52];
  assign out[27] = in[55] | in[54];
  assign out[28] = in[57] | in[56];
  assign out[29] = in[59] | in[58];
  assign out[30] = in[61] | in[60];
  assign out[31] = in[63] | in[62];
  assign out[32] = in[65] | in[64];
  assign out[33] = in[67] | in[66];
  assign out[34] = in[69] | in[68];
  assign out[35] = in[71] | in[70];
  assign out[36] = in[73] | in[72];
  assign out[37] = in[75] | in[74];
  assign out[38] = in[77] | in[76];
  assign out[39] = in[79] | in[78];
  assign out[40] = in[81] | in[80];
  assign out[41] = in[83] | in[82];
  assign out[42] = in[85] | in[84];
  assign out[43] = in[87] | in[86];
  assign out[44] = in[89] | in[88];
  assign out[45] = in[91] | in[90];
  assign out[46] = in[93] | in[92];
  assign out[47] = in[95] | in[94];
  assign out[48] = in[97] | in[96];
  assign out[49] = in[99] | in[98];
  assign out[50] = in[101] | in[100];
  assign out[51] = in[103] | in[102];
  assign out[52] = in[105] | in[104];
  assign out[53] = in[107] | in[106];

endmodule



module bsg_scan_width_p56_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [55:0] i;
  output [55:0] o;
  wire [55:0] o;
  wire t_5__55_,t_5__54_,t_5__53_,t_5__52_,t_5__51_,t_5__50_,t_5__49_,t_5__48_,
  t_5__47_,t_5__46_,t_5__45_,t_5__44_,t_5__43_,t_5__42_,t_5__41_,t_5__40_,t_5__39_,
  t_5__38_,t_5__37_,t_5__36_,t_5__35_,t_5__34_,t_5__33_,t_5__32_,t_5__31_,t_5__30_,
  t_5__29_,t_5__28_,t_5__27_,t_5__26_,t_5__25_,t_5__24_,t_5__23_,t_5__22_,t_5__21_,
  t_5__20_,t_5__19_,t_5__18_,t_5__17_,t_5__16_,t_5__15_,t_5__14_,t_5__13_,t_5__12_,
  t_5__11_,t_5__10_,t_5__9_,t_5__8_,t_5__7_,t_5__6_,t_5__5_,t_5__4_,t_5__3_,t_5__2_,
  t_5__1_,t_5__0_,t_4__55_,t_4__54_,t_4__53_,t_4__52_,t_4__51_,t_4__50_,t_4__49_,
  t_4__48_,t_4__47_,t_4__46_,t_4__45_,t_4__44_,t_4__43_,t_4__42_,t_4__41_,t_4__40_,
  t_4__39_,t_4__38_,t_4__37_,t_4__36_,t_4__35_,t_4__34_,t_4__33_,t_4__32_,t_4__31_,
  t_4__30_,t_4__29_,t_4__28_,t_4__27_,t_4__26_,t_4__25_,t_4__24_,t_4__23_,t_4__22_,
  t_4__21_,t_4__20_,t_4__19_,t_4__18_,t_4__17_,t_4__16_,t_4__15_,t_4__14_,
  t_4__13_,t_4__12_,t_4__11_,t_4__10_,t_4__9_,t_4__8_,t_4__7_,t_4__6_,t_4__5_,t_4__4_,
  t_4__3_,t_4__2_,t_4__1_,t_4__0_,t_3__55_,t_3__54_,t_3__53_,t_3__52_,t_3__51_,
  t_3__50_,t_3__49_,t_3__48_,t_3__47_,t_3__46_,t_3__45_,t_3__44_,t_3__43_,t_3__42_,
  t_3__41_,t_3__40_,t_3__39_,t_3__38_,t_3__37_,t_3__36_,t_3__35_,t_3__34_,t_3__33_,
  t_3__32_,t_3__31_,t_3__30_,t_3__29_,t_3__28_,t_3__27_,t_3__26_,t_3__25_,t_3__24_,
  t_3__23_,t_3__22_,t_3__21_,t_3__20_,t_3__19_,t_3__18_,t_3__17_,t_3__16_,t_3__15_,
  t_3__14_,t_3__13_,t_3__12_,t_3__11_,t_3__10_,t_3__9_,t_3__8_,t_3__7_,t_3__6_,
  t_3__5_,t_3__4_,t_3__3_,t_3__2_,t_3__1_,t_3__0_,t_2__55_,t_2__54_,t_2__53_,t_2__52_,
  t_2__51_,t_2__50_,t_2__49_,t_2__48_,t_2__47_,t_2__46_,t_2__45_,t_2__44_,t_2__43_,
  t_2__42_,t_2__41_,t_2__40_,t_2__39_,t_2__38_,t_2__37_,t_2__36_,t_2__35_,t_2__34_,
  t_2__33_,t_2__32_,t_2__31_,t_2__30_,t_2__29_,t_2__28_,t_2__27_,t_2__26_,
  t_2__25_,t_2__24_,t_2__23_,t_2__22_,t_2__21_,t_2__20_,t_2__19_,t_2__18_,t_2__17_,
  t_2__16_,t_2__15_,t_2__14_,t_2__13_,t_2__12_,t_2__11_,t_2__10_,t_2__9_,t_2__8_,t_2__7_,
  t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__55_,t_1__54_,
  t_1__53_,t_1__52_,t_1__51_,t_1__50_,t_1__49_,t_1__48_,t_1__47_,t_1__46_,t_1__45_,
  t_1__44_,t_1__43_,t_1__42_,t_1__41_,t_1__40_,t_1__39_,t_1__38_,t_1__37_,t_1__36_,
  t_1__35_,t_1__34_,t_1__33_,t_1__32_,t_1__31_,t_1__30_,t_1__29_,t_1__28_,t_1__27_,
  t_1__26_,t_1__25_,t_1__24_,t_1__23_,t_1__22_,t_1__21_,t_1__20_,t_1__19_,t_1__18_,
  t_1__17_,t_1__16_,t_1__15_,t_1__14_,t_1__13_,t_1__12_,t_1__11_,t_1__10_,t_1__9_,
  t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__55_ = i[0] | 1'b0;
  assign t_1__54_ = i[1] | i[0];
  assign t_1__53_ = i[2] | i[1];
  assign t_1__52_ = i[3] | i[2];
  assign t_1__51_ = i[4] | i[3];
  assign t_1__50_ = i[5] | i[4];
  assign t_1__49_ = i[6] | i[5];
  assign t_1__48_ = i[7] | i[6];
  assign t_1__47_ = i[8] | i[7];
  assign t_1__46_ = i[9] | i[8];
  assign t_1__45_ = i[10] | i[9];
  assign t_1__44_ = i[11] | i[10];
  assign t_1__43_ = i[12] | i[11];
  assign t_1__42_ = i[13] | i[12];
  assign t_1__41_ = i[14] | i[13];
  assign t_1__40_ = i[15] | i[14];
  assign t_1__39_ = i[16] | i[15];
  assign t_1__38_ = i[17] | i[16];
  assign t_1__37_ = i[18] | i[17];
  assign t_1__36_ = i[19] | i[18];
  assign t_1__35_ = i[20] | i[19];
  assign t_1__34_ = i[21] | i[20];
  assign t_1__33_ = i[22] | i[21];
  assign t_1__32_ = i[23] | i[22];
  assign t_1__31_ = i[24] | i[23];
  assign t_1__30_ = i[25] | i[24];
  assign t_1__29_ = i[26] | i[25];
  assign t_1__28_ = i[27] | i[26];
  assign t_1__27_ = i[28] | i[27];
  assign t_1__26_ = i[29] | i[28];
  assign t_1__25_ = i[30] | i[29];
  assign t_1__24_ = i[31] | i[30];
  assign t_1__23_ = i[32] | i[31];
  assign t_1__22_ = i[33] | i[32];
  assign t_1__21_ = i[34] | i[33];
  assign t_1__20_ = i[35] | i[34];
  assign t_1__19_ = i[36] | i[35];
  assign t_1__18_ = i[37] | i[36];
  assign t_1__17_ = i[38] | i[37];
  assign t_1__16_ = i[39] | i[38];
  assign t_1__15_ = i[40] | i[39];
  assign t_1__14_ = i[41] | i[40];
  assign t_1__13_ = i[42] | i[41];
  assign t_1__12_ = i[43] | i[42];
  assign t_1__11_ = i[44] | i[43];
  assign t_1__10_ = i[45] | i[44];
  assign t_1__9_ = i[46] | i[45];
  assign t_1__8_ = i[47] | i[46];
  assign t_1__7_ = i[48] | i[47];
  assign t_1__6_ = i[49] | i[48];
  assign t_1__5_ = i[50] | i[49];
  assign t_1__4_ = i[51] | i[50];
  assign t_1__3_ = i[52] | i[51];
  assign t_1__2_ = i[53] | i[52];
  assign t_1__1_ = i[54] | i[53];
  assign t_1__0_ = i[55] | i[54];
  assign t_2__55_ = t_1__55_ | 1'b0;
  assign t_2__54_ = t_1__54_ | 1'b0;
  assign t_2__53_ = t_1__53_ | t_1__55_;
  assign t_2__52_ = t_1__52_ | t_1__54_;
  assign t_2__51_ = t_1__51_ | t_1__53_;
  assign t_2__50_ = t_1__50_ | t_1__52_;
  assign t_2__49_ = t_1__49_ | t_1__51_;
  assign t_2__48_ = t_1__48_ | t_1__50_;
  assign t_2__47_ = t_1__47_ | t_1__49_;
  assign t_2__46_ = t_1__46_ | t_1__48_;
  assign t_2__45_ = t_1__45_ | t_1__47_;
  assign t_2__44_ = t_1__44_ | t_1__46_;
  assign t_2__43_ = t_1__43_ | t_1__45_;
  assign t_2__42_ = t_1__42_ | t_1__44_;
  assign t_2__41_ = t_1__41_ | t_1__43_;
  assign t_2__40_ = t_1__40_ | t_1__42_;
  assign t_2__39_ = t_1__39_ | t_1__41_;
  assign t_2__38_ = t_1__38_ | t_1__40_;
  assign t_2__37_ = t_1__37_ | t_1__39_;
  assign t_2__36_ = t_1__36_ | t_1__38_;
  assign t_2__35_ = t_1__35_ | t_1__37_;
  assign t_2__34_ = t_1__34_ | t_1__36_;
  assign t_2__33_ = t_1__33_ | t_1__35_;
  assign t_2__32_ = t_1__32_ | t_1__34_;
  assign t_2__31_ = t_1__31_ | t_1__33_;
  assign t_2__30_ = t_1__30_ | t_1__32_;
  assign t_2__29_ = t_1__29_ | t_1__31_;
  assign t_2__28_ = t_1__28_ | t_1__30_;
  assign t_2__27_ = t_1__27_ | t_1__29_;
  assign t_2__26_ = t_1__26_ | t_1__28_;
  assign t_2__25_ = t_1__25_ | t_1__27_;
  assign t_2__24_ = t_1__24_ | t_1__26_;
  assign t_2__23_ = t_1__23_ | t_1__25_;
  assign t_2__22_ = t_1__22_ | t_1__24_;
  assign t_2__21_ = t_1__21_ | t_1__23_;
  assign t_2__20_ = t_1__20_ | t_1__22_;
  assign t_2__19_ = t_1__19_ | t_1__21_;
  assign t_2__18_ = t_1__18_ | t_1__20_;
  assign t_2__17_ = t_1__17_ | t_1__19_;
  assign t_2__16_ = t_1__16_ | t_1__18_;
  assign t_2__15_ = t_1__15_ | t_1__17_;
  assign t_2__14_ = t_1__14_ | t_1__16_;
  assign t_2__13_ = t_1__13_ | t_1__15_;
  assign t_2__12_ = t_1__12_ | t_1__14_;
  assign t_2__11_ = t_1__11_ | t_1__13_;
  assign t_2__10_ = t_1__10_ | t_1__12_;
  assign t_2__9_ = t_1__9_ | t_1__11_;
  assign t_2__8_ = t_1__8_ | t_1__10_;
  assign t_2__7_ = t_1__7_ | t_1__9_;
  assign t_2__6_ = t_1__6_ | t_1__8_;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign t_3__55_ = t_2__55_ | 1'b0;
  assign t_3__54_ = t_2__54_ | 1'b0;
  assign t_3__53_ = t_2__53_ | 1'b0;
  assign t_3__52_ = t_2__52_ | 1'b0;
  assign t_3__51_ = t_2__51_ | t_2__55_;
  assign t_3__50_ = t_2__50_ | t_2__54_;
  assign t_3__49_ = t_2__49_ | t_2__53_;
  assign t_3__48_ = t_2__48_ | t_2__52_;
  assign t_3__47_ = t_2__47_ | t_2__51_;
  assign t_3__46_ = t_2__46_ | t_2__50_;
  assign t_3__45_ = t_2__45_ | t_2__49_;
  assign t_3__44_ = t_2__44_ | t_2__48_;
  assign t_3__43_ = t_2__43_ | t_2__47_;
  assign t_3__42_ = t_2__42_ | t_2__46_;
  assign t_3__41_ = t_2__41_ | t_2__45_;
  assign t_3__40_ = t_2__40_ | t_2__44_;
  assign t_3__39_ = t_2__39_ | t_2__43_;
  assign t_3__38_ = t_2__38_ | t_2__42_;
  assign t_3__37_ = t_2__37_ | t_2__41_;
  assign t_3__36_ = t_2__36_ | t_2__40_;
  assign t_3__35_ = t_2__35_ | t_2__39_;
  assign t_3__34_ = t_2__34_ | t_2__38_;
  assign t_3__33_ = t_2__33_ | t_2__37_;
  assign t_3__32_ = t_2__32_ | t_2__36_;
  assign t_3__31_ = t_2__31_ | t_2__35_;
  assign t_3__30_ = t_2__30_ | t_2__34_;
  assign t_3__29_ = t_2__29_ | t_2__33_;
  assign t_3__28_ = t_2__28_ | t_2__32_;
  assign t_3__27_ = t_2__27_ | t_2__31_;
  assign t_3__26_ = t_2__26_ | t_2__30_;
  assign t_3__25_ = t_2__25_ | t_2__29_;
  assign t_3__24_ = t_2__24_ | t_2__28_;
  assign t_3__23_ = t_2__23_ | t_2__27_;
  assign t_3__22_ = t_2__22_ | t_2__26_;
  assign t_3__21_ = t_2__21_ | t_2__25_;
  assign t_3__20_ = t_2__20_ | t_2__24_;
  assign t_3__19_ = t_2__19_ | t_2__23_;
  assign t_3__18_ = t_2__18_ | t_2__22_;
  assign t_3__17_ = t_2__17_ | t_2__21_;
  assign t_3__16_ = t_2__16_ | t_2__20_;
  assign t_3__15_ = t_2__15_ | t_2__19_;
  assign t_3__14_ = t_2__14_ | t_2__18_;
  assign t_3__13_ = t_2__13_ | t_2__17_;
  assign t_3__12_ = t_2__12_ | t_2__16_;
  assign t_3__11_ = t_2__11_ | t_2__15_;
  assign t_3__10_ = t_2__10_ | t_2__14_;
  assign t_3__9_ = t_2__9_ | t_2__13_;
  assign t_3__8_ = t_2__8_ | t_2__12_;
  assign t_3__7_ = t_2__7_ | t_2__11_;
  assign t_3__6_ = t_2__6_ | t_2__10_;
  assign t_3__5_ = t_2__5_ | t_2__9_;
  assign t_3__4_ = t_2__4_ | t_2__8_;
  assign t_3__3_ = t_2__3_ | t_2__7_;
  assign t_3__2_ = t_2__2_ | t_2__6_;
  assign t_3__1_ = t_2__1_ | t_2__5_;
  assign t_3__0_ = t_2__0_ | t_2__4_;
  assign t_4__55_ = t_3__55_ | 1'b0;
  assign t_4__54_ = t_3__54_ | 1'b0;
  assign t_4__53_ = t_3__53_ | 1'b0;
  assign t_4__52_ = t_3__52_ | 1'b0;
  assign t_4__51_ = t_3__51_ | 1'b0;
  assign t_4__50_ = t_3__50_ | 1'b0;
  assign t_4__49_ = t_3__49_ | 1'b0;
  assign t_4__48_ = t_3__48_ | 1'b0;
  assign t_4__47_ = t_3__47_ | t_3__55_;
  assign t_4__46_ = t_3__46_ | t_3__54_;
  assign t_4__45_ = t_3__45_ | t_3__53_;
  assign t_4__44_ = t_3__44_ | t_3__52_;
  assign t_4__43_ = t_3__43_ | t_3__51_;
  assign t_4__42_ = t_3__42_ | t_3__50_;
  assign t_4__41_ = t_3__41_ | t_3__49_;
  assign t_4__40_ = t_3__40_ | t_3__48_;
  assign t_4__39_ = t_3__39_ | t_3__47_;
  assign t_4__38_ = t_3__38_ | t_3__46_;
  assign t_4__37_ = t_3__37_ | t_3__45_;
  assign t_4__36_ = t_3__36_ | t_3__44_;
  assign t_4__35_ = t_3__35_ | t_3__43_;
  assign t_4__34_ = t_3__34_ | t_3__42_;
  assign t_4__33_ = t_3__33_ | t_3__41_;
  assign t_4__32_ = t_3__32_ | t_3__40_;
  assign t_4__31_ = t_3__31_ | t_3__39_;
  assign t_4__30_ = t_3__30_ | t_3__38_;
  assign t_4__29_ = t_3__29_ | t_3__37_;
  assign t_4__28_ = t_3__28_ | t_3__36_;
  assign t_4__27_ = t_3__27_ | t_3__35_;
  assign t_4__26_ = t_3__26_ | t_3__34_;
  assign t_4__25_ = t_3__25_ | t_3__33_;
  assign t_4__24_ = t_3__24_ | t_3__32_;
  assign t_4__23_ = t_3__23_ | t_3__31_;
  assign t_4__22_ = t_3__22_ | t_3__30_;
  assign t_4__21_ = t_3__21_ | t_3__29_;
  assign t_4__20_ = t_3__20_ | t_3__28_;
  assign t_4__19_ = t_3__19_ | t_3__27_;
  assign t_4__18_ = t_3__18_ | t_3__26_;
  assign t_4__17_ = t_3__17_ | t_3__25_;
  assign t_4__16_ = t_3__16_ | t_3__24_;
  assign t_4__15_ = t_3__15_ | t_3__23_;
  assign t_4__14_ = t_3__14_ | t_3__22_;
  assign t_4__13_ = t_3__13_ | t_3__21_;
  assign t_4__12_ = t_3__12_ | t_3__20_;
  assign t_4__11_ = t_3__11_ | t_3__19_;
  assign t_4__10_ = t_3__10_ | t_3__18_;
  assign t_4__9_ = t_3__9_ | t_3__17_;
  assign t_4__8_ = t_3__8_ | t_3__16_;
  assign t_4__7_ = t_3__7_ | t_3__15_;
  assign t_4__6_ = t_3__6_ | t_3__14_;
  assign t_4__5_ = t_3__5_ | t_3__13_;
  assign t_4__4_ = t_3__4_ | t_3__12_;
  assign t_4__3_ = t_3__3_ | t_3__11_;
  assign t_4__2_ = t_3__2_ | t_3__10_;
  assign t_4__1_ = t_3__1_ | t_3__9_;
  assign t_4__0_ = t_3__0_ | t_3__8_;
  assign t_5__55_ = t_4__55_ | 1'b0;
  assign t_5__54_ = t_4__54_ | 1'b0;
  assign t_5__53_ = t_4__53_ | 1'b0;
  assign t_5__52_ = t_4__52_ | 1'b0;
  assign t_5__51_ = t_4__51_ | 1'b0;
  assign t_5__50_ = t_4__50_ | 1'b0;
  assign t_5__49_ = t_4__49_ | 1'b0;
  assign t_5__48_ = t_4__48_ | 1'b0;
  assign t_5__47_ = t_4__47_ | 1'b0;
  assign t_5__46_ = t_4__46_ | 1'b0;
  assign t_5__45_ = t_4__45_ | 1'b0;
  assign t_5__44_ = t_4__44_ | 1'b0;
  assign t_5__43_ = t_4__43_ | 1'b0;
  assign t_5__42_ = t_4__42_ | 1'b0;
  assign t_5__41_ = t_4__41_ | 1'b0;
  assign t_5__40_ = t_4__40_ | 1'b0;
  assign t_5__39_ = t_4__39_ | t_4__55_;
  assign t_5__38_ = t_4__38_ | t_4__54_;
  assign t_5__37_ = t_4__37_ | t_4__53_;
  assign t_5__36_ = t_4__36_ | t_4__52_;
  assign t_5__35_ = t_4__35_ | t_4__51_;
  assign t_5__34_ = t_4__34_ | t_4__50_;
  assign t_5__33_ = t_4__33_ | t_4__49_;
  assign t_5__32_ = t_4__32_ | t_4__48_;
  assign t_5__31_ = t_4__31_ | t_4__47_;
  assign t_5__30_ = t_4__30_ | t_4__46_;
  assign t_5__29_ = t_4__29_ | t_4__45_;
  assign t_5__28_ = t_4__28_ | t_4__44_;
  assign t_5__27_ = t_4__27_ | t_4__43_;
  assign t_5__26_ = t_4__26_ | t_4__42_;
  assign t_5__25_ = t_4__25_ | t_4__41_;
  assign t_5__24_ = t_4__24_ | t_4__40_;
  assign t_5__23_ = t_4__23_ | t_4__39_;
  assign t_5__22_ = t_4__22_ | t_4__38_;
  assign t_5__21_ = t_4__21_ | t_4__37_;
  assign t_5__20_ = t_4__20_ | t_4__36_;
  assign t_5__19_ = t_4__19_ | t_4__35_;
  assign t_5__18_ = t_4__18_ | t_4__34_;
  assign t_5__17_ = t_4__17_ | t_4__33_;
  assign t_5__16_ = t_4__16_ | t_4__32_;
  assign t_5__15_ = t_4__15_ | t_4__31_;
  assign t_5__14_ = t_4__14_ | t_4__30_;
  assign t_5__13_ = t_4__13_ | t_4__29_;
  assign t_5__12_ = t_4__12_ | t_4__28_;
  assign t_5__11_ = t_4__11_ | t_4__27_;
  assign t_5__10_ = t_4__10_ | t_4__26_;
  assign t_5__9_ = t_4__9_ | t_4__25_;
  assign t_5__8_ = t_4__8_ | t_4__24_;
  assign t_5__7_ = t_4__7_ | t_4__23_;
  assign t_5__6_ = t_4__6_ | t_4__22_;
  assign t_5__5_ = t_4__5_ | t_4__21_;
  assign t_5__4_ = t_4__4_ | t_4__20_;
  assign t_5__3_ = t_4__3_ | t_4__19_;
  assign t_5__2_ = t_4__2_ | t_4__18_;
  assign t_5__1_ = t_4__1_ | t_4__17_;
  assign t_5__0_ = t_4__0_ | t_4__16_;
  assign o[0] = t_5__55_ | 1'b0;
  assign o[1] = t_5__54_ | 1'b0;
  assign o[2] = t_5__53_ | 1'b0;
  assign o[3] = t_5__52_ | 1'b0;
  assign o[4] = t_5__51_ | 1'b0;
  assign o[5] = t_5__50_ | 1'b0;
  assign o[6] = t_5__49_ | 1'b0;
  assign o[7] = t_5__48_ | 1'b0;
  assign o[8] = t_5__47_ | 1'b0;
  assign o[9] = t_5__46_ | 1'b0;
  assign o[10] = t_5__45_ | 1'b0;
  assign o[11] = t_5__44_ | 1'b0;
  assign o[12] = t_5__43_ | 1'b0;
  assign o[13] = t_5__42_ | 1'b0;
  assign o[14] = t_5__41_ | 1'b0;
  assign o[15] = t_5__40_ | 1'b0;
  assign o[16] = t_5__39_ | 1'b0;
  assign o[17] = t_5__38_ | 1'b0;
  assign o[18] = t_5__37_ | 1'b0;
  assign o[19] = t_5__36_ | 1'b0;
  assign o[20] = t_5__35_ | 1'b0;
  assign o[21] = t_5__34_ | 1'b0;
  assign o[22] = t_5__33_ | 1'b0;
  assign o[23] = t_5__32_ | 1'b0;
  assign o[24] = t_5__31_ | 1'b0;
  assign o[25] = t_5__30_ | 1'b0;
  assign o[26] = t_5__29_ | 1'b0;
  assign o[27] = t_5__28_ | 1'b0;
  assign o[28] = t_5__27_ | 1'b0;
  assign o[29] = t_5__26_ | 1'b0;
  assign o[30] = t_5__25_ | 1'b0;
  assign o[31] = t_5__24_ | 1'b0;
  assign o[32] = t_5__23_ | t_5__55_;
  assign o[33] = t_5__22_ | t_5__54_;
  assign o[34] = t_5__21_ | t_5__53_;
  assign o[35] = t_5__20_ | t_5__52_;
  assign o[36] = t_5__19_ | t_5__51_;
  assign o[37] = t_5__18_ | t_5__50_;
  assign o[38] = t_5__17_ | t_5__49_;
  assign o[39] = t_5__16_ | t_5__48_;
  assign o[40] = t_5__15_ | t_5__47_;
  assign o[41] = t_5__14_ | t_5__46_;
  assign o[42] = t_5__13_ | t_5__45_;
  assign o[43] = t_5__12_ | t_5__44_;
  assign o[44] = t_5__11_ | t_5__43_;
  assign o[45] = t_5__10_ | t_5__42_;
  assign o[46] = t_5__9_ | t_5__41_;
  assign o[47] = t_5__8_ | t_5__40_;
  assign o[48] = t_5__7_ | t_5__39_;
  assign o[49] = t_5__6_ | t_5__38_;
  assign o[50] = t_5__5_ | t_5__37_;
  assign o[51] = t_5__4_ | t_5__36_;
  assign o[52] = t_5__3_ | t_5__35_;
  assign o[53] = t_5__2_ | t_5__34_;
  assign o[54] = t_5__1_ | t_5__33_;
  assign o[55] = t_5__0_ | t_5__32_;

endmodule



module bsg_priority_encode_one_hot_out_width_p56_lo_to_hi_p1
(
  i,
  o,
  v_o
);

  input [55:0] i;
  output [55:0] o;
  output v_o;
  wire [55:0] o;
  wire v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54;
  wire [54:1] scan_lo;

  bsg_scan_width_p56_or_p1_lo_to_hi_p1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, scan_lo, o[0:0] })
  );

  assign o[55] = v_o & N0;
  assign N0 = ~scan_lo[54];
  assign o[54] = scan_lo[54] & N1;
  assign N1 = ~scan_lo[53];
  assign o[53] = scan_lo[53] & N2;
  assign N2 = ~scan_lo[52];
  assign o[52] = scan_lo[52] & N3;
  assign N3 = ~scan_lo[51];
  assign o[51] = scan_lo[51] & N4;
  assign N4 = ~scan_lo[50];
  assign o[50] = scan_lo[50] & N5;
  assign N5 = ~scan_lo[49];
  assign o[49] = scan_lo[49] & N6;
  assign N6 = ~scan_lo[48];
  assign o[48] = scan_lo[48] & N7;
  assign N7 = ~scan_lo[47];
  assign o[47] = scan_lo[47] & N8;
  assign N8 = ~scan_lo[46];
  assign o[46] = scan_lo[46] & N9;
  assign N9 = ~scan_lo[45];
  assign o[45] = scan_lo[45] & N10;
  assign N10 = ~scan_lo[44];
  assign o[44] = scan_lo[44] & N11;
  assign N11 = ~scan_lo[43];
  assign o[43] = scan_lo[43] & N12;
  assign N12 = ~scan_lo[42];
  assign o[42] = scan_lo[42] & N13;
  assign N13 = ~scan_lo[41];
  assign o[41] = scan_lo[41] & N14;
  assign N14 = ~scan_lo[40];
  assign o[40] = scan_lo[40] & N15;
  assign N15 = ~scan_lo[39];
  assign o[39] = scan_lo[39] & N16;
  assign N16 = ~scan_lo[38];
  assign o[38] = scan_lo[38] & N17;
  assign N17 = ~scan_lo[37];
  assign o[37] = scan_lo[37] & N18;
  assign N18 = ~scan_lo[36];
  assign o[36] = scan_lo[36] & N19;
  assign N19 = ~scan_lo[35];
  assign o[35] = scan_lo[35] & N20;
  assign N20 = ~scan_lo[34];
  assign o[34] = scan_lo[34] & N21;
  assign N21 = ~scan_lo[33];
  assign o[33] = scan_lo[33] & N22;
  assign N22 = ~scan_lo[32];
  assign o[32] = scan_lo[32] & N23;
  assign N23 = ~scan_lo[31];
  assign o[31] = scan_lo[31] & N24;
  assign N24 = ~scan_lo[30];
  assign o[30] = scan_lo[30] & N25;
  assign N25 = ~scan_lo[29];
  assign o[29] = scan_lo[29] & N26;
  assign N26 = ~scan_lo[28];
  assign o[28] = scan_lo[28] & N27;
  assign N27 = ~scan_lo[27];
  assign o[27] = scan_lo[27] & N28;
  assign N28 = ~scan_lo[26];
  assign o[26] = scan_lo[26] & N29;
  assign N29 = ~scan_lo[25];
  assign o[25] = scan_lo[25] & N30;
  assign N30 = ~scan_lo[24];
  assign o[24] = scan_lo[24] & N31;
  assign N31 = ~scan_lo[23];
  assign o[23] = scan_lo[23] & N32;
  assign N32 = ~scan_lo[22];
  assign o[22] = scan_lo[22] & N33;
  assign N33 = ~scan_lo[21];
  assign o[21] = scan_lo[21] & N34;
  assign N34 = ~scan_lo[20];
  assign o[20] = scan_lo[20] & N35;
  assign N35 = ~scan_lo[19];
  assign o[19] = scan_lo[19] & N36;
  assign N36 = ~scan_lo[18];
  assign o[18] = scan_lo[18] & N37;
  assign N37 = ~scan_lo[17];
  assign o[17] = scan_lo[17] & N38;
  assign N38 = ~scan_lo[16];
  assign o[16] = scan_lo[16] & N39;
  assign N39 = ~scan_lo[15];
  assign o[15] = scan_lo[15] & N40;
  assign N40 = ~scan_lo[14];
  assign o[14] = scan_lo[14] & N41;
  assign N41 = ~scan_lo[13];
  assign o[13] = scan_lo[13] & N42;
  assign N42 = ~scan_lo[12];
  assign o[12] = scan_lo[12] & N43;
  assign N43 = ~scan_lo[11];
  assign o[11] = scan_lo[11] & N44;
  assign N44 = ~scan_lo[10];
  assign o[10] = scan_lo[10] & N45;
  assign N45 = ~scan_lo[9];
  assign o[9] = scan_lo[9] & N46;
  assign N46 = ~scan_lo[8];
  assign o[8] = scan_lo[8] & N47;
  assign N47 = ~scan_lo[7];
  assign o[7] = scan_lo[7] & N48;
  assign N48 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N49;
  assign N49 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N50;
  assign N50 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N51;
  assign N51 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N52;
  assign N52 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N53;
  assign N53 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N54;
  assign N54 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p56_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [55:0] i;
  output [5:0] addr_o;
  output v_o;
  wire [5:0] addr_o;
  wire v_o,v_5__0_,v_4__48_,v_4__32_,v_4__16_,v_4__0_,v_3__56_,v_3__48_,v_3__40_,
  v_3__32_,v_3__24_,v_3__16_,v_3__8_,v_3__0_,v_2__60_,v_2__56_,v_2__52_,v_2__48_,
  v_2__44_,v_2__40_,v_2__36_,v_2__32_,v_2__28_,v_2__24_,v_2__20_,v_2__16_,v_2__12_,
  v_2__8_,v_2__4_,v_2__0_,v_1__62_,v_1__60_,v_1__58_,v_1__56_,v_1__54_,v_1__52_,
  v_1__50_,v_1__48_,v_1__46_,v_1__44_,v_1__42_,v_1__40_,v_1__38_,v_1__36_,v_1__34_,
  v_1__32_,v_1__30_,v_1__28_,v_1__26_,v_1__24_,v_1__22_,v_1__20_,v_1__18_,v_1__16_,
  v_1__14_,v_1__12_,v_1__10_,v_1__8_,v_1__6_,v_1__4_,v_1__2_,v_1__0_,addr_5__35_,
  addr_5__34_,addr_5__33_,addr_5__32_,addr_5__3_,addr_5__2_,addr_5__1_,addr_5__0_,
  addr_4__50_,addr_4__49_,addr_4__48_,addr_4__34_,addr_4__33_,addr_4__32_,addr_4__18_,
  addr_4__17_,addr_4__16_,addr_4__2_,addr_4__1_,addr_4__0_,addr_3__57_,addr_3__56_,
  addr_3__49_,addr_3__48_,addr_3__41_,addr_3__40_,addr_3__33_,addr_3__32_,
  addr_3__25_,addr_3__24_,addr_3__17_,addr_3__16_,addr_3__9_,addr_3__8_,addr_3__1_,
  addr_3__0_,addr_2__60_,addr_2__56_,addr_2__52_,addr_2__48_,addr_2__44_,addr_2__40_,
  addr_2__36_,addr_2__32_,addr_2__28_,addr_2__24_,addr_2__20_,addr_2__16_,addr_2__12_,
  addr_2__8_,addr_2__4_,addr_2__0_;
  assign v_1__0_ = i[1] | i[0];
  assign v_1__2_ = i[3] | i[2];
  assign v_1__4_ = i[5] | i[4];
  assign v_1__6_ = i[7] | i[6];
  assign v_1__8_ = i[9] | i[8];
  assign v_1__10_ = i[11] | i[10];
  assign v_1__12_ = i[13] | i[12];
  assign v_1__14_ = i[15] | i[14];
  assign v_1__16_ = i[17] | i[16];
  assign v_1__18_ = i[19] | i[18];
  assign v_1__20_ = i[21] | i[20];
  assign v_1__22_ = i[23] | i[22];
  assign v_1__24_ = i[25] | i[24];
  assign v_1__26_ = i[27] | i[26];
  assign v_1__28_ = i[29] | i[28];
  assign v_1__30_ = i[31] | i[30];
  assign v_1__32_ = i[33] | i[32];
  assign v_1__34_ = i[35] | i[34];
  assign v_1__36_ = i[37] | i[36];
  assign v_1__38_ = i[39] | i[38];
  assign v_1__40_ = i[41] | i[40];
  assign v_1__42_ = i[43] | i[42];
  assign v_1__44_ = i[45] | i[44];
  assign v_1__46_ = i[47] | i[46];
  assign v_1__48_ = i[49] | i[48];
  assign v_1__50_ = i[51] | i[50];
  assign v_1__52_ = i[53] | i[52];
  assign v_1__54_ = i[55] | i[54];
  assign v_1__56_ = 1'b0 | 1'b0;
  assign v_1__58_ = 1'b0 | 1'b0;
  assign v_1__60_ = 1'b0 | 1'b0;
  assign v_1__62_ = 1'b0 | 1'b0;
  assign v_2__0_ = v_1__2_ | v_1__0_;
  assign addr_2__0_ = i[1] | i[3];
  assign v_2__4_ = v_1__6_ | v_1__4_;
  assign addr_2__4_ = i[5] | i[7];
  assign v_2__8_ = v_1__10_ | v_1__8_;
  assign addr_2__8_ = i[9] | i[11];
  assign v_2__12_ = v_1__14_ | v_1__12_;
  assign addr_2__12_ = i[13] | i[15];
  assign v_2__16_ = v_1__18_ | v_1__16_;
  assign addr_2__16_ = i[17] | i[19];
  assign v_2__20_ = v_1__22_ | v_1__20_;
  assign addr_2__20_ = i[21] | i[23];
  assign v_2__24_ = v_1__26_ | v_1__24_;
  assign addr_2__24_ = i[25] | i[27];
  assign v_2__28_ = v_1__30_ | v_1__28_;
  assign addr_2__28_ = i[29] | i[31];
  assign v_2__32_ = v_1__34_ | v_1__32_;
  assign addr_2__32_ = i[33] | i[35];
  assign v_2__36_ = v_1__38_ | v_1__36_;
  assign addr_2__36_ = i[37] | i[39];
  assign v_2__40_ = v_1__42_ | v_1__40_;
  assign addr_2__40_ = i[41] | i[43];
  assign v_2__44_ = v_1__46_ | v_1__44_;
  assign addr_2__44_ = i[45] | i[47];
  assign v_2__48_ = v_1__50_ | v_1__48_;
  assign addr_2__48_ = i[49] | i[51];
  assign v_2__52_ = v_1__54_ | v_1__52_;
  assign addr_2__52_ = i[53] | i[55];
  assign v_2__56_ = v_1__58_ | v_1__56_;
  assign addr_2__56_ = 1'b0 | 1'b0;
  assign v_2__60_ = v_1__62_ | v_1__60_;
  assign addr_2__60_ = 1'b0 | 1'b0;
  assign v_3__0_ = v_2__4_ | v_2__0_;
  assign addr_3__1_ = v_1__2_ | v_1__6_;
  assign addr_3__0_ = addr_2__0_ | addr_2__4_;
  assign v_3__8_ = v_2__12_ | v_2__8_;
  assign addr_3__9_ = v_1__10_ | v_1__14_;
  assign addr_3__8_ = addr_2__8_ | addr_2__12_;
  assign v_3__16_ = v_2__20_ | v_2__16_;
  assign addr_3__17_ = v_1__18_ | v_1__22_;
  assign addr_3__16_ = addr_2__16_ | addr_2__20_;
  assign v_3__24_ = v_2__28_ | v_2__24_;
  assign addr_3__25_ = v_1__26_ | v_1__30_;
  assign addr_3__24_ = addr_2__24_ | addr_2__28_;
  assign v_3__32_ = v_2__36_ | v_2__32_;
  assign addr_3__33_ = v_1__34_ | v_1__38_;
  assign addr_3__32_ = addr_2__32_ | addr_2__36_;
  assign v_3__40_ = v_2__44_ | v_2__40_;
  assign addr_3__41_ = v_1__42_ | v_1__46_;
  assign addr_3__40_ = addr_2__40_ | addr_2__44_;
  assign v_3__48_ = v_2__52_ | v_2__48_;
  assign addr_3__49_ = v_1__50_ | v_1__54_;
  assign addr_3__48_ = addr_2__48_ | addr_2__52_;
  assign v_3__56_ = v_2__60_ | v_2__56_;
  assign addr_3__57_ = v_1__58_ | v_1__62_;
  assign addr_3__56_ = addr_2__56_ | addr_2__60_;
  assign v_4__0_ = v_3__8_ | v_3__0_;
  assign addr_4__2_ = v_2__4_ | v_2__12_;
  assign addr_4__1_ = addr_3__1_ | addr_3__9_;
  assign addr_4__0_ = addr_3__0_ | addr_3__8_;
  assign v_4__16_ = v_3__24_ | v_3__16_;
  assign addr_4__18_ = v_2__20_ | v_2__28_;
  assign addr_4__17_ = addr_3__17_ | addr_3__25_;
  assign addr_4__16_ = addr_3__16_ | addr_3__24_;
  assign v_4__32_ = v_3__40_ | v_3__32_;
  assign addr_4__34_ = v_2__36_ | v_2__44_;
  assign addr_4__33_ = addr_3__33_ | addr_3__41_;
  assign addr_4__32_ = addr_3__32_ | addr_3__40_;
  assign v_4__48_ = v_3__56_ | v_3__48_;
  assign addr_4__50_ = v_2__52_ | v_2__60_;
  assign addr_4__49_ = addr_3__49_ | addr_3__57_;
  assign addr_4__48_ = addr_3__48_ | addr_3__56_;
  assign v_5__0_ = v_4__16_ | v_4__0_;
  assign addr_5__3_ = v_3__8_ | v_3__24_;
  assign addr_5__2_ = addr_4__2_ | addr_4__18_;
  assign addr_5__1_ = addr_4__1_ | addr_4__17_;
  assign addr_5__0_ = addr_4__0_ | addr_4__16_;
  assign addr_o[5] = v_4__48_ | v_4__32_;
  assign addr_5__35_ = v_3__40_ | v_3__56_;
  assign addr_5__34_ = addr_4__34_ | addr_4__50_;
  assign addr_5__33_ = addr_4__33_ | addr_4__49_;
  assign addr_5__32_ = addr_4__32_ | addr_4__48_;
  assign v_o = addr_o[5] | v_5__0_;
  assign addr_o[4] = v_4__16_ | v_4__48_;
  assign addr_o[3] = addr_5__3_ | addr_5__35_;
  assign addr_o[2] = addr_5__2_ | addr_5__34_;
  assign addr_o[1] = addr_5__1_ | addr_5__33_;
  assign addr_o[0] = addr_5__0_ | addr_5__32_;

endmodule



module bsg_priority_encode_width_p56_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [55:0] i;
  output [5:0] addr_o;
  output v_o;
  wire [5:0] addr_o;
  wire v_o;
  wire [55:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p56_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_width_p56_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o)
  );


endmodule



module bsg_counting_leading_zeros_width_p55
(
  a_i,
  num_zero_o
);

  input [54:0] a_i;
  output [5:0] num_zero_o;
  wire [5:0] num_zero_o;

  bsg_priority_encode_width_p56_lo_to_hi_p1
  pe0
  (
    .i({ 1'b1, a_i[0:0], a_i[1:1], a_i[2:2], a_i[3:3], a_i[4:4], a_i[5:5], a_i[6:6], a_i[7:7], a_i[8:8], a_i[9:9], a_i[10:10], a_i[11:11], a_i[12:12], a_i[13:13], a_i[14:14], a_i[15:15], a_i[16:16], a_i[17:17], a_i[18:18], a_i[19:19], a_i[20:20], a_i[21:21], a_i[22:22], a_i[23:23], a_i[24:24], a_i[25:25], a_i[26:26], a_i[27:27], a_i[28:28], a_i[29:29], a_i[30:30], a_i[31:31], a_i[32:32], a_i[33:33], a_i[34:34], a_i[35:35], a_i[36:36], a_i[37:37], a_i[38:38], a_i[39:39], a_i[40:40], a_i[41:41], a_i[42:42], a_i[43:43], a_i[44:44], a_i[45:45], a_i[46:46], a_i[47:47], a_i[48:48], a_i[49:49], a_i[50:50], a_i[51:51], a_i[52:52], a_i[53:53], a_i[54:54] }),
    .addr_o(num_zero_o)
  );


endmodule



module compressBy2_inWidth27
(
  in,
  out
);

  input [26:0] in;
  output [13:0] out;
  wire [13:0] out;
  wire out_13_;
  assign out_13_ = in[26];
  assign out[13] = out_13_;
  assign out[0] = in[1] | in[0];
  assign out[1] = in[3] | in[2];
  assign out[2] = in[5] | in[4];
  assign out[3] = in[7] | in[6];
  assign out[4] = in[9] | in[8];
  assign out[5] = in[11] | in[10];
  assign out[6] = in[13] | in[12];
  assign out[7] = in[15] | in[14];
  assign out[8] = in[17] | in[16];
  assign out[9] = in[19] | in[18];
  assign out[10] = in[21] | in[20];
  assign out[11] = in[23] | in[22];
  assign out[12] = in[25] | in[24];

endmodule



module lowMaskLoHi_inWidth5_topBound0_bottomBound13
(
  in,
  out
);

  input [4:0] in;
  output [12:0] out;
  wire [12:0] out,reverseOut;
  wire N0,N1,N2,N3,N4,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,
  sv2v_dc_7,sv2v_dc_8,sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,
  sv2v_dc_15,sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19;

  reverse_width13
  reverse
  (
    .in(reverseOut),
    .out(out)
  );

  assign { sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, reverseOut } = $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) >>> { N0, N1, N2, N3, N4 };
  assign N0 = ~in[4];
  assign N1 = ~in[3];
  assign N2 = ~in[2];
  assign N3 = ~in[1];
  assign N4 = ~in[0];

endmodule



module mulAddRecFNToRaw_postMul_expWidth11_sigWidth53
(
  intermed_compactState,
  intermed_sExp,
  intermed_CDom_CAlignDist,
  intermed_highAlignedSigC,
  mulAddResult,
  roundingMode,
  invalidExc,
  out_isNaN,
  out_isInf,
  out_isZero,
  out_sign,
  out_sExp,
  out_sig
);

  input [5:0] intermed_compactState;
  input [12:0] intermed_sExp;
  input [5:0] intermed_CDom_CAlignDist;
  input [54:0] intermed_highAlignedSigC;
  input [106:0] mulAddResult;
  input [2:0] roundingMode;
  output [12:0] out_sExp;
  output [55:0] out_sig;
  output invalidExc;
  output out_isNaN;
  output out_isInf;
  output out_isZero;
  output out_sign;
  wire [12:0] out_sExp,CDom_sExp,CDom_sigExtraMask,notCDom_sExp,notCDom_sigExtraMask;
  wire [55:0] out_sig;
  wire invalidExc,out_isNaN,out_isInf,out_isZero,out_sign,N0,N1,N2,N3,N4,N5,N6,N7,N8,
  notNaN_addZeros,opSignC,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,
  N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,
  N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,
  N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,
  N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,
  N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,
  N119,CDom_absSigSumExtra,N120,CDom_reduced4SigExtra,N121,N122,N123,N124,N125,
  N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,
  N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,
  N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,
  N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,
  N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,
  N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,
  N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,
  N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,
  N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
  N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,
  notCDom_reduced4SigExtra,notCDom_completeCancellation,N284,notCDom_sign,N285,N286,N287,N288,
  N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,
  N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,
  N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
  N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,
  N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
  N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,
  N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,
  N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,
  N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,
  N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,
  N449,N450,N451,N452,N453,N454,N455,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,
  sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,
  sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,
  sv2v_dc_20,sv2v_dc_21,sv2v_dc_22,sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,
  sv2v_dc_27,sv2v_dc_28,sv2v_dc_29,sv2v_dc_30,sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,sv2v_dc_34,
  sv2v_dc_35,sv2v_dc_36,sv2v_dc_37,sv2v_dc_38,sv2v_dc_39,sv2v_dc_40,sv2v_dc_41,
  sv2v_dc_42,sv2v_dc_43,sv2v_dc_44,sv2v_dc_45,sv2v_dc_46,sv2v_dc_47,sv2v_dc_48,
  sv2v_dc_49,sv2v_dc_50,sv2v_dc_51,sv2v_dc_52,sv2v_dc_53,sv2v_dc_54,sv2v_dc_55,
  sv2v_dc_56,sv2v_dc_57,sv2v_dc_58,sv2v_dc_59,sv2v_dc_60,sv2v_dc_61,sv2v_dc_62,sv2v_dc_63,
  sv2v_dc_64,sv2v_dc_65,sv2v_dc_66,sv2v_dc_67,sv2v_dc_68,sv2v_dc_69,sv2v_dc_70,
  sv2v_dc_71,sv2v_dc_72,sv2v_dc_73,sv2v_dc_74,sv2v_dc_75,sv2v_dc_76,sv2v_dc_77,
  sv2v_dc_78,sv2v_dc_79,sv2v_dc_80,sv2v_dc_81,sv2v_dc_82,sv2v_dc_83,sv2v_dc_84,sv2v_dc_85,
  sv2v_dc_86,sv2v_dc_87,sv2v_dc_88,sv2v_dc_89,sv2v_dc_90,sv2v_dc_91,sv2v_dc_92,
  sv2v_dc_93,sv2v_dc_94,sv2v_dc_95,sv2v_dc_96,sv2v_dc_97,sv2v_dc_98,sv2v_dc_99,
  sv2v_dc_100,sv2v_dc_101,sv2v_dc_102;
  wire [54:0] incHighAlignedSigC,notCDom_reduced2AbsSigSum;
  wire [161:107] sigSum;
  wire [107:0] CDom_absSigSum;
  wire [57:0] CDom_mainSig,notCDom_mainSig;
  wire [13:0] CDom_reduced4LowSig,notCDom_reduced4AbsSigSum;
  wire [0:0] CDom_sig,notCDom_sig;
  wire [108:0] notCDom_absSigSum;
  wire [5:0] notCDom_normDistReduced2;
  assign { CDom_mainSig, sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36, sv2v_dc_37, sv2v_dc_38, sv2v_dc_39, sv2v_dc_40, sv2v_dc_41, sv2v_dc_42, sv2v_dc_43, sv2v_dc_44, sv2v_dc_45, sv2v_dc_46, sv2v_dc_47, sv2v_dc_48, sv2v_dc_49, sv2v_dc_50 } = CDom_absSigSum << intermed_CDom_CAlignDist;

  compressBy4_inWidth55
  compressBy4_CDom_absSigSum
  (
    .in({ CDom_absSigSum[52:0], 1'b0, 1'b0 }),
    .out(CDom_reduced4LowSig)
  );


  lowMaskLoHi_inWidth4_topBound0_bottomBound13
  lowMask_CDom_sigExtraMask
  (
    .in(intermed_CDom_CAlignDist[5:2]),
    .out(CDom_sigExtraMask)
  );


  compressBy2_inWidth109
  compressBy2_notCDom_absSigSum
  (
    .in(notCDom_absSigSum),
    .out(notCDom_reduced2AbsSigSum)
  );


  bsg_counting_leading_zeros_width_p55
  clz
  (
    .a_i(notCDom_reduced2AbsSigSum),
    .num_zero_o(notCDom_normDistReduced2)
  );

  assign { notCDom_mainSig, sv2v_dc_51, sv2v_dc_52, sv2v_dc_53, sv2v_dc_54, sv2v_dc_55, sv2v_dc_56, sv2v_dc_57, sv2v_dc_58, sv2v_dc_59, sv2v_dc_60, sv2v_dc_61, sv2v_dc_62, sv2v_dc_63, sv2v_dc_64, sv2v_dc_65, sv2v_dc_66, sv2v_dc_67, sv2v_dc_68, sv2v_dc_69, sv2v_dc_70, sv2v_dc_71, sv2v_dc_72, sv2v_dc_73, sv2v_dc_74, sv2v_dc_75, sv2v_dc_76, sv2v_dc_77, sv2v_dc_78, sv2v_dc_79, sv2v_dc_80, sv2v_dc_81, sv2v_dc_82, sv2v_dc_83, sv2v_dc_84, sv2v_dc_85, sv2v_dc_86, sv2v_dc_87, sv2v_dc_88, sv2v_dc_89, sv2v_dc_90, sv2v_dc_91, sv2v_dc_92, sv2v_dc_93, sv2v_dc_94, sv2v_dc_95, sv2v_dc_96, sv2v_dc_97, sv2v_dc_98, sv2v_dc_99, sv2v_dc_100, sv2v_dc_101, sv2v_dc_102 } = { 1'b0, notCDom_absSigSum } << { notCDom_normDistReduced2, 1'b0 };

  compressBy2_inWidth27
  compressBy2_notCDom_reduced2AbsSigSum
  (
    .in(notCDom_reduced2AbsSigSum[26:0]),
    .out(notCDom_reduced4AbsSigSum)
  );


  lowMaskLoHi_inWidth5_topBound0_bottomBound13
  lowMask_notCDom_sigExtraMask
  (
    .in(notCDom_normDistReduced2[5:1]),
    .out(notCDom_sigExtraMask)
  );

  assign notCDom_completeCancellation = notCDom_mainSig[57:56] == 1'b0;
  assign N286 = ~roundingMode[1];
  assign N287 = N286 | roundingMode[2];
  assign N288 = roundingMode[0] | N287;
  assign N289 = ~N288;
  assign CDom_sExp = intermed_sExp - intermed_compactState[3];
  assign notCDom_sExp = intermed_sExp - { notCDom_normDistReduced2, 1'b0 };
  assign incHighAlignedSigC = intermed_highAlignedSigC + 1'b1;
  assign { N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175 } = { sigSum[108:107], mulAddResult[105:0], intermed_compactState[1:1] } + intermed_compactState[3];
  assign sigSum = (N0)? incHighAlignedSigC : 
                  (N9)? intermed_highAlignedSigC : 1'b0;
  assign N0 = mulAddResult[106];
  assign CDom_absSigSum = (N1)? { N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117 } : 
                          (N2)? { 1'b0, intermed_highAlignedSigC[54:53], sigSum[159:107], mulAddResult[105:54] } : 1'b0;
  assign N1 = intermed_compactState[3];
  assign N2 = N118;
  assign CDom_absSigSumExtra = (N1)? N119 : 
                               (N2)? N120 : 1'b0;
  assign notCDom_absSigSum = (N3)? { N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174 } : 
                             (N4)? { N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175 } : 1'b0;
  assign N3 = sigSum[109];
  assign N4 = N62;
  assign notCDom_sign = (N5)? N289 : 
                        (N6)? N285 : 1'b0;
  assign N5 = notCDom_completeCancellation;
  assign N6 = N284;
  assign out_sExp = (N7)? CDom_sExp : 
                    (N8)? notCDom_sExp : 1'b0;
  assign N7 = intermed_compactState[2];
  assign N8 = N447;
  assign out_sig = (N7)? { CDom_mainSig[57:3], CDom_sig[0:0] } : 
                   (N8)? { notCDom_mainSig[57:3], notCDom_sig[0:0] } : 1'b0;
  assign invalidExc = intermed_compactState[5] & intermed_compactState[4];
  assign out_isNaN = intermed_compactState[5] & intermed_compactState[3];
  assign out_isInf = intermed_compactState[5] & intermed_compactState[2];
  assign notNaN_addZeros = intermed_compactState[5] & intermed_compactState[1];
  assign opSignC = intermed_compactState[4] ^ intermed_compactState[3];
  assign N9 = ~mulAddResult[106];
  assign N10 = ~sigSum[161];
  assign N11 = ~sigSum[160];
  assign N12 = ~sigSum[159];
  assign N13 = ~sigSum[158];
  assign N14 = ~sigSum[157];
  assign N15 = ~sigSum[156];
  assign N16 = ~sigSum[155];
  assign N17 = ~sigSum[154];
  assign N18 = ~sigSum[153];
  assign N19 = ~sigSum[152];
  assign N20 = ~sigSum[151];
  assign N21 = ~sigSum[150];
  assign N22 = ~sigSum[149];
  assign N23 = ~sigSum[148];
  assign N24 = ~sigSum[147];
  assign N25 = ~sigSum[146];
  assign N26 = ~sigSum[145];
  assign N27 = ~sigSum[144];
  assign N28 = ~sigSum[143];
  assign N29 = ~sigSum[142];
  assign N30 = ~sigSum[141];
  assign N31 = ~sigSum[140];
  assign N32 = ~sigSum[139];
  assign N33 = ~sigSum[138];
  assign N34 = ~sigSum[137];
  assign N35 = ~sigSum[136];
  assign N36 = ~sigSum[135];
  assign N37 = ~sigSum[134];
  assign N38 = ~sigSum[133];
  assign N39 = ~sigSum[132];
  assign N40 = ~sigSum[131];
  assign N41 = ~sigSum[130];
  assign N42 = ~sigSum[129];
  assign N43 = ~sigSum[128];
  assign N44 = ~sigSum[127];
  assign N45 = ~sigSum[126];
  assign N46 = ~sigSum[125];
  assign N47 = ~sigSum[124];
  assign N48 = ~sigSum[123];
  assign N49 = ~sigSum[122];
  assign N50 = ~sigSum[121];
  assign N51 = ~sigSum[120];
  assign N52 = ~sigSum[119];
  assign N53 = ~sigSum[118];
  assign N54 = ~sigSum[117];
  assign N55 = ~sigSum[116];
  assign N56 = ~sigSum[115];
  assign N57 = ~sigSum[114];
  assign N58 = ~sigSum[113];
  assign N59 = ~sigSum[112];
  assign N60 = ~sigSum[111];
  assign N61 = ~sigSum[110];
  assign N62 = ~sigSum[109];
  assign N63 = ~sigSum[108];
  assign N64 = ~sigSum[107];
  assign N65 = ~mulAddResult[105];
  assign N66 = ~mulAddResult[104];
  assign N67 = ~mulAddResult[103];
  assign N68 = ~mulAddResult[102];
  assign N69 = ~mulAddResult[101];
  assign N70 = ~mulAddResult[100];
  assign N71 = ~mulAddResult[99];
  assign N72 = ~mulAddResult[98];
  assign N73 = ~mulAddResult[97];
  assign N74 = ~mulAddResult[96];
  assign N75 = ~mulAddResult[95];
  assign N76 = ~mulAddResult[94];
  assign N77 = ~mulAddResult[93];
  assign N78 = ~mulAddResult[92];
  assign N79 = ~mulAddResult[91];
  assign N80 = ~mulAddResult[90];
  assign N81 = ~mulAddResult[89];
  assign N82 = ~mulAddResult[88];
  assign N83 = ~mulAddResult[87];
  assign N84 = ~mulAddResult[86];
  assign N85 = ~mulAddResult[85];
  assign N86 = ~mulAddResult[84];
  assign N87 = ~mulAddResult[83];
  assign N88 = ~mulAddResult[82];
  assign N89 = ~mulAddResult[81];
  assign N90 = ~mulAddResult[80];
  assign N91 = ~mulAddResult[79];
  assign N92 = ~mulAddResult[78];
  assign N93 = ~mulAddResult[77];
  assign N94 = ~mulAddResult[76];
  assign N95 = ~mulAddResult[75];
  assign N96 = ~mulAddResult[74];
  assign N97 = ~mulAddResult[73];
  assign N98 = ~mulAddResult[72];
  assign N99 = ~mulAddResult[71];
  assign N100 = ~mulAddResult[70];
  assign N101 = ~mulAddResult[69];
  assign N102 = ~mulAddResult[68];
  assign N103 = ~mulAddResult[67];
  assign N104 = ~mulAddResult[66];
  assign N105 = ~mulAddResult[65];
  assign N106 = ~mulAddResult[64];
  assign N107 = ~mulAddResult[63];
  assign N108 = ~mulAddResult[62];
  assign N109 = ~mulAddResult[61];
  assign N110 = ~mulAddResult[60];
  assign N111 = ~mulAddResult[59];
  assign N112 = ~mulAddResult[58];
  assign N113 = ~mulAddResult[57];
  assign N114 = ~mulAddResult[56];
  assign N115 = ~mulAddResult[55];
  assign N116 = ~mulAddResult[54];
  assign N117 = ~mulAddResult[53];
  assign N118 = ~intermed_compactState[3];
  assign N119 = ~N341;
  assign N341 = N340 & mulAddResult[0];
  assign N340 = N339 & mulAddResult[1];
  assign N339 = N338 & mulAddResult[2];
  assign N338 = N337 & mulAddResult[3];
  assign N337 = N336 & mulAddResult[4];
  assign N336 = N335 & mulAddResult[5];
  assign N335 = N334 & mulAddResult[6];
  assign N334 = N333 & mulAddResult[7];
  assign N333 = N332 & mulAddResult[8];
  assign N332 = N331 & mulAddResult[9];
  assign N331 = N330 & mulAddResult[10];
  assign N330 = N329 & mulAddResult[11];
  assign N329 = N328 & mulAddResult[12];
  assign N328 = N327 & mulAddResult[13];
  assign N327 = N326 & mulAddResult[14];
  assign N326 = N325 & mulAddResult[15];
  assign N325 = N324 & mulAddResult[16];
  assign N324 = N323 & mulAddResult[17];
  assign N323 = N322 & mulAddResult[18];
  assign N322 = N321 & mulAddResult[19];
  assign N321 = N320 & mulAddResult[20];
  assign N320 = N319 & mulAddResult[21];
  assign N319 = N318 & mulAddResult[22];
  assign N318 = N317 & mulAddResult[23];
  assign N317 = N316 & mulAddResult[24];
  assign N316 = N315 & mulAddResult[25];
  assign N315 = N314 & mulAddResult[26];
  assign N314 = N313 & mulAddResult[27];
  assign N313 = N312 & mulAddResult[28];
  assign N312 = N311 & mulAddResult[29];
  assign N311 = N310 & mulAddResult[30];
  assign N310 = N309 & mulAddResult[31];
  assign N309 = N308 & mulAddResult[32];
  assign N308 = N307 & mulAddResult[33];
  assign N307 = N306 & mulAddResult[34];
  assign N306 = N305 & mulAddResult[35];
  assign N305 = N304 & mulAddResult[36];
  assign N304 = N303 & mulAddResult[37];
  assign N303 = N302 & mulAddResult[38];
  assign N302 = N301 & mulAddResult[39];
  assign N301 = N300 & mulAddResult[40];
  assign N300 = N299 & mulAddResult[41];
  assign N299 = N298 & mulAddResult[42];
  assign N298 = N297 & mulAddResult[43];
  assign N297 = N296 & mulAddResult[44];
  assign N296 = N295 & mulAddResult[45];
  assign N295 = N294 & mulAddResult[46];
  assign N294 = N293 & mulAddResult[47];
  assign N293 = N292 & mulAddResult[48];
  assign N292 = N291 & mulAddResult[49];
  assign N291 = N290 & mulAddResult[50];
  assign N290 = mulAddResult[52] & mulAddResult[51];
  assign N120 = N393 | mulAddResult[0];
  assign N393 = N392 | mulAddResult[1];
  assign N392 = N391 | mulAddResult[2];
  assign N391 = N390 | mulAddResult[3];
  assign N390 = N389 | mulAddResult[4];
  assign N389 = N388 | mulAddResult[5];
  assign N388 = N387 | mulAddResult[6];
  assign N387 = N386 | mulAddResult[7];
  assign N386 = N385 | mulAddResult[8];
  assign N385 = N384 | mulAddResult[9];
  assign N384 = N383 | mulAddResult[10];
  assign N383 = N382 | mulAddResult[11];
  assign N382 = N381 | mulAddResult[12];
  assign N381 = N380 | mulAddResult[13];
  assign N380 = N379 | mulAddResult[14];
  assign N379 = N378 | mulAddResult[15];
  assign N378 = N377 | mulAddResult[16];
  assign N377 = N376 | mulAddResult[17];
  assign N376 = N375 | mulAddResult[18];
  assign N375 = N374 | mulAddResult[19];
  assign N374 = N373 | mulAddResult[20];
  assign N373 = N372 | mulAddResult[21];
  assign N372 = N371 | mulAddResult[22];
  assign N371 = N370 | mulAddResult[23];
  assign N370 = N369 | mulAddResult[24];
  assign N369 = N368 | mulAddResult[25];
  assign N368 = N367 | mulAddResult[26];
  assign N367 = N366 | mulAddResult[27];
  assign N366 = N365 | mulAddResult[28];
  assign N365 = N364 | mulAddResult[29];
  assign N364 = N363 | mulAddResult[30];
  assign N363 = N362 | mulAddResult[31];
  assign N362 = N361 | mulAddResult[32];
  assign N361 = N360 | mulAddResult[33];
  assign N360 = N359 | mulAddResult[34];
  assign N359 = N358 | mulAddResult[35];
  assign N358 = N357 | mulAddResult[36];
  assign N357 = N356 | mulAddResult[37];
  assign N356 = N355 | mulAddResult[38];
  assign N355 = N354 | mulAddResult[39];
  assign N354 = N353 | mulAddResult[40];
  assign N353 = N352 | mulAddResult[41];
  assign N352 = N351 | mulAddResult[42];
  assign N351 = N350 | mulAddResult[43];
  assign N350 = N349 | mulAddResult[44];
  assign N349 = N348 | mulAddResult[45];
  assign N348 = N347 | mulAddResult[46];
  assign N347 = N346 | mulAddResult[47];
  assign N346 = N345 | mulAddResult[48];
  assign N345 = N344 | mulAddResult[49];
  assign N344 = N343 | mulAddResult[50];
  assign N343 = N342 | mulAddResult[51];
  assign N342 = mulAddResult[53] | mulAddResult[52];
  assign CDom_reduced4SigExtra = N416 | N417;
  assign N416 = N414 | N415;
  assign N414 = N412 | N413;
  assign N412 = N410 | N411;
  assign N410 = N408 | N409;
  assign N408 = N406 | N407;
  assign N406 = N404 | N405;
  assign N404 = N402 | N403;
  assign N402 = N400 | N401;
  assign N400 = N398 | N399;
  assign N398 = N396 | N397;
  assign N396 = N394 | N395;
  assign N394 = CDom_reduced4LowSig[12] & CDom_sigExtraMask[12];
  assign N395 = CDom_reduced4LowSig[11] & CDom_sigExtraMask[11];
  assign N397 = CDom_reduced4LowSig[10] & CDom_sigExtraMask[10];
  assign N399 = CDom_reduced4LowSig[9] & CDom_sigExtraMask[9];
  assign N401 = CDom_reduced4LowSig[8] & CDom_sigExtraMask[8];
  assign N403 = CDom_reduced4LowSig[7] & CDom_sigExtraMask[7];
  assign N405 = CDom_reduced4LowSig[6] & CDom_sigExtraMask[6];
  assign N407 = CDom_reduced4LowSig[5] & CDom_sigExtraMask[5];
  assign N409 = CDom_reduced4LowSig[4] & CDom_sigExtraMask[4];
  assign N411 = CDom_reduced4LowSig[3] & CDom_sigExtraMask[3];
  assign N413 = CDom_reduced4LowSig[2] & CDom_sigExtraMask[2];
  assign N415 = CDom_reduced4LowSig[1] & CDom_sigExtraMask[1];
  assign N417 = CDom_reduced4LowSig[0] & CDom_sigExtraMask[0];
  assign CDom_sig[0] = N420 | CDom_absSigSumExtra;
  assign N420 = N419 | CDom_reduced4SigExtra;
  assign N419 = N418 | CDom_mainSig[0];
  assign N418 = CDom_mainSig[2] | CDom_mainSig[1];
  assign N121 = ~mulAddResult[52];
  assign N122 = ~mulAddResult[51];
  assign N123 = ~mulAddResult[50];
  assign N124 = ~mulAddResult[49];
  assign N125 = ~mulAddResult[48];
  assign N126 = ~mulAddResult[47];
  assign N127 = ~mulAddResult[46];
  assign N128 = ~mulAddResult[45];
  assign N129 = ~mulAddResult[44];
  assign N130 = ~mulAddResult[43];
  assign N131 = ~mulAddResult[42];
  assign N132 = ~mulAddResult[41];
  assign N133 = ~mulAddResult[40];
  assign N134 = ~mulAddResult[39];
  assign N135 = ~mulAddResult[38];
  assign N136 = ~mulAddResult[37];
  assign N137 = ~mulAddResult[36];
  assign N138 = ~mulAddResult[35];
  assign N139 = ~mulAddResult[34];
  assign N140 = ~mulAddResult[33];
  assign N141 = ~mulAddResult[32];
  assign N142 = ~mulAddResult[31];
  assign N143 = ~mulAddResult[30];
  assign N144 = ~mulAddResult[29];
  assign N145 = ~mulAddResult[28];
  assign N146 = ~mulAddResult[27];
  assign N147 = ~mulAddResult[26];
  assign N148 = ~mulAddResult[25];
  assign N149 = ~mulAddResult[24];
  assign N150 = ~mulAddResult[23];
  assign N151 = ~mulAddResult[22];
  assign N152 = ~mulAddResult[21];
  assign N153 = ~mulAddResult[20];
  assign N154 = ~mulAddResult[19];
  assign N155 = ~mulAddResult[18];
  assign N156 = ~mulAddResult[17];
  assign N157 = ~mulAddResult[16];
  assign N158 = ~mulAddResult[15];
  assign N159 = ~mulAddResult[14];
  assign N160 = ~mulAddResult[13];
  assign N161 = ~mulAddResult[12];
  assign N162 = ~mulAddResult[11];
  assign N163 = ~mulAddResult[10];
  assign N164 = ~mulAddResult[9];
  assign N165 = ~mulAddResult[8];
  assign N166 = ~mulAddResult[7];
  assign N167 = ~mulAddResult[6];
  assign N168 = ~mulAddResult[5];
  assign N169 = ~mulAddResult[4];
  assign N170 = ~mulAddResult[3];
  assign N171 = ~mulAddResult[2];
  assign N172 = ~mulAddResult[1];
  assign N173 = ~mulAddResult[0];
  assign N174 = ~intermed_compactState[1];
  assign notCDom_reduced4SigExtra = N443 | N444;
  assign N443 = N441 | N442;
  assign N441 = N439 | N440;
  assign N439 = N437 | N438;
  assign N437 = N435 | N436;
  assign N435 = N433 | N434;
  assign N433 = N431 | N432;
  assign N431 = N429 | N430;
  assign N429 = N427 | N428;
  assign N427 = N425 | N426;
  assign N425 = N423 | N424;
  assign N423 = N421 | N422;
  assign N421 = notCDom_reduced4AbsSigSum[12] & notCDom_sigExtraMask[12];
  assign N422 = notCDom_reduced4AbsSigSum[11] & notCDom_sigExtraMask[11];
  assign N424 = notCDom_reduced4AbsSigSum[10] & notCDom_sigExtraMask[10];
  assign N426 = notCDom_reduced4AbsSigSum[9] & notCDom_sigExtraMask[9];
  assign N428 = notCDom_reduced4AbsSigSum[8] & notCDom_sigExtraMask[8];
  assign N430 = notCDom_reduced4AbsSigSum[7] & notCDom_sigExtraMask[7];
  assign N432 = notCDom_reduced4AbsSigSum[6] & notCDom_sigExtraMask[6];
  assign N434 = notCDom_reduced4AbsSigSum[5] & notCDom_sigExtraMask[5];
  assign N436 = notCDom_reduced4AbsSigSum[4] & notCDom_sigExtraMask[4];
  assign N438 = notCDom_reduced4AbsSigSum[3] & notCDom_sigExtraMask[3];
  assign N440 = notCDom_reduced4AbsSigSum[2] & notCDom_sigExtraMask[2];
  assign N442 = notCDom_reduced4AbsSigSum[1] & notCDom_sigExtraMask[1];
  assign N444 = notCDom_reduced4AbsSigSum[0] & notCDom_sigExtraMask[0];
  assign notCDom_sig[0] = N446 | notCDom_reduced4SigExtra;
  assign N446 = N445 | notCDom_mainSig[0];
  assign N445 = notCDom_mainSig[2] | notCDom_mainSig[1];
  assign N284 = ~notCDom_completeCancellation;
  assign N285 = intermed_compactState[4] ^ sigSum[109];
  assign out_isZero = notNaN_addZeros | N448;
  assign N448 = N447 & notCDom_completeCancellation;
  assign N447 = ~intermed_compactState[2];
  assign out_sign = N453 | N455;
  assign N453 = N449 | N452;
  assign N449 = intermed_compactState[5] & intermed_compactState[0];
  assign N452 = N451 & opSignC;
  assign N451 = N450 & intermed_compactState[2];
  assign N450 = ~intermed_compactState[5];
  assign N455 = N454 & notCDom_sign;
  assign N454 = N450 & N447;

endmodule



module mulAddRecFNToRaw_expWidth11_sigWidth53_pipelineStages0_imulEn1
(
  clock,
  control,
  op,
  a,
  b,
  c,
  roundingMode,
  invalidExc,
  out_isNaN,
  out_isInf,
  out_isZero,
  out_sign,
  out_sExp,
  out_sig,
  out_imul
);

  input [0:0] control;
  input [2:0] op;
  input [64:0] a;
  input [64:0] b;
  input [64:0] c;
  input [2:0] roundingMode;
  output [12:0] out_sExp;
  output [55:0] out_sig;
  output [63:0] out_imul;
  input clock;
  output invalidExc;
  output out_isNaN;
  output out_isInf;
  output out_isZero;
  output out_sign;
  wire [12:0] out_sExp,intermed_sExp,intermed_sExp_Z;
  wire [55:0] out_sig;
  wire [63:0] out_imul;
  wire invalidExc,out_isNaN,out_isInf,out_isZero,out_sign;
  wire [52:0] mulAddA,mulAddB;
  wire [105:0] mulAddC;
  wire [5:0] intermed_compactState,intermed_CDom_CAlignDist,intermed_compactState_Z,
  intermed_CDom_CAlignDist_Z;
  wire [54:0] intermed_highAlignedSigC,intermed_highAlignedSigC_Z;
  wire [106:64] mulAddResult;
  wire [2:0] roundingMode_Z;

  mulAddRecFNToRaw_preMul_expWidth11_sigWidth53_imulEn1
  mulAddToRaw_preMul
  (
    .control(control[0]),
    .op(op),
    .a(a),
    .b(b),
    .c(c),
    .roundingMode(roundingMode),
    .mulAddA(mulAddA),
    .mulAddB(mulAddB),
    .mulAddC(mulAddC),
    .intermed_compactState(intermed_compactState),
    .intermed_sExp(intermed_sExp),
    .intermed_CDom_CAlignDist(intermed_CDom_CAlignDist),
    .intermed_highAlignedSigC(intermed_highAlignedSigC)
  );


  bsg_mul_add_unsigned_width_a_p53_width_b_p53_width_c_p106_width_o_p107_pipeline_p0
  mulAdd
  (
    .clk_i(clock),
    .a_i(mulAddA),
    .b_i(mulAddB),
    .c_i(mulAddC),
    .o({ mulAddResult, out_imul })
  );


  bsg_dff_chain_width_p83_num_stages_p0
  shuntMulAdd
  (
    .clk_i(clock),
    .data_i({ intermed_compactState, intermed_sExp, intermed_CDom_CAlignDist, intermed_highAlignedSigC, roundingMode }),
    .data_o({ intermed_compactState_Z, intermed_sExp_Z, intermed_CDom_CAlignDist_Z, intermed_highAlignedSigC_Z, roundingMode_Z })
  );


  mulAddRecFNToRaw_postMul_expWidth11_sigWidth53
  mulAddToRaw_postMul
  (
    .intermed_compactState(intermed_compactState_Z),
    .intermed_sExp(intermed_sExp_Z),
    .intermed_CDom_CAlignDist(intermed_CDom_CAlignDist_Z),
    .intermed_highAlignedSigC(intermed_highAlignedSigC_Z),
    .mulAddResult({ mulAddResult, out_imul }),
    .roundingMode(roundingMode_Z),
    .invalidExc(invalidExc),
    .out_isNaN(out_isNaN),
    .out_isInf(out_isInf),
    .out_isZero(out_isZero),
    .out_sign(out_sign),
    .out_sExp(out_sExp),
    .out_sig(out_sig)
  );


endmodule



module bsg_dff_chain_width_p76_num_stages_p0
(
  clk_i,
  data_i,
  data_o
);

  input [75:0] data_i;
  output [75:0] data_o;
  input clk_i;
  wire [75:0] data_o;
  assign data_o[75] = data_i[75];
  assign data_o[74] = data_i[74];
  assign data_o[73] = data_i[73];
  assign data_o[72] = data_i[72];
  assign data_o[71] = data_i[71];
  assign data_o[70] = data_i[70];
  assign data_o[69] = data_i[69];
  assign data_o[68] = data_i[68];
  assign data_o[67] = data_i[67];
  assign data_o[66] = data_i[66];
  assign data_o[65] = data_i[65];
  assign data_o[64] = data_i[64];
  assign data_o[63] = data_i[63];
  assign data_o[62] = data_i[62];
  assign data_o[61] = data_i[61];
  assign data_o[60] = data_i[60];
  assign data_o[59] = data_i[59];
  assign data_o[58] = data_i[58];
  assign data_o[57] = data_i[57];
  assign data_o[56] = data_i[56];
  assign data_o[55] = data_i[55];
  assign data_o[54] = data_i[54];
  assign data_o[53] = data_i[53];
  assign data_o[52] = data_i[52];
  assign data_o[51] = data_i[51];
  assign data_o[50] = data_i[50];
  assign data_o[49] = data_i[49];
  assign data_o[48] = data_i[48];
  assign data_o[47] = data_i[47];
  assign data_o[46] = data_i[46];
  assign data_o[45] = data_i[45];
  assign data_o[44] = data_i[44];
  assign data_o[43] = data_i[43];
  assign data_o[42] = data_i[42];
  assign data_o[41] = data_i[41];
  assign data_o[40] = data_i[40];
  assign data_o[39] = data_i[39];
  assign data_o[38] = data_i[38];
  assign data_o[37] = data_i[37];
  assign data_o[36] = data_i[36];
  assign data_o[35] = data_i[35];
  assign data_o[34] = data_i[34];
  assign data_o[33] = data_i[33];
  assign data_o[32] = data_i[32];
  assign data_o[31] = data_i[31];
  assign data_o[30] = data_i[30];
  assign data_o[29] = data_i[29];
  assign data_o[28] = data_i[28];
  assign data_o[27] = data_i[27];
  assign data_o[26] = data_i[26];
  assign data_o[25] = data_i[25];
  assign data_o[24] = data_i[24];
  assign data_o[23] = data_i[23];
  assign data_o[22] = data_i[22];
  assign data_o[21] = data_i[21];
  assign data_o[20] = data_i[20];
  assign data_o[19] = data_i[19];
  assign data_o[18] = data_i[18];
  assign data_o[17] = data_i[17];
  assign data_o[16] = data_i[16];
  assign data_o[15] = data_i[15];
  assign data_o[14] = data_i[14];
  assign data_o[13] = data_i[13];
  assign data_o[12] = data_i[12];
  assign data_o[11] = data_i[11];
  assign data_o[10] = data_i[10];
  assign data_o[9] = data_i[9];
  assign data_o[8] = data_i[8];
  assign data_o[7] = data_i[7];
  assign data_o[6] = data_i[6];
  assign data_o[5] = data_i[5];
  assign data_o[4] = data_i[4];
  assign data_o[3] = data_i[3];
  assign data_o[2] = data_i[2];
  assign data_o[1] = data_i[1];
  assign data_o[0] = data_i[0];

endmodule



module bsg_dff_chain_width_p66_num_stages_p2
(
  clk_i,
  data_i,
  data_o
);

  input [65:0] data_i;
  output [65:0] data_o;
  input clk_i;
  wire [65:0] data_o;
  wire \chained.data_delayed_1__65_ ,\chained.data_delayed_1__64_ ,
  \chained.data_delayed_1__63_ ,\chained.data_delayed_1__62_ ,\chained.data_delayed_1__61_ ,
  \chained.data_delayed_1__60_ ,\chained.data_delayed_1__59_ ,\chained.data_delayed_1__58_ ,
  \chained.data_delayed_1__57_ ,\chained.data_delayed_1__56_ ,
  \chained.data_delayed_1__55_ ,\chained.data_delayed_1__54_ ,\chained.data_delayed_1__53_ ,
  \chained.data_delayed_1__52_ ,\chained.data_delayed_1__51_ ,\chained.data_delayed_1__50_ ,
  \chained.data_delayed_1__49_ ,\chained.data_delayed_1__48_ ,
  \chained.data_delayed_1__47_ ,\chained.data_delayed_1__46_ ,\chained.data_delayed_1__45_ ,
  \chained.data_delayed_1__44_ ,\chained.data_delayed_1__43_ ,\chained.data_delayed_1__42_ ,
  \chained.data_delayed_1__41_ ,\chained.data_delayed_1__40_ ,
  \chained.data_delayed_1__39_ ,\chained.data_delayed_1__38_ ,\chained.data_delayed_1__37_ ,
  \chained.data_delayed_1__36_ ,\chained.data_delayed_1__35_ ,\chained.data_delayed_1__34_ ,
  \chained.data_delayed_1__33_ ,\chained.data_delayed_1__32_ ,
  \chained.data_delayed_1__31_ ,\chained.data_delayed_1__30_ ,\chained.data_delayed_1__29_ ,
  \chained.data_delayed_1__28_ ,\chained.data_delayed_1__27_ ,\chained.data_delayed_1__26_ ,
  \chained.data_delayed_1__25_ ,\chained.data_delayed_1__24_ ,
  \chained.data_delayed_1__23_ ,\chained.data_delayed_1__22_ ,\chained.data_delayed_1__21_ ,
  \chained.data_delayed_1__20_ ,\chained.data_delayed_1__19_ ,\chained.data_delayed_1__18_ ,
  \chained.data_delayed_1__17_ ,\chained.data_delayed_1__16_ ,
  \chained.data_delayed_1__15_ ,\chained.data_delayed_1__14_ ,\chained.data_delayed_1__13_ ,
  \chained.data_delayed_1__12_ ,\chained.data_delayed_1__11_ ,\chained.data_delayed_1__10_ ,
  \chained.data_delayed_1__9_ ,\chained.data_delayed_1__8_ ,
  \chained.data_delayed_1__7_ ,\chained.data_delayed_1__6_ ,\chained.data_delayed_1__5_ ,
  \chained.data_delayed_1__4_ ,\chained.data_delayed_1__3_ ,\chained.data_delayed_1__2_ ,
  \chained.data_delayed_1__1_ ,\chained.data_delayed_1__0_ ;

  bsg_dff_width_p66
  \chained.genblk1_1_.ch_reg 
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .data_o({ \chained.data_delayed_1__65_ , \chained.data_delayed_1__64_ , \chained.data_delayed_1__63_ , \chained.data_delayed_1__62_ , \chained.data_delayed_1__61_ , \chained.data_delayed_1__60_ , \chained.data_delayed_1__59_ , \chained.data_delayed_1__58_ , \chained.data_delayed_1__57_ , \chained.data_delayed_1__56_ , \chained.data_delayed_1__55_ , \chained.data_delayed_1__54_ , \chained.data_delayed_1__53_ , \chained.data_delayed_1__52_ , \chained.data_delayed_1__51_ , \chained.data_delayed_1__50_ , \chained.data_delayed_1__49_ , \chained.data_delayed_1__48_ , \chained.data_delayed_1__47_ , \chained.data_delayed_1__46_ , \chained.data_delayed_1__45_ , \chained.data_delayed_1__44_ , \chained.data_delayed_1__43_ , \chained.data_delayed_1__42_ , \chained.data_delayed_1__41_ , \chained.data_delayed_1__40_ , \chained.data_delayed_1__39_ , \chained.data_delayed_1__38_ , \chained.data_delayed_1__37_ , \chained.data_delayed_1__36_ , \chained.data_delayed_1__35_ , \chained.data_delayed_1__34_ , \chained.data_delayed_1__33_ , \chained.data_delayed_1__32_ , \chained.data_delayed_1__31_ , \chained.data_delayed_1__30_ , \chained.data_delayed_1__29_ , \chained.data_delayed_1__28_ , \chained.data_delayed_1__27_ , \chained.data_delayed_1__26_ , \chained.data_delayed_1__25_ , \chained.data_delayed_1__24_ , \chained.data_delayed_1__23_ , \chained.data_delayed_1__22_ , \chained.data_delayed_1__21_ , \chained.data_delayed_1__20_ , \chained.data_delayed_1__19_ , \chained.data_delayed_1__18_ , \chained.data_delayed_1__17_ , \chained.data_delayed_1__16_ , \chained.data_delayed_1__15_ , \chained.data_delayed_1__14_ , \chained.data_delayed_1__13_ , \chained.data_delayed_1__12_ , \chained.data_delayed_1__11_ , \chained.data_delayed_1__10_ , \chained.data_delayed_1__9_ , \chained.data_delayed_1__8_ , \chained.data_delayed_1__7_ , \chained.data_delayed_1__6_ , \chained.data_delayed_1__5_ , \chained.data_delayed_1__4_ , \chained.data_delayed_1__3_ , \chained.data_delayed_1__2_ , \chained.data_delayed_1__1_ , \chained.data_delayed_1__0_  })
  );


  bsg_dff_width_p66
  \chained.genblk1_2_.ch_reg 
  (
    .clk_i(clk_i),
    .data_i({ \chained.data_delayed_1__65_ , \chained.data_delayed_1__64_ , \chained.data_delayed_1__63_ , \chained.data_delayed_1__62_ , \chained.data_delayed_1__61_ , \chained.data_delayed_1__60_ , \chained.data_delayed_1__59_ , \chained.data_delayed_1__58_ , \chained.data_delayed_1__57_ , \chained.data_delayed_1__56_ , \chained.data_delayed_1__55_ , \chained.data_delayed_1__54_ , \chained.data_delayed_1__53_ , \chained.data_delayed_1__52_ , \chained.data_delayed_1__51_ , \chained.data_delayed_1__50_ , \chained.data_delayed_1__49_ , \chained.data_delayed_1__48_ , \chained.data_delayed_1__47_ , \chained.data_delayed_1__46_ , \chained.data_delayed_1__45_ , \chained.data_delayed_1__44_ , \chained.data_delayed_1__43_ , \chained.data_delayed_1__42_ , \chained.data_delayed_1__41_ , \chained.data_delayed_1__40_ , \chained.data_delayed_1__39_ , \chained.data_delayed_1__38_ , \chained.data_delayed_1__37_ , \chained.data_delayed_1__36_ , \chained.data_delayed_1__35_ , \chained.data_delayed_1__34_ , \chained.data_delayed_1__33_ , \chained.data_delayed_1__32_ , \chained.data_delayed_1__31_ , \chained.data_delayed_1__30_ , \chained.data_delayed_1__29_ , \chained.data_delayed_1__28_ , \chained.data_delayed_1__27_ , \chained.data_delayed_1__26_ , \chained.data_delayed_1__25_ , \chained.data_delayed_1__24_ , \chained.data_delayed_1__23_ , \chained.data_delayed_1__22_ , \chained.data_delayed_1__21_ , \chained.data_delayed_1__20_ , \chained.data_delayed_1__19_ , \chained.data_delayed_1__18_ , \chained.data_delayed_1__17_ , \chained.data_delayed_1__16_ , \chained.data_delayed_1__15_ , \chained.data_delayed_1__14_ , \chained.data_delayed_1__13_ , \chained.data_delayed_1__12_ , \chained.data_delayed_1__11_ , \chained.data_delayed_1__10_ , \chained.data_delayed_1__9_ , \chained.data_delayed_1__8_ , \chained.data_delayed_1__7_ , \chained.data_delayed_1__6_ , \chained.data_delayed_1__5_ , \chained.data_delayed_1__4_ , \chained.data_delayed_1__3_ , \chained.data_delayed_1__2_ , \chained.data_delayed_1__1_ , \chained.data_delayed_1__0_  }),
    .data_o(data_o)
  );


endmodule



module bsg_dff_chain_width_p71_num_stages_p3
(
  clk_i,
  data_i,
  data_o
);

  input [70:0] data_i;
  output [70:0] data_o;
  input clk_i;
  wire [70:0] data_o;
  wire \chained.data_delayed_2__70_ ,\chained.data_delayed_2__69_ ,
  \chained.data_delayed_2__68_ ,\chained.data_delayed_2__67_ ,\chained.data_delayed_2__66_ ,
  \chained.data_delayed_2__65_ ,\chained.data_delayed_2__64_ ,\chained.data_delayed_2__63_ ,
  \chained.data_delayed_2__62_ ,\chained.data_delayed_2__61_ ,
  \chained.data_delayed_2__60_ ,\chained.data_delayed_2__59_ ,\chained.data_delayed_2__58_ ,
  \chained.data_delayed_2__57_ ,\chained.data_delayed_2__56_ ,\chained.data_delayed_2__55_ ,
  \chained.data_delayed_2__54_ ,\chained.data_delayed_2__53_ ,
  \chained.data_delayed_2__52_ ,\chained.data_delayed_2__51_ ,\chained.data_delayed_2__50_ ,
  \chained.data_delayed_2__49_ ,\chained.data_delayed_2__48_ ,\chained.data_delayed_2__47_ ,
  \chained.data_delayed_2__46_ ,\chained.data_delayed_2__45_ ,
  \chained.data_delayed_2__44_ ,\chained.data_delayed_2__43_ ,\chained.data_delayed_2__42_ ,
  \chained.data_delayed_2__41_ ,\chained.data_delayed_2__40_ ,\chained.data_delayed_2__39_ ,
  \chained.data_delayed_2__38_ ,\chained.data_delayed_2__37_ ,
  \chained.data_delayed_2__36_ ,\chained.data_delayed_2__35_ ,\chained.data_delayed_2__34_ ,
  \chained.data_delayed_2__33_ ,\chained.data_delayed_2__32_ ,\chained.data_delayed_2__31_ ,
  \chained.data_delayed_2__30_ ,\chained.data_delayed_2__29_ ,
  \chained.data_delayed_2__28_ ,\chained.data_delayed_2__27_ ,\chained.data_delayed_2__26_ ,
  \chained.data_delayed_2__25_ ,\chained.data_delayed_2__24_ ,\chained.data_delayed_2__23_ ,
  \chained.data_delayed_2__22_ ,\chained.data_delayed_2__21_ ,
  \chained.data_delayed_2__20_ ,\chained.data_delayed_2__19_ ,\chained.data_delayed_2__18_ ,
  \chained.data_delayed_2__17_ ,\chained.data_delayed_2__16_ ,\chained.data_delayed_2__15_ ,
  \chained.data_delayed_2__14_ ,\chained.data_delayed_2__13_ ,
  \chained.data_delayed_2__12_ ,\chained.data_delayed_2__11_ ,\chained.data_delayed_2__10_ ,
  \chained.data_delayed_2__9_ ,\chained.data_delayed_2__8_ ,\chained.data_delayed_2__7_ ,
  \chained.data_delayed_2__6_ ,\chained.data_delayed_2__5_ ,
  \chained.data_delayed_2__4_ ,\chained.data_delayed_2__3_ ,\chained.data_delayed_2__2_ ,
  \chained.data_delayed_2__1_ ,\chained.data_delayed_2__0_ ,\chained.data_delayed_1__70_ ,
  \chained.data_delayed_1__69_ ,\chained.data_delayed_1__68_ ,\chained.data_delayed_1__67_ ,
  \chained.data_delayed_1__66_ ,\chained.data_delayed_1__65_ ,
  \chained.data_delayed_1__64_ ,\chained.data_delayed_1__63_ ,\chained.data_delayed_1__62_ ,
  \chained.data_delayed_1__61_ ,\chained.data_delayed_1__60_ ,\chained.data_delayed_1__59_ ,
  \chained.data_delayed_1__58_ ,\chained.data_delayed_1__57_ ,
  \chained.data_delayed_1__56_ ,\chained.data_delayed_1__55_ ,\chained.data_delayed_1__54_ ,
  \chained.data_delayed_1__53_ ,\chained.data_delayed_1__52_ ,\chained.data_delayed_1__51_ ,
  \chained.data_delayed_1__50_ ,\chained.data_delayed_1__49_ ,
  \chained.data_delayed_1__48_ ,\chained.data_delayed_1__47_ ,\chained.data_delayed_1__46_ ,
  \chained.data_delayed_1__45_ ,\chained.data_delayed_1__44_ ,\chained.data_delayed_1__43_ ,
  \chained.data_delayed_1__42_ ,\chained.data_delayed_1__41_ ,
  \chained.data_delayed_1__40_ ,\chained.data_delayed_1__39_ ,\chained.data_delayed_1__38_ ,
  \chained.data_delayed_1__37_ ,\chained.data_delayed_1__36_ ,\chained.data_delayed_1__35_ ,
  \chained.data_delayed_1__34_ ,\chained.data_delayed_1__33_ ,
  \chained.data_delayed_1__32_ ,\chained.data_delayed_1__31_ ,\chained.data_delayed_1__30_ ,
  \chained.data_delayed_1__29_ ,\chained.data_delayed_1__28_ ,\chained.data_delayed_1__27_ ,
  \chained.data_delayed_1__26_ ,\chained.data_delayed_1__25_ ,
  \chained.data_delayed_1__24_ ,\chained.data_delayed_1__23_ ,\chained.data_delayed_1__22_ ,
  \chained.data_delayed_1__21_ ,\chained.data_delayed_1__20_ ,\chained.data_delayed_1__19_ ,
  \chained.data_delayed_1__18_ ,\chained.data_delayed_1__17_ ,
  \chained.data_delayed_1__16_ ,\chained.data_delayed_1__15_ ,\chained.data_delayed_1__14_ ,
  \chained.data_delayed_1__13_ ,\chained.data_delayed_1__12_ ,\chained.data_delayed_1__11_ ,
  \chained.data_delayed_1__10_ ,\chained.data_delayed_1__9_ ,
  \chained.data_delayed_1__8_ ,\chained.data_delayed_1__7_ ,\chained.data_delayed_1__6_ ,
  \chained.data_delayed_1__5_ ,\chained.data_delayed_1__4_ ,\chained.data_delayed_1__3_ ,
  \chained.data_delayed_1__2_ ,\chained.data_delayed_1__1_ ,\chained.data_delayed_1__0_ ;

  bsg_dff_width_p71
  \chained.genblk1_1_.ch_reg 
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .data_o({ \chained.data_delayed_1__70_ , \chained.data_delayed_1__69_ , \chained.data_delayed_1__68_ , \chained.data_delayed_1__67_ , \chained.data_delayed_1__66_ , \chained.data_delayed_1__65_ , \chained.data_delayed_1__64_ , \chained.data_delayed_1__63_ , \chained.data_delayed_1__62_ , \chained.data_delayed_1__61_ , \chained.data_delayed_1__60_ , \chained.data_delayed_1__59_ , \chained.data_delayed_1__58_ , \chained.data_delayed_1__57_ , \chained.data_delayed_1__56_ , \chained.data_delayed_1__55_ , \chained.data_delayed_1__54_ , \chained.data_delayed_1__53_ , \chained.data_delayed_1__52_ , \chained.data_delayed_1__51_ , \chained.data_delayed_1__50_ , \chained.data_delayed_1__49_ , \chained.data_delayed_1__48_ , \chained.data_delayed_1__47_ , \chained.data_delayed_1__46_ , \chained.data_delayed_1__45_ , \chained.data_delayed_1__44_ , \chained.data_delayed_1__43_ , \chained.data_delayed_1__42_ , \chained.data_delayed_1__41_ , \chained.data_delayed_1__40_ , \chained.data_delayed_1__39_ , \chained.data_delayed_1__38_ , \chained.data_delayed_1__37_ , \chained.data_delayed_1__36_ , \chained.data_delayed_1__35_ , \chained.data_delayed_1__34_ , \chained.data_delayed_1__33_ , \chained.data_delayed_1__32_ , \chained.data_delayed_1__31_ , \chained.data_delayed_1__30_ , \chained.data_delayed_1__29_ , \chained.data_delayed_1__28_ , \chained.data_delayed_1__27_ , \chained.data_delayed_1__26_ , \chained.data_delayed_1__25_ , \chained.data_delayed_1__24_ , \chained.data_delayed_1__23_ , \chained.data_delayed_1__22_ , \chained.data_delayed_1__21_ , \chained.data_delayed_1__20_ , \chained.data_delayed_1__19_ , \chained.data_delayed_1__18_ , \chained.data_delayed_1__17_ , \chained.data_delayed_1__16_ , \chained.data_delayed_1__15_ , \chained.data_delayed_1__14_ , \chained.data_delayed_1__13_ , \chained.data_delayed_1__12_ , \chained.data_delayed_1__11_ , \chained.data_delayed_1__10_ , \chained.data_delayed_1__9_ , \chained.data_delayed_1__8_ , \chained.data_delayed_1__7_ , \chained.data_delayed_1__6_ , \chained.data_delayed_1__5_ , \chained.data_delayed_1__4_ , \chained.data_delayed_1__3_ , \chained.data_delayed_1__2_ , \chained.data_delayed_1__1_ , \chained.data_delayed_1__0_  })
  );


  bsg_dff_width_p71
  \chained.genblk1_2_.ch_reg 
  (
    .clk_i(clk_i),
    .data_i({ \chained.data_delayed_1__70_ , \chained.data_delayed_1__69_ , \chained.data_delayed_1__68_ , \chained.data_delayed_1__67_ , \chained.data_delayed_1__66_ , \chained.data_delayed_1__65_ , \chained.data_delayed_1__64_ , \chained.data_delayed_1__63_ , \chained.data_delayed_1__62_ , \chained.data_delayed_1__61_ , \chained.data_delayed_1__60_ , \chained.data_delayed_1__59_ , \chained.data_delayed_1__58_ , \chained.data_delayed_1__57_ , \chained.data_delayed_1__56_ , \chained.data_delayed_1__55_ , \chained.data_delayed_1__54_ , \chained.data_delayed_1__53_ , \chained.data_delayed_1__52_ , \chained.data_delayed_1__51_ , \chained.data_delayed_1__50_ , \chained.data_delayed_1__49_ , \chained.data_delayed_1__48_ , \chained.data_delayed_1__47_ , \chained.data_delayed_1__46_ , \chained.data_delayed_1__45_ , \chained.data_delayed_1__44_ , \chained.data_delayed_1__43_ , \chained.data_delayed_1__42_ , \chained.data_delayed_1__41_ , \chained.data_delayed_1__40_ , \chained.data_delayed_1__39_ , \chained.data_delayed_1__38_ , \chained.data_delayed_1__37_ , \chained.data_delayed_1__36_ , \chained.data_delayed_1__35_ , \chained.data_delayed_1__34_ , \chained.data_delayed_1__33_ , \chained.data_delayed_1__32_ , \chained.data_delayed_1__31_ , \chained.data_delayed_1__30_ , \chained.data_delayed_1__29_ , \chained.data_delayed_1__28_ , \chained.data_delayed_1__27_ , \chained.data_delayed_1__26_ , \chained.data_delayed_1__25_ , \chained.data_delayed_1__24_ , \chained.data_delayed_1__23_ , \chained.data_delayed_1__22_ , \chained.data_delayed_1__21_ , \chained.data_delayed_1__20_ , \chained.data_delayed_1__19_ , \chained.data_delayed_1__18_ , \chained.data_delayed_1__17_ , \chained.data_delayed_1__16_ , \chained.data_delayed_1__15_ , \chained.data_delayed_1__14_ , \chained.data_delayed_1__13_ , \chained.data_delayed_1__12_ , \chained.data_delayed_1__11_ , \chained.data_delayed_1__10_ , \chained.data_delayed_1__9_ , \chained.data_delayed_1__8_ , \chained.data_delayed_1__7_ , \chained.data_delayed_1__6_ , \chained.data_delayed_1__5_ , \chained.data_delayed_1__4_ , \chained.data_delayed_1__3_ , \chained.data_delayed_1__2_ , \chained.data_delayed_1__1_ , \chained.data_delayed_1__0_  }),
    .data_o({ \chained.data_delayed_2__70_ , \chained.data_delayed_2__69_ , \chained.data_delayed_2__68_ , \chained.data_delayed_2__67_ , \chained.data_delayed_2__66_ , \chained.data_delayed_2__65_ , \chained.data_delayed_2__64_ , \chained.data_delayed_2__63_ , \chained.data_delayed_2__62_ , \chained.data_delayed_2__61_ , \chained.data_delayed_2__60_ , \chained.data_delayed_2__59_ , \chained.data_delayed_2__58_ , \chained.data_delayed_2__57_ , \chained.data_delayed_2__56_ , \chained.data_delayed_2__55_ , \chained.data_delayed_2__54_ , \chained.data_delayed_2__53_ , \chained.data_delayed_2__52_ , \chained.data_delayed_2__51_ , \chained.data_delayed_2__50_ , \chained.data_delayed_2__49_ , \chained.data_delayed_2__48_ , \chained.data_delayed_2__47_ , \chained.data_delayed_2__46_ , \chained.data_delayed_2__45_ , \chained.data_delayed_2__44_ , \chained.data_delayed_2__43_ , \chained.data_delayed_2__42_ , \chained.data_delayed_2__41_ , \chained.data_delayed_2__40_ , \chained.data_delayed_2__39_ , \chained.data_delayed_2__38_ , \chained.data_delayed_2__37_ , \chained.data_delayed_2__36_ , \chained.data_delayed_2__35_ , \chained.data_delayed_2__34_ , \chained.data_delayed_2__33_ , \chained.data_delayed_2__32_ , \chained.data_delayed_2__31_ , \chained.data_delayed_2__30_ , \chained.data_delayed_2__29_ , \chained.data_delayed_2__28_ , \chained.data_delayed_2__27_ , \chained.data_delayed_2__26_ , \chained.data_delayed_2__25_ , \chained.data_delayed_2__24_ , \chained.data_delayed_2__23_ , \chained.data_delayed_2__22_ , \chained.data_delayed_2__21_ , \chained.data_delayed_2__20_ , \chained.data_delayed_2__19_ , \chained.data_delayed_2__18_ , \chained.data_delayed_2__17_ , \chained.data_delayed_2__16_ , \chained.data_delayed_2__15_ , \chained.data_delayed_2__14_ , \chained.data_delayed_2__13_ , \chained.data_delayed_2__12_ , \chained.data_delayed_2__11_ , \chained.data_delayed_2__10_ , \chained.data_delayed_2__9_ , \chained.data_delayed_2__8_ , \chained.data_delayed_2__7_ , \chained.data_delayed_2__6_ , \chained.data_delayed_2__5_ , \chained.data_delayed_2__4_ , \chained.data_delayed_2__3_ , \chained.data_delayed_2__2_ , \chained.data_delayed_2__1_ , \chained.data_delayed_2__0_  })
  );


  bsg_dff_width_p71
  \chained.genblk1_3_.ch_reg 
  (
    .clk_i(clk_i),
    .data_i({ \chained.data_delayed_2__70_ , \chained.data_delayed_2__69_ , \chained.data_delayed_2__68_ , \chained.data_delayed_2__67_ , \chained.data_delayed_2__66_ , \chained.data_delayed_2__65_ , \chained.data_delayed_2__64_ , \chained.data_delayed_2__63_ , \chained.data_delayed_2__62_ , \chained.data_delayed_2__61_ , \chained.data_delayed_2__60_ , \chained.data_delayed_2__59_ , \chained.data_delayed_2__58_ , \chained.data_delayed_2__57_ , \chained.data_delayed_2__56_ , \chained.data_delayed_2__55_ , \chained.data_delayed_2__54_ , \chained.data_delayed_2__53_ , \chained.data_delayed_2__52_ , \chained.data_delayed_2__51_ , \chained.data_delayed_2__50_ , \chained.data_delayed_2__49_ , \chained.data_delayed_2__48_ , \chained.data_delayed_2__47_ , \chained.data_delayed_2__46_ , \chained.data_delayed_2__45_ , \chained.data_delayed_2__44_ , \chained.data_delayed_2__43_ , \chained.data_delayed_2__42_ , \chained.data_delayed_2__41_ , \chained.data_delayed_2__40_ , \chained.data_delayed_2__39_ , \chained.data_delayed_2__38_ , \chained.data_delayed_2__37_ , \chained.data_delayed_2__36_ , \chained.data_delayed_2__35_ , \chained.data_delayed_2__34_ , \chained.data_delayed_2__33_ , \chained.data_delayed_2__32_ , \chained.data_delayed_2__31_ , \chained.data_delayed_2__30_ , \chained.data_delayed_2__29_ , \chained.data_delayed_2__28_ , \chained.data_delayed_2__27_ , \chained.data_delayed_2__26_ , \chained.data_delayed_2__25_ , \chained.data_delayed_2__24_ , \chained.data_delayed_2__23_ , \chained.data_delayed_2__22_ , \chained.data_delayed_2__21_ , \chained.data_delayed_2__20_ , \chained.data_delayed_2__19_ , \chained.data_delayed_2__18_ , \chained.data_delayed_2__17_ , \chained.data_delayed_2__16_ , \chained.data_delayed_2__15_ , \chained.data_delayed_2__14_ , \chained.data_delayed_2__13_ , \chained.data_delayed_2__12_ , \chained.data_delayed_2__11_ , \chained.data_delayed_2__10_ , \chained.data_delayed_2__9_ , \chained.data_delayed_2__8_ , \chained.data_delayed_2__7_ , \chained.data_delayed_2__6_ , \chained.data_delayed_2__5_ , \chained.data_delayed_2__4_ , \chained.data_delayed_2__3_ , \chained.data_delayed_2__2_ , \chained.data_delayed_2__1_ , \chained.data_delayed_2__0_  }),
    .data_o(data_o)
  );


endmodule



module bsg_dff_chain_width_p1_num_stages_p3
(
  clk_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  wire [0:0] data_o;
  wire \chained.data_delayed_2__0_ ,\chained.data_delayed_1__0_ ;

  bsg_dff_width_p1
  \chained.genblk1_1_.ch_reg 
  (
    .clk_i(clk_i),
    .data_i(data_i[0]),
    .data_o(\chained.data_delayed_1__0_ )
  );


  bsg_dff_width_p1
  \chained.genblk1_2_.ch_reg 
  (
    .clk_i(clk_i),
    .data_i(\chained.data_delayed_1__0_ ),
    .data_o(\chained.data_delayed_2__0_ )
  );


  bsg_dff_width_p1
  \chained.genblk1_3_.ch_reg 
  (
    .clk_i(clk_i),
    .data_i(\chained.data_delayed_2__0_ ),
    .data_o(data_o[0])
  );


endmodule



module bp_be_pipe_fma_00
(
  clk_i,
  reset_i,
  reservation_i,
  flush_i,
  frm_dyn_i,
  imul_data_o,
  imul_v_o,
  fma_data_o,
  fma_v_o,
  fma_fflags_o_nv_,
  fma_fflags_o_dz_,
  fma_fflags_o_of_,
  fma_fflags_o_uf_,
  fma_fflags_o_nx_
);

  input [520:0] reservation_i;
  input [2:0] frm_dyn_i;
  output [65:0] imul_data_o;
  output [65:0] fma_data_o;
  input clk_i;
  input reset_i;
  input flush_i;
  output imul_v_o;
  output fma_v_o;
  output fma_fflags_o_nv_;
  output fma_fflags_o_dz_;
  output fma_fflags_o_of_;
  output fma_fflags_o_uf_;
  output fma_fflags_o_nx_;
  wire [65:0] imul_data_o,fma_data_o,ird_data_lo,frd_data_lo;
  wire imul_v_o,fma_v_o,fma_fflags_o_nv_,fma_fflags_o_dz_,fma_fflags_o_of_,
  fma_fflags_o_uf_,fma_fflags_o_nx_,N0,N1,N2,N3,N4,N5,is_faddsub_li,N6,N7,N8,N9,N10,N11,N12,
  N13,N14,N15,N16,N17,N18,negate_sign,N19,N20,N21,N22,N23,N24,N25,N26,N27,frd_tag_r,
  invalid_exc,invalid_exc_r,fflags_lo_nv_,fflags_lo_dz_,fflags_lo_of_,
  fflags_lo_uf_,fflags_lo_nx_,imul_v_li,fma_v_li,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75;
  wire [2:0] frm_li,fma_op_li,frm_r;
  wire [64:64] fma_zero;
  wire [64:0] fma_a_li,fma_b_li,fma_c_li;
  wire [1:0] ird_tag_r;
  wire [63:0] imul_out;
  wire [74:0] fma_raw_lo,fma_raw_r;

  bsg_dff_chain_width_p4_num_stages_p0
  fma_info_chain
  (
    .clk_i(clk_i),
    .data_i({ frm_li, reservation_i[403:403] }),
    .data_o({ frm_r, frd_tag_r })
  );


  bsg_dff_chain_width_p2_num_stages_p0
  mul_info_chain
  (
    .clk_i(clk_i),
    .data_i(reservation_i[402:401]),
    .data_o(ird_tag_r)
  );


  mulAddRecFNToRaw_expWidth11_sigWidth53_pipelineStages0_imulEn1
  fma
  (
    .clock(clk_i),
    .control(1'b1),
    .op(fma_op_li),
    .a(fma_a_li),
    .b(fma_b_li),
    .c(fma_c_li),
    .roundingMode(frm_li),
    .invalidExc(invalid_exc),
    .out_isNaN(fma_raw_lo[74]),
    .out_isInf(fma_raw_lo[73]),
    .out_isZero(fma_raw_lo[72]),
    .out_sign(fma_raw_lo[69]),
    .out_sExp(fma_raw_lo[68:56]),
    .out_sig(fma_raw_lo[55:0]),
    .out_imul(imul_out)
  );


  bp_be_int_box_00
  imul_box
  (
    .raw_i(imul_out),
    .tag_i(ird_tag_r),
    .unsigned_i(1'b0),
    .reg_o(ird_data_lo)
  );


  bsg_dff_chain_width_p76_num_stages_p0
  round_info_chain
  (
    .clk_i(clk_i),
    .data_i({ invalid_exc, fma_raw_lo }),
    .data_o({ invalid_exc_r, fma_raw_r })
  );


  bp_be_fp_rebox_00
  rebox
  (
    .raw_i(fma_raw_r),
    .tag_i(frd_tag_r),
    .frm_i(frm_r),
    .invalid_exc_i(invalid_exc_r),
    .infinite_exc_i(1'b0),
    .reg_o(frd_data_lo),
    .fflags_o({ fflags_lo_nv_, fflags_lo_dz_, fflags_lo_of_, fflags_lo_uf_, fflags_lo_nx_ })
  );


  bsg_dff_chain_width_p66_num_stages_p2
  imul_retiming_chain
  (
    .clk_i(clk_i),
    .data_i(ird_data_lo),
    .data_o(imul_data_o)
  );


  bsg_dff_chain_width_p71_num_stages_p3
  fma_retiming_chain
  (
    .clk_i(clk_i),
    .data_i({ fflags_lo_nv_, fflags_lo_dz_, fflags_lo_of_, fflags_lo_uf_, fflags_lo_nx_, frd_data_lo }),
    .data_o({ fma_fflags_o_nv_, fma_fflags_o_dz_, fma_fflags_o_of_, fma_fflags_o_uf_, fma_fflags_o_nx_, fma_data_o })
  );


  bsg_dff_chain_width_p1_num_stages_p2
  imul_v_chain
  (
    .clk_i(clk_i),
    .data_i(imul_v_li),
    .data_o(imul_v_o)
  );


  bsg_dff_chain_width_p1_num_stages_p3
  fma_v_chain
  (
    .clk_i(clk_i),
    .data_i(fma_v_li),
    .data_o(fma_v_o)
  );

  assign N28 = reservation_i[462] & reservation_i[463];
  assign N29 = reservation_i[461] & N28;
  assign N30 = ~reservation_i[406];
  assign N31 = ~reservation_i[405];
  assign N32 = reservation_i[408] | reservation_i[409];
  assign N33 = reservation_i[407] | N32;
  assign N34 = N30 | N33;
  assign N35 = N31 | N34;
  assign N36 = reservation_i[404] | N35;
  assign N37 = ~N36;
  assign N38 = ~reservation_i[404];
  assign N39 = reservation_i[408] | reservation_i[409];
  assign N40 = reservation_i[407] | N39;
  assign N41 = N30 | N40;
  assign N42 = reservation_i[405] | N41;
  assign N43 = N38 | N42;
  assign N44 = ~N43;
  assign N45 = reservation_i[408] | reservation_i[409];
  assign N46 = reservation_i[407] | N45;
  assign N47 = N30 | N46;
  assign N48 = reservation_i[405] | N47;
  assign N49 = reservation_i[404] | N48;
  assign N50 = ~N49;
  assign N51 = reservation_i[408] | reservation_i[409];
  assign N52 = reservation_i[407] | N51;
  assign N53 = reservation_i[406] | N52;
  assign N54 = reservation_i[405] | N53;
  assign N55 = N38 | N54;
  assign N56 = ~N55;
  assign N57 = reservation_i[408] | reservation_i[409];
  assign N58 = reservation_i[407] | N57;
  assign N59 = reservation_i[406] | N58;
  assign N60 = N31 | N59;
  assign N61 = N38 | N60;
  assign N62 = ~N61;
  assign N63 = reservation_i[408] | reservation_i[409];
  assign N64 = reservation_i[407] | N63;
  assign N65 = reservation_i[406] | N64;
  assign N66 = reservation_i[405] | N65;
  assign N67 = reservation_i[404] | N66;
  assign N68 = ~N67;
  assign N69 = reservation_i[408] | reservation_i[409];
  assign N70 = reservation_i[407] | N69;
  assign N71 = reservation_i[406] | N70;
  assign N72 = N31 | N71;
  assign N73 = reservation_i[404] | N72;
  assign N74 = ~N73;
  assign frm_li = (N0)? frm_dyn_i : 
                  (N5)? reservation_i[463:461] : 1'b0;
  assign N0 = N29;
  assign fma_op_li = (N1)? { 1'b0, 1'b0, 1'b0 } : 
                     (N13)? { 1'b0, 1'b0, 1'b1 } : 
                     (N16)? { 1'b0, 1'b1, 1'b0 } : 
                     (N18)? { 1'b0, 1'b1, 1'b1 } : 
                     (N11)? { 1'b1, 1'b0, 1'b0 } : 1'b0;
  assign N1 = N6;
  assign fma_a_li = (N2)? { 1'b0, reservation_i[388:325] } : 
                    (N19)? reservation_i[194:130] : 1'b0;
  assign N2 = reservation_i[440];
  assign fma_b_li = (N3)? { 1'b0, reservation_i[323:260] } : 
                    (N23)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                    (N21)? reservation_i[129:65] : 1'b0;
  assign N3 = reservation_i[439];
  assign fma_c_li = (N4)? reservation_i[129:65] : 
                    (N27)? { fma_zero[64:64], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                    (N25)? reservation_i[64:0] : 1'b0;
  assign N4 = is_faddsub_li;
  assign N5 = ~N29;
  assign is_faddsub_li = N68 | N56;
  assign N6 = N75 | N74;
  assign N75 = N62 | N68;
  assign N7 = N50 | N56;
  assign N8 = N7 | N6;
  assign N9 = N44 | N8;
  assign N10 = N37 | N9;
  assign N11 = ~N10;
  assign N12 = ~N6;
  assign N13 = N7 & N12;
  assign N14 = ~N7;
  assign N15 = N12 & N14;
  assign N16 = N44 & N15;
  assign N17 = N15 & N43;
  assign N18 = N37 & N17;
  assign negate_sign = reservation_i[194] ^ reservation_i[129];
  assign fma_zero[64] = negate_sign;
  assign N19 = ~reservation_i[440];
  assign N20 = is_faddsub_li | reservation_i[439];
  assign N21 = ~N20;
  assign N22 = ~reservation_i[439];
  assign N23 = is_faddsub_li & N22;
  assign N24 = N74 | is_faddsub_li;
  assign N25 = ~N24;
  assign N26 = ~is_faddsub_li;
  assign N27 = N74 & N26;
  assign imul_v_li = reservation_i[520] & reservation_i[443];
  assign fma_v_li = reservation_i[520] & reservation_i[442];

endmodule



module bsg_imul_iterative_width_p64
(
  clk_i,
  reset_i,
  v_i,
  ready_and_o,
  opA_i,
  signed_opA_i,
  opB_i,
  signed_opB_i,
  gets_high_part_i,
  v_o,
  result_o,
  yumi_i
);

  input [63:0] opA_i;
  input [63:0] opB_i;
  output [63:0] result_o;
  input clk_i;
  input reset_i;
  input v_i;
  input signed_opA_i;
  input signed_opB_i;
  input gets_high_part_i;
  input yumi_i;
  output ready_and_o;
  output v_o;
  wire [63:0] result_o,opA_r,adder_a,opB_r,adder_b;
  wire ready_and_o,v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,
  N18,N19,N20,N21,N22,N23,N24,N25,gets_high_part_r,N26,shift_counter_full,N27,N28,
  N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,
  N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,
  N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,
  N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,
  N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,
  N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,
  N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,
  N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,
  N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
  N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,
  N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,
  N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,
  N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,
  N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,adder_neg_op,
  N265,latch_input,signed_opA,signed_opB,signed_opA_r,signed_opB_r,
  need_neg_result_r,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,
  N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,
  N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,
  N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,
  N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,
  N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,
  N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,
  N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,
  N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
  N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,
  N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,
  N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,
  N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,
  N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,
  N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,
  N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,
  N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,
  shifted_lsb,all_sh_lsb_zero_r,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,
  N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,
  N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,
  N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,
  N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,
  N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,
  N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,
  N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,
  N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,
  N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,
  N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,
  N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,
  N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,
  N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,
  N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,
  N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,
  N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,
  N803,N804,N805,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,
  N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,
  N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,
  N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N863,N864,N865,N866,N867,N868,
  N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,
  N885,N886;
  wire [6:0] shift_counter_r;
  wire [2:0] curr_state_r,next_state;
  wire [64:0] adder_result;
  reg curr_state_r_2_sv2v_reg,curr_state_r_1_sv2v_reg,curr_state_r_0_sv2v_reg,
  shift_counter_r_6_sv2v_reg,shift_counter_r_5_sv2v_reg,shift_counter_r_4_sv2v_reg,
  shift_counter_r_3_sv2v_reg,shift_counter_r_2_sv2v_reg,shift_counter_r_1_sv2v_reg,
  shift_counter_r_0_sv2v_reg,signed_opA_r_sv2v_reg,signed_opB_r_sv2v_reg,
  need_neg_result_r_sv2v_reg,gets_high_part_r_sv2v_reg,opA_r_63_sv2v_reg,opA_r_62_sv2v_reg,
  opA_r_61_sv2v_reg,opA_r_60_sv2v_reg,opA_r_59_sv2v_reg,opA_r_58_sv2v_reg,
  opA_r_57_sv2v_reg,opA_r_56_sv2v_reg,opA_r_55_sv2v_reg,opA_r_54_sv2v_reg,opA_r_53_sv2v_reg,
  opA_r_52_sv2v_reg,opA_r_51_sv2v_reg,opA_r_50_sv2v_reg,opA_r_49_sv2v_reg,
  opA_r_48_sv2v_reg,opA_r_47_sv2v_reg,opA_r_46_sv2v_reg,opA_r_45_sv2v_reg,opA_r_44_sv2v_reg,
  opA_r_43_sv2v_reg,opA_r_42_sv2v_reg,opA_r_41_sv2v_reg,opA_r_40_sv2v_reg,
  opA_r_39_sv2v_reg,opA_r_38_sv2v_reg,opA_r_37_sv2v_reg,opA_r_36_sv2v_reg,opA_r_35_sv2v_reg,
  opA_r_34_sv2v_reg,opA_r_33_sv2v_reg,opA_r_32_sv2v_reg,opA_r_31_sv2v_reg,
  opA_r_30_sv2v_reg,opA_r_29_sv2v_reg,opA_r_28_sv2v_reg,opA_r_27_sv2v_reg,
  opA_r_26_sv2v_reg,opA_r_25_sv2v_reg,opA_r_24_sv2v_reg,opA_r_23_sv2v_reg,opA_r_22_sv2v_reg,
  opA_r_21_sv2v_reg,opA_r_20_sv2v_reg,opA_r_19_sv2v_reg,opA_r_18_sv2v_reg,
  opA_r_17_sv2v_reg,opA_r_16_sv2v_reg,opA_r_15_sv2v_reg,opA_r_14_sv2v_reg,opA_r_13_sv2v_reg,
  opA_r_12_sv2v_reg,opA_r_11_sv2v_reg,opA_r_10_sv2v_reg,opA_r_9_sv2v_reg,
  opA_r_8_sv2v_reg,opA_r_7_sv2v_reg,opA_r_6_sv2v_reg,opA_r_5_sv2v_reg,opA_r_4_sv2v_reg,
  opA_r_3_sv2v_reg,opA_r_2_sv2v_reg,opA_r_1_sv2v_reg,opA_r_0_sv2v_reg,opB_r_63_sv2v_reg,
  opB_r_62_sv2v_reg,opB_r_61_sv2v_reg,opB_r_60_sv2v_reg,opB_r_59_sv2v_reg,
  opB_r_58_sv2v_reg,opB_r_57_sv2v_reg,opB_r_56_sv2v_reg,opB_r_55_sv2v_reg,opB_r_54_sv2v_reg,
  opB_r_53_sv2v_reg,opB_r_52_sv2v_reg,opB_r_51_sv2v_reg,opB_r_50_sv2v_reg,
  opB_r_49_sv2v_reg,opB_r_48_sv2v_reg,opB_r_47_sv2v_reg,opB_r_46_sv2v_reg,
  opB_r_45_sv2v_reg,opB_r_44_sv2v_reg,opB_r_43_sv2v_reg,opB_r_42_sv2v_reg,opB_r_41_sv2v_reg,
  opB_r_40_sv2v_reg,opB_r_39_sv2v_reg,opB_r_38_sv2v_reg,opB_r_37_sv2v_reg,
  opB_r_36_sv2v_reg,opB_r_35_sv2v_reg,opB_r_34_sv2v_reg,opB_r_33_sv2v_reg,opB_r_32_sv2v_reg,
  opB_r_31_sv2v_reg,opB_r_30_sv2v_reg,opB_r_29_sv2v_reg,opB_r_28_sv2v_reg,
  opB_r_27_sv2v_reg,opB_r_26_sv2v_reg,opB_r_25_sv2v_reg,opB_r_24_sv2v_reg,opB_r_23_sv2v_reg,
  opB_r_22_sv2v_reg,opB_r_21_sv2v_reg,opB_r_20_sv2v_reg,opB_r_19_sv2v_reg,
  opB_r_18_sv2v_reg,opB_r_17_sv2v_reg,opB_r_16_sv2v_reg,opB_r_15_sv2v_reg,opB_r_14_sv2v_reg,
  opB_r_13_sv2v_reg,opB_r_12_sv2v_reg,opB_r_11_sv2v_reg,opB_r_10_sv2v_reg,
  opB_r_9_sv2v_reg,opB_r_8_sv2v_reg,opB_r_7_sv2v_reg,opB_r_6_sv2v_reg,opB_r_5_sv2v_reg,
  opB_r_4_sv2v_reg,opB_r_3_sv2v_reg,opB_r_2_sv2v_reg,opB_r_1_sv2v_reg,
  opB_r_0_sv2v_reg,all_sh_lsb_zero_r_sv2v_reg,result_o_63_sv2v_reg,result_o_62_sv2v_reg,
  result_o_61_sv2v_reg,result_o_60_sv2v_reg,result_o_59_sv2v_reg,result_o_58_sv2v_reg,
  result_o_57_sv2v_reg,result_o_56_sv2v_reg,result_o_55_sv2v_reg,result_o_54_sv2v_reg,
  result_o_53_sv2v_reg,result_o_52_sv2v_reg,result_o_51_sv2v_reg,
  result_o_50_sv2v_reg,result_o_49_sv2v_reg,result_o_48_sv2v_reg,result_o_47_sv2v_reg,
  result_o_46_sv2v_reg,result_o_45_sv2v_reg,result_o_44_sv2v_reg,result_o_43_sv2v_reg,
  result_o_42_sv2v_reg,result_o_41_sv2v_reg,result_o_40_sv2v_reg,result_o_39_sv2v_reg,
  result_o_38_sv2v_reg,result_o_37_sv2v_reg,result_o_36_sv2v_reg,result_o_35_sv2v_reg,
  result_o_34_sv2v_reg,result_o_33_sv2v_reg,result_o_32_sv2v_reg,
  result_o_31_sv2v_reg,result_o_30_sv2v_reg,result_o_29_sv2v_reg,result_o_28_sv2v_reg,
  result_o_27_sv2v_reg,result_o_26_sv2v_reg,result_o_25_sv2v_reg,result_o_24_sv2v_reg,
  result_o_23_sv2v_reg,result_o_22_sv2v_reg,result_o_21_sv2v_reg,result_o_20_sv2v_reg,
  result_o_19_sv2v_reg,result_o_18_sv2v_reg,result_o_17_sv2v_reg,result_o_16_sv2v_reg,
  result_o_15_sv2v_reg,result_o_14_sv2v_reg,result_o_13_sv2v_reg,
  result_o_12_sv2v_reg,result_o_11_sv2v_reg,result_o_10_sv2v_reg,result_o_9_sv2v_reg,
  result_o_8_sv2v_reg,result_o_7_sv2v_reg,result_o_6_sv2v_reg,result_o_5_sv2v_reg,
  result_o_4_sv2v_reg,result_o_3_sv2v_reg,result_o_2_sv2v_reg,result_o_1_sv2v_reg,
  result_o_0_sv2v_reg;
  assign curr_state_r[2] = curr_state_r_2_sv2v_reg;
  assign curr_state_r[1] = curr_state_r_1_sv2v_reg;
  assign curr_state_r[0] = curr_state_r_0_sv2v_reg;
  assign shift_counter_r[6] = shift_counter_r_6_sv2v_reg;
  assign shift_counter_r[5] = shift_counter_r_5_sv2v_reg;
  assign shift_counter_r[4] = shift_counter_r_4_sv2v_reg;
  assign shift_counter_r[3] = shift_counter_r_3_sv2v_reg;
  assign shift_counter_r[2] = shift_counter_r_2_sv2v_reg;
  assign shift_counter_r[1] = shift_counter_r_1_sv2v_reg;
  assign shift_counter_r[0] = shift_counter_r_0_sv2v_reg;
  assign signed_opA_r = signed_opA_r_sv2v_reg;
  assign signed_opB_r = signed_opB_r_sv2v_reg;
  assign need_neg_result_r = need_neg_result_r_sv2v_reg;
  assign gets_high_part_r = gets_high_part_r_sv2v_reg;
  assign opA_r[63] = opA_r_63_sv2v_reg;
  assign opA_r[62] = opA_r_62_sv2v_reg;
  assign opA_r[61] = opA_r_61_sv2v_reg;
  assign opA_r[60] = opA_r_60_sv2v_reg;
  assign opA_r[59] = opA_r_59_sv2v_reg;
  assign opA_r[58] = opA_r_58_sv2v_reg;
  assign opA_r[57] = opA_r_57_sv2v_reg;
  assign opA_r[56] = opA_r_56_sv2v_reg;
  assign opA_r[55] = opA_r_55_sv2v_reg;
  assign opA_r[54] = opA_r_54_sv2v_reg;
  assign opA_r[53] = opA_r_53_sv2v_reg;
  assign opA_r[52] = opA_r_52_sv2v_reg;
  assign opA_r[51] = opA_r_51_sv2v_reg;
  assign opA_r[50] = opA_r_50_sv2v_reg;
  assign opA_r[49] = opA_r_49_sv2v_reg;
  assign opA_r[48] = opA_r_48_sv2v_reg;
  assign opA_r[47] = opA_r_47_sv2v_reg;
  assign opA_r[46] = opA_r_46_sv2v_reg;
  assign opA_r[45] = opA_r_45_sv2v_reg;
  assign opA_r[44] = opA_r_44_sv2v_reg;
  assign opA_r[43] = opA_r_43_sv2v_reg;
  assign opA_r[42] = opA_r_42_sv2v_reg;
  assign opA_r[41] = opA_r_41_sv2v_reg;
  assign opA_r[40] = opA_r_40_sv2v_reg;
  assign opA_r[39] = opA_r_39_sv2v_reg;
  assign opA_r[38] = opA_r_38_sv2v_reg;
  assign opA_r[37] = opA_r_37_sv2v_reg;
  assign opA_r[36] = opA_r_36_sv2v_reg;
  assign opA_r[35] = opA_r_35_sv2v_reg;
  assign opA_r[34] = opA_r_34_sv2v_reg;
  assign opA_r[33] = opA_r_33_sv2v_reg;
  assign opA_r[32] = opA_r_32_sv2v_reg;
  assign opA_r[31] = opA_r_31_sv2v_reg;
  assign opA_r[30] = opA_r_30_sv2v_reg;
  assign opA_r[29] = opA_r_29_sv2v_reg;
  assign opA_r[28] = opA_r_28_sv2v_reg;
  assign opA_r[27] = opA_r_27_sv2v_reg;
  assign opA_r[26] = opA_r_26_sv2v_reg;
  assign opA_r[25] = opA_r_25_sv2v_reg;
  assign opA_r[24] = opA_r_24_sv2v_reg;
  assign opA_r[23] = opA_r_23_sv2v_reg;
  assign opA_r[22] = opA_r_22_sv2v_reg;
  assign opA_r[21] = opA_r_21_sv2v_reg;
  assign opA_r[20] = opA_r_20_sv2v_reg;
  assign opA_r[19] = opA_r_19_sv2v_reg;
  assign opA_r[18] = opA_r_18_sv2v_reg;
  assign opA_r[17] = opA_r_17_sv2v_reg;
  assign opA_r[16] = opA_r_16_sv2v_reg;
  assign opA_r[15] = opA_r_15_sv2v_reg;
  assign opA_r[14] = opA_r_14_sv2v_reg;
  assign opA_r[13] = opA_r_13_sv2v_reg;
  assign opA_r[12] = opA_r_12_sv2v_reg;
  assign opA_r[11] = opA_r_11_sv2v_reg;
  assign opA_r[10] = opA_r_10_sv2v_reg;
  assign opA_r[9] = opA_r_9_sv2v_reg;
  assign opA_r[8] = opA_r_8_sv2v_reg;
  assign opA_r[7] = opA_r_7_sv2v_reg;
  assign opA_r[6] = opA_r_6_sv2v_reg;
  assign opA_r[5] = opA_r_5_sv2v_reg;
  assign opA_r[4] = opA_r_4_sv2v_reg;
  assign opA_r[3] = opA_r_3_sv2v_reg;
  assign opA_r[2] = opA_r_2_sv2v_reg;
  assign opA_r[1] = opA_r_1_sv2v_reg;
  assign opA_r[0] = opA_r_0_sv2v_reg;
  assign opB_r[63] = opB_r_63_sv2v_reg;
  assign opB_r[62] = opB_r_62_sv2v_reg;
  assign opB_r[61] = opB_r_61_sv2v_reg;
  assign opB_r[60] = opB_r_60_sv2v_reg;
  assign opB_r[59] = opB_r_59_sv2v_reg;
  assign opB_r[58] = opB_r_58_sv2v_reg;
  assign opB_r[57] = opB_r_57_sv2v_reg;
  assign opB_r[56] = opB_r_56_sv2v_reg;
  assign opB_r[55] = opB_r_55_sv2v_reg;
  assign opB_r[54] = opB_r_54_sv2v_reg;
  assign opB_r[53] = opB_r_53_sv2v_reg;
  assign opB_r[52] = opB_r_52_sv2v_reg;
  assign opB_r[51] = opB_r_51_sv2v_reg;
  assign opB_r[50] = opB_r_50_sv2v_reg;
  assign opB_r[49] = opB_r_49_sv2v_reg;
  assign opB_r[48] = opB_r_48_sv2v_reg;
  assign opB_r[47] = opB_r_47_sv2v_reg;
  assign opB_r[46] = opB_r_46_sv2v_reg;
  assign opB_r[45] = opB_r_45_sv2v_reg;
  assign opB_r[44] = opB_r_44_sv2v_reg;
  assign opB_r[43] = opB_r_43_sv2v_reg;
  assign opB_r[42] = opB_r_42_sv2v_reg;
  assign opB_r[41] = opB_r_41_sv2v_reg;
  assign opB_r[40] = opB_r_40_sv2v_reg;
  assign opB_r[39] = opB_r_39_sv2v_reg;
  assign opB_r[38] = opB_r_38_sv2v_reg;
  assign opB_r[37] = opB_r_37_sv2v_reg;
  assign opB_r[36] = opB_r_36_sv2v_reg;
  assign opB_r[35] = opB_r_35_sv2v_reg;
  assign opB_r[34] = opB_r_34_sv2v_reg;
  assign opB_r[33] = opB_r_33_sv2v_reg;
  assign opB_r[32] = opB_r_32_sv2v_reg;
  assign opB_r[31] = opB_r_31_sv2v_reg;
  assign opB_r[30] = opB_r_30_sv2v_reg;
  assign opB_r[29] = opB_r_29_sv2v_reg;
  assign opB_r[28] = opB_r_28_sv2v_reg;
  assign opB_r[27] = opB_r_27_sv2v_reg;
  assign opB_r[26] = opB_r_26_sv2v_reg;
  assign opB_r[25] = opB_r_25_sv2v_reg;
  assign opB_r[24] = opB_r_24_sv2v_reg;
  assign opB_r[23] = opB_r_23_sv2v_reg;
  assign opB_r[22] = opB_r_22_sv2v_reg;
  assign opB_r[21] = opB_r_21_sv2v_reg;
  assign opB_r[20] = opB_r_20_sv2v_reg;
  assign opB_r[19] = opB_r_19_sv2v_reg;
  assign opB_r[18] = opB_r_18_sv2v_reg;
  assign opB_r[17] = opB_r_17_sv2v_reg;
  assign opB_r[16] = opB_r_16_sv2v_reg;
  assign opB_r[15] = opB_r_15_sv2v_reg;
  assign opB_r[14] = opB_r_14_sv2v_reg;
  assign opB_r[13] = opB_r_13_sv2v_reg;
  assign opB_r[12] = opB_r_12_sv2v_reg;
  assign opB_r[11] = opB_r_11_sv2v_reg;
  assign opB_r[10] = opB_r_10_sv2v_reg;
  assign opB_r[9] = opB_r_9_sv2v_reg;
  assign opB_r[8] = opB_r_8_sv2v_reg;
  assign opB_r[7] = opB_r_7_sv2v_reg;
  assign opB_r[6] = opB_r_6_sv2v_reg;
  assign opB_r[5] = opB_r_5_sv2v_reg;
  assign opB_r[4] = opB_r_4_sv2v_reg;
  assign opB_r[3] = opB_r_3_sv2v_reg;
  assign opB_r[2] = opB_r_2_sv2v_reg;
  assign opB_r[1] = opB_r_1_sv2v_reg;
  assign opB_r[0] = opB_r_0_sv2v_reg;
  assign all_sh_lsb_zero_r = all_sh_lsb_zero_r_sv2v_reg;
  assign result_o[63] = result_o_63_sv2v_reg;
  assign result_o[62] = result_o_62_sv2v_reg;
  assign result_o[61] = result_o_61_sv2v_reg;
  assign result_o[60] = result_o_60_sv2v_reg;
  assign result_o[59] = result_o_59_sv2v_reg;
  assign result_o[58] = result_o_58_sv2v_reg;
  assign result_o[57] = result_o_57_sv2v_reg;
  assign result_o[56] = result_o_56_sv2v_reg;
  assign result_o[55] = result_o_55_sv2v_reg;
  assign result_o[54] = result_o_54_sv2v_reg;
  assign result_o[53] = result_o_53_sv2v_reg;
  assign result_o[52] = result_o_52_sv2v_reg;
  assign result_o[51] = result_o_51_sv2v_reg;
  assign result_o[50] = result_o_50_sv2v_reg;
  assign result_o[49] = result_o_49_sv2v_reg;
  assign result_o[48] = result_o_48_sv2v_reg;
  assign result_o[47] = result_o_47_sv2v_reg;
  assign result_o[46] = result_o_46_sv2v_reg;
  assign result_o[45] = result_o_45_sv2v_reg;
  assign result_o[44] = result_o_44_sv2v_reg;
  assign result_o[43] = result_o_43_sv2v_reg;
  assign result_o[42] = result_o_42_sv2v_reg;
  assign result_o[41] = result_o_41_sv2v_reg;
  assign result_o[40] = result_o_40_sv2v_reg;
  assign result_o[39] = result_o_39_sv2v_reg;
  assign result_o[38] = result_o_38_sv2v_reg;
  assign result_o[37] = result_o_37_sv2v_reg;
  assign result_o[36] = result_o_36_sv2v_reg;
  assign result_o[35] = result_o_35_sv2v_reg;
  assign result_o[34] = result_o_34_sv2v_reg;
  assign result_o[33] = result_o_33_sv2v_reg;
  assign result_o[32] = result_o_32_sv2v_reg;
  assign result_o[31] = result_o_31_sv2v_reg;
  assign result_o[30] = result_o_30_sv2v_reg;
  assign result_o[29] = result_o_29_sv2v_reg;
  assign result_o[28] = result_o_28_sv2v_reg;
  assign result_o[27] = result_o_27_sv2v_reg;
  assign result_o[26] = result_o_26_sv2v_reg;
  assign result_o[25] = result_o_25_sv2v_reg;
  assign result_o[24] = result_o_24_sv2v_reg;
  assign result_o[23] = result_o_23_sv2v_reg;
  assign result_o[22] = result_o_22_sv2v_reg;
  assign result_o[21] = result_o_21_sv2v_reg;
  assign result_o[20] = result_o_20_sv2v_reg;
  assign result_o[19] = result_o_19_sv2v_reg;
  assign result_o[18] = result_o_18_sv2v_reg;
  assign result_o[17] = result_o_17_sv2v_reg;
  assign result_o[16] = result_o_16_sv2v_reg;
  assign result_o[15] = result_o_15_sv2v_reg;
  assign result_o[14] = result_o_14_sv2v_reg;
  assign result_o[13] = result_o_13_sv2v_reg;
  assign result_o[12] = result_o_12_sv2v_reg;
  assign result_o[11] = result_o_11_sv2v_reg;
  assign result_o[10] = result_o_10_sv2v_reg;
  assign result_o[9] = result_o_9_sv2v_reg;
  assign result_o[8] = result_o_8_sv2v_reg;
  assign result_o[7] = result_o_7_sv2v_reg;
  assign result_o[6] = result_o_6_sv2v_reg;
  assign result_o[5] = result_o_5_sv2v_reg;
  assign result_o[4] = result_o_4_sv2v_reg;
  assign result_o[3] = result_o_3_sv2v_reg;
  assign result_o[2] = result_o_2_sv2v_reg;
  assign result_o[1] = result_o_1_sv2v_reg;
  assign result_o[0] = result_o_0_sv2v_reg;
  assign N27 = N802 & N807;
  assign N28 = N27 & N803;
  assign N29 = curr_state_r[2] | curr_state_r[1];
  assign N30 = N29 | N803;
  assign N32 = curr_state_r[2] | N807;
  assign N33 = N32 | curr_state_r[0];
  assign N35 = curr_state_r[2] | N807;
  assign N36 = N35 | N803;
  assign N38 = N802 | curr_state_r[1];
  assign N39 = N38 | curr_state_r[0];
  assign N41 = N802 | curr_state_r[1];
  assign N42 = N41 | N803;
  assign N44 = curr_state_r[2] & curr_state_r[1];
  assign N738 = reset_i | latch_input;
  assign N739 = reset_i | latch_input;
  assign N740 = reset_i | latch_input;
  assign N741 = reset_i | latch_input;
  assign N742 = reset_i | latch_input;
  assign N743 = reset_i | latch_input;
  assign N744 = reset_i | latch_input;
  assign N745 = reset_i | latch_input;
  assign N746 = reset_i | latch_input;
  assign N747 = reset_i | latch_input;
  assign N748 = reset_i | latch_input;
  assign N749 = reset_i | latch_input;
  assign N750 = reset_i | latch_input;
  assign N751 = reset_i | latch_input;
  assign N752 = reset_i | latch_input;
  assign N753 = reset_i | latch_input;
  assign N754 = reset_i | latch_input;
  assign N755 = reset_i | latch_input;
  assign N756 = reset_i | latch_input;
  assign N757 = reset_i | latch_input;
  assign N758 = reset_i | latch_input;
  assign N759 = reset_i | latch_input;
  assign N760 = reset_i | latch_input;
  assign N761 = reset_i | latch_input;
  assign N762 = reset_i | latch_input;
  assign N763 = reset_i | latch_input;
  assign N764 = reset_i | latch_input;
  assign N765 = reset_i | latch_input;
  assign N766 = reset_i | latch_input;
  assign N767 = reset_i | latch_input;
  assign N768 = reset_i | latch_input;
  assign N769 = reset_i | latch_input;
  assign N770 = reset_i | latch_input;
  assign N771 = reset_i | latch_input;
  assign N772 = reset_i | latch_input;
  assign N773 = reset_i | latch_input;
  assign N774 = reset_i | latch_input;
  assign N775 = reset_i | latch_input;
  assign N776 = reset_i | latch_input;
  assign N777 = reset_i | latch_input;
  assign N778 = reset_i | latch_input;
  assign N779 = reset_i | latch_input;
  assign N780 = reset_i | latch_input;
  assign N781 = reset_i | latch_input;
  assign N782 = reset_i | latch_input;
  assign N783 = reset_i | latch_input;
  assign N784 = reset_i | latch_input;
  assign N785 = reset_i | latch_input;
  assign N786 = reset_i | latch_input;
  assign N787 = reset_i | latch_input;
  assign N788 = reset_i | latch_input;
  assign N789 = reset_i | latch_input;
  assign N790 = reset_i | latch_input;
  assign N791 = reset_i | latch_input;
  assign N792 = reset_i | latch_input;
  assign N793 = reset_i | latch_input;
  assign N794 = reset_i | latch_input;
  assign N795 = reset_i | latch_input;
  assign N796 = reset_i | latch_input;
  assign N797 = reset_i | latch_input;
  assign N798 = reset_i | latch_input;
  assign N799 = reset_i | latch_input;
  assign N800 = reset_i | latch_input;
  assign N801 = reset_i | latch_input;
  assign N802 = ~curr_state_r[2];
  assign N803 = ~curr_state_r[0];
  assign N804 = curr_state_r[1] | N802;
  assign N805 = N803 | N804;
  assign v_o = ~N805;
  assign N807 = ~curr_state_r[1];
  assign N808 = N807 | curr_state_r[2];
  assign N809 = N803 | N808;
  assign N810 = ~N809;
  assign N811 = N807 | curr_state_r[2];
  assign N812 = N803 | N811;
  assign N813 = ~N812;
  assign N814 = N807 | curr_state_r[2];
  assign N815 = N803 | N814;
  assign N816 = ~N815;
  assign N817 = N807 | curr_state_r[2];
  assign N818 = N803 | N817;
  assign N819 = ~N818;
  assign N820 = curr_state_r[1] | curr_state_r[2];
  assign N821 = N803 | N820;
  assign N822 = ~N821;
  assign N823 = N807 | curr_state_r[2];
  assign N824 = N803 | N823;
  assign N825 = ~N824;
  assign N826 = N807 | curr_state_r[2];
  assign N827 = curr_state_r[0] | N826;
  assign N828 = ~N827;
  assign N829 = N807 | curr_state_r[2];
  assign N830 = N803 | N829;
  assign N831 = ~N830;
  assign N832 = curr_state_r[1] | N802;
  assign N833 = curr_state_r[0] | N832;
  assign N834 = ~N833;
  assign N835 = N807 | curr_state_r[2];
  assign N836 = N803 | N835;
  assign N837 = ~next_state[1];
  assign N838 = ~next_state[0];
  assign N839 = N837 | next_state[2];
  assign N840 = N838 | N839;
  assign N841 = ~N840;
  assign N842 = curr_state_r[1] | N802;
  assign N843 = curr_state_r[0] | N842;
  assign N844 = ~N843;
  assign N845 = curr_state_r[1] | curr_state_r[2];
  assign N846 = N803 | N845;
  assign N847 = ~N846;
  assign N848 = N807 | curr_state_r[2];
  assign N849 = curr_state_r[0] | N848;
  assign N850 = ~N849;
  assign N851 = curr_state_r[1] | N802;
  assign N852 = curr_state_r[0] | N851;
  assign N853 = ~N852;
  assign N854 = N807 | curr_state_r[2];
  assign N855 = curr_state_r[0] | N854;
  assign N856 = ~N855;
  assign N857 = curr_state_r[1] | curr_state_r[2];
  assign N858 = N803 | N857;
  assign N859 = ~N858;
  assign N860 = curr_state_r[1] | curr_state_r[2];
  assign N861 = curr_state_r[0] | N860;
  assign ready_and_o = ~N861;
  assign N863 = ~shift_counter_r[5];
  assign N864 = ~shift_counter_r[4];
  assign N865 = ~shift_counter_r[3];
  assign N866 = ~shift_counter_r[2];
  assign N867 = ~shift_counter_r[1];
  assign N868 = ~shift_counter_r[0];
  assign N869 = N863 | shift_counter_r[6];
  assign N870 = N864 | N869;
  assign N871 = N865 | N870;
  assign N872 = N866 | N871;
  assign N873 = N867 | N872;
  assign N874 = N868 | N873;
  assign N875 = ~N874;
  assign N876 = ~shift_counter_r[6];
  assign N877 = shift_counter_r[5] | N876;
  assign N878 = shift_counter_r[4] | N877;
  assign N879 = shift_counter_r[3] | N878;
  assign N880 = shift_counter_r[2] | N879;
  assign N881 = shift_counter_r[1] | N880;
  assign N882 = shift_counter_r[0] | N881;
  assign N883 = ~N882;
  assign adder_result = adder_a + adder_b;
  assign { N59, N58, N57, N56, N55, N54, N53 } = shift_counter_r + 1'b1;
  assign shift_counter_full = (N0)? N875 : 
                              (N1)? N883 : 1'b0;
  assign N0 = gets_high_part_r;
  assign N1 = N26;
  assign next_state = (N2)? { 1'b0, 1'b0, v_i } : 
                      (N3)? { 1'b0, 1'b1, 1'b0 } : 
                      (N4)? { 1'b0, 1'b1, 1'b1 } : 
                      (N5)? { shift_counter_full, N45, N45 } : 
                      (N6)? { 1'b1, 1'b0, 1'b1 } : 
                      (N7)? { N46, 1'b0, N46 } : 
                      (N8)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2 = N28;
  assign N3 = N31;
  assign N4 = N34;
  assign N5 = N37;
  assign N6 = N40;
  assign N7 = N43;
  assign N8 = N44;
  assign N60 = (N9)? 1'b1 : 
               (N69)? 1'b1 : 
               (N51)? 1'b0 : 1'b0;
  assign N9 = N49;
  assign { N67, N66, N65, N64, N63, N62, N61 } = (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                 (N69)? { N59, N58, N57, N56, N55, N54, N53 } : 1'b0;
  assign adder_a = (N10)? { N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136 } : 
                   (N11)? { N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200 } : 
                   (N12)? { N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264 } : 
                   (N72)? result_o : 1'b0;
  assign N10 = N859;
  assign N11 = N856;
  assign N12 = N844;
  assign adder_b = (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                   (N14)? opA_r : 1'b0;
  assign N13 = adder_neg_op;
  assign N14 = N265;
  assign N272 = (N15)? 1'b1 : 
                (N16)? 1'b1 : 
                (N271)? 1'b0 : 1'b0;
  assign N15 = N268;
  assign N16 = N269;
  assign { N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273 } = (N15)? { opA_r[62:0], 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N16)? adder_result[63:0] : 1'b0;
  assign N337 = (N17)? 1'b1 : 
                (N18)? N272 : 1'b0;
  assign N17 = latch_input;
  assign N18 = N267;
  assign { N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338 } = (N17)? opA_i : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N18)? { N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273 } : 1'b0;
  assign N405 = (N19)? 1'b1 : 
                (N20)? 1'b1 : 
                (N404)? 1'b0 : 1'b0;
  assign N19 = N813;
  assign N20 = N402;
  assign { N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406 } = (N19)? { 1'b0, opB_r[63:1] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N20)? adder_result[63:0] : 1'b0;
  assign N470 = (N17)? 1'b1 : 
                (N18)? N405 : 1'b0;
  assign { N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471 } = (N17)? opB_i : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N18)? { N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406 } : 1'b0;
  assign shifted_lsb = (N21)? adder_result[0] : 
                       (N535)? result_o[0] : 1'b0;
  assign N21 = opB_r[0];
  assign { N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545 } = (N22)? { N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N544)? adder_result[63:0] : 1'b0;
  assign N22 = N543;
  assign { N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609 } = (N0)? adder_result[64:1] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N1)? adder_result[63:0] : 1'b0;
  assign N673 = (N23)? 1'b1 : 
                (N24)? 1'b1 : 
                (N25)? gets_high_part_r : 
                (N542)? 1'b0 : 1'b0;
  assign N23 = N537;
  assign N24 = N538;
  assign N25 = N539;
  assign { N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674 } = (N23)? { N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N24)? { N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N25)? { 1'b0, result_o[63:1] } : 1'b0;
  assign N26 = ~gets_high_part_r;
  assign N31 = ~N30;
  assign N34 = ~N33;
  assign N37 = ~N36;
  assign N40 = ~N39;
  assign N43 = ~N42;
  assign N45 = ~shift_counter_full;
  assign N46 = ~yumi_i;
  assign N47 = ~reset_i;
  assign N48 = N47;
  assign N49 = N836 & N841;
  assign N50 = N819 | N49;
  assign N51 = ~N50;
  assign N52 = N48 & N69;
  assign N68 = ~N49;
  assign N69 = N819 & N68;
  assign N70 = N856 | N859;
  assign N71 = N844 | N70;
  assign N72 = ~N71;
  assign N73 = ~opA_r[63];
  assign N74 = ~opA_r[62];
  assign N75 = ~opA_r[61];
  assign N76 = ~opA_r[60];
  assign N77 = ~opA_r[59];
  assign N78 = ~opA_r[58];
  assign N79 = ~opA_r[57];
  assign N80 = ~opA_r[56];
  assign N81 = ~opA_r[55];
  assign N82 = ~opA_r[54];
  assign N83 = ~opA_r[53];
  assign N84 = ~opA_r[52];
  assign N85 = ~opA_r[51];
  assign N86 = ~opA_r[50];
  assign N87 = ~opA_r[49];
  assign N88 = ~opA_r[48];
  assign N89 = ~opA_r[47];
  assign N90 = ~opA_r[46];
  assign N91 = ~opA_r[45];
  assign N92 = ~opA_r[44];
  assign N93 = ~opA_r[43];
  assign N94 = ~opA_r[42];
  assign N95 = ~opA_r[41];
  assign N96 = ~opA_r[40];
  assign N97 = ~opA_r[39];
  assign N98 = ~opA_r[38];
  assign N99 = ~opA_r[37];
  assign N100 = ~opA_r[36];
  assign N101 = ~opA_r[35];
  assign N102 = ~opA_r[34];
  assign N103 = ~opA_r[33];
  assign N104 = ~opA_r[32];
  assign N105 = ~opA_r[31];
  assign N106 = ~opA_r[30];
  assign N107 = ~opA_r[29];
  assign N108 = ~opA_r[28];
  assign N109 = ~opA_r[27];
  assign N110 = ~opA_r[26];
  assign N111 = ~opA_r[25];
  assign N112 = ~opA_r[24];
  assign N113 = ~opA_r[23];
  assign N114 = ~opA_r[22];
  assign N115 = ~opA_r[21];
  assign N116 = ~opA_r[20];
  assign N117 = ~opA_r[19];
  assign N118 = ~opA_r[18];
  assign N119 = ~opA_r[17];
  assign N120 = ~opA_r[16];
  assign N121 = ~opA_r[15];
  assign N122 = ~opA_r[14];
  assign N123 = ~opA_r[13];
  assign N124 = ~opA_r[12];
  assign N125 = ~opA_r[11];
  assign N126 = ~opA_r[10];
  assign N127 = ~opA_r[9];
  assign N128 = ~opA_r[8];
  assign N129 = ~opA_r[7];
  assign N130 = ~opA_r[6];
  assign N131 = ~opA_r[5];
  assign N132 = ~opA_r[4];
  assign N133 = ~opA_r[3];
  assign N134 = ~opA_r[2];
  assign N135 = ~opA_r[1];
  assign N136 = ~opA_r[0];
  assign N137 = ~opB_r[63];
  assign N138 = ~opB_r[62];
  assign N139 = ~opB_r[61];
  assign N140 = ~opB_r[60];
  assign N141 = ~opB_r[59];
  assign N142 = ~opB_r[58];
  assign N143 = ~opB_r[57];
  assign N144 = ~opB_r[56];
  assign N145 = ~opB_r[55];
  assign N146 = ~opB_r[54];
  assign N147 = ~opB_r[53];
  assign N148 = ~opB_r[52];
  assign N149 = ~opB_r[51];
  assign N150 = ~opB_r[50];
  assign N151 = ~opB_r[49];
  assign N152 = ~opB_r[48];
  assign N153 = ~opB_r[47];
  assign N154 = ~opB_r[46];
  assign N155 = ~opB_r[45];
  assign N156 = ~opB_r[44];
  assign N157 = ~opB_r[43];
  assign N158 = ~opB_r[42];
  assign N159 = ~opB_r[41];
  assign N160 = ~opB_r[40];
  assign N161 = ~opB_r[39];
  assign N162 = ~opB_r[38];
  assign N163 = ~opB_r[37];
  assign N164 = ~opB_r[36];
  assign N165 = ~opB_r[35];
  assign N166 = ~opB_r[34];
  assign N167 = ~opB_r[33];
  assign N168 = ~opB_r[32];
  assign N169 = ~opB_r[31];
  assign N170 = ~opB_r[30];
  assign N171 = ~opB_r[29];
  assign N172 = ~opB_r[28];
  assign N173 = ~opB_r[27];
  assign N174 = ~opB_r[26];
  assign N175 = ~opB_r[25];
  assign N176 = ~opB_r[24];
  assign N177 = ~opB_r[23];
  assign N178 = ~opB_r[22];
  assign N179 = ~opB_r[21];
  assign N180 = ~opB_r[20];
  assign N181 = ~opB_r[19];
  assign N182 = ~opB_r[18];
  assign N183 = ~opB_r[17];
  assign N184 = ~opB_r[16];
  assign N185 = ~opB_r[15];
  assign N186 = ~opB_r[14];
  assign N187 = ~opB_r[13];
  assign N188 = ~opB_r[12];
  assign N189 = ~opB_r[11];
  assign N190 = ~opB_r[10];
  assign N191 = ~opB_r[9];
  assign N192 = ~opB_r[8];
  assign N193 = ~opB_r[7];
  assign N194 = ~opB_r[6];
  assign N195 = ~opB_r[5];
  assign N196 = ~opB_r[4];
  assign N197 = ~opB_r[3];
  assign N198 = ~opB_r[2];
  assign N199 = ~opB_r[1];
  assign N200 = ~opB_r[0];
  assign N201 = ~result_o[63];
  assign N202 = ~result_o[62];
  assign N203 = ~result_o[61];
  assign N204 = ~result_o[60];
  assign N205 = ~result_o[59];
  assign N206 = ~result_o[58];
  assign N207 = ~result_o[57];
  assign N208 = ~result_o[56];
  assign N209 = ~result_o[55];
  assign N210 = ~result_o[54];
  assign N211 = ~result_o[53];
  assign N212 = ~result_o[52];
  assign N213 = ~result_o[51];
  assign N214 = ~result_o[50];
  assign N215 = ~result_o[49];
  assign N216 = ~result_o[48];
  assign N217 = ~result_o[47];
  assign N218 = ~result_o[46];
  assign N219 = ~result_o[45];
  assign N220 = ~result_o[44];
  assign N221 = ~result_o[43];
  assign N222 = ~result_o[42];
  assign N223 = ~result_o[41];
  assign N224 = ~result_o[40];
  assign N225 = ~result_o[39];
  assign N226 = ~result_o[38];
  assign N227 = ~result_o[37];
  assign N228 = ~result_o[36];
  assign N229 = ~result_o[35];
  assign N230 = ~result_o[34];
  assign N231 = ~result_o[33];
  assign N232 = ~result_o[32];
  assign N233 = ~result_o[31];
  assign N234 = ~result_o[30];
  assign N235 = ~result_o[29];
  assign N236 = ~result_o[28];
  assign N237 = ~result_o[27];
  assign N238 = ~result_o[26];
  assign N239 = ~result_o[25];
  assign N240 = ~result_o[24];
  assign N241 = ~result_o[23];
  assign N242 = ~result_o[22];
  assign N243 = ~result_o[21];
  assign N244 = ~result_o[20];
  assign N245 = ~result_o[19];
  assign N246 = ~result_o[18];
  assign N247 = ~result_o[17];
  assign N248 = ~result_o[16];
  assign N249 = ~result_o[15];
  assign N250 = ~result_o[14];
  assign N251 = ~result_o[13];
  assign N252 = ~result_o[12];
  assign N253 = ~result_o[11];
  assign N254 = ~result_o[10];
  assign N255 = ~result_o[9];
  assign N256 = ~result_o[8];
  assign N257 = ~result_o[7];
  assign N258 = ~result_o[6];
  assign N259 = ~result_o[5];
  assign N260 = ~result_o[4];
  assign N261 = ~result_o[3];
  assign N262 = ~result_o[2];
  assign N263 = ~result_o[1];
  assign N264 = ~result_o[0];
  assign adder_neg_op = N884 | N853;
  assign N884 = N847 | N850;
  assign N265 = ~adder_neg_op;
  assign latch_input = v_i & ready_and_o;
  assign signed_opA = signed_opA_i & opA_i[63];
  assign signed_opB = signed_opB_i & opB_i[63];
  assign N266 = signed_opA ^ signed_opB;
  assign N267 = ~latch_input;
  assign N268 = N825 & N26;
  assign N269 = N822 & signed_opA_r;
  assign N270 = N269 | N268;
  assign N271 = ~N270;
  assign N402 = N828 & signed_opB_r;
  assign N403 = N402 | N813;
  assign N404 = ~N403;
  assign N535 = ~opB_r[0];
  assign N536 = all_sh_lsb_zero_r & N885;
  assign N885 = ~shifted_lsb;
  assign N537 = N834 & need_neg_result_r;
  assign N538 = N831 & opB_r[0];
  assign N539 = N816 & N200;
  assign N540 = N538 | N537;
  assign N541 = N539 | N540;
  assign N542 = ~N541;
  assign N543 = gets_high_part_r & N886;
  assign N886 = ~all_sh_lsb_zero_r;
  assign N544 = ~N543;

  always @(posedge clk_i) begin
    if(reset_i) begin
      curr_state_r_2_sv2v_reg <= 1'b0;
      curr_state_r_1_sv2v_reg <= 1'b0;
      curr_state_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      curr_state_r_2_sv2v_reg <= next_state[2];
      curr_state_r_1_sv2v_reg <= next_state[1];
      curr_state_r_0_sv2v_reg <= next_state[0];
    end 
    if(reset_i) begin
      shift_counter_r_6_sv2v_reg <= 1'b0;
      shift_counter_r_5_sv2v_reg <= 1'b0;
      shift_counter_r_4_sv2v_reg <= 1'b0;
      shift_counter_r_3_sv2v_reg <= 1'b0;
      shift_counter_r_2_sv2v_reg <= 1'b0;
      shift_counter_r_1_sv2v_reg <= 1'b0;
      shift_counter_r_0_sv2v_reg <= 1'b0;
    end else if(N60) begin
      shift_counter_r_6_sv2v_reg <= N67;
      shift_counter_r_5_sv2v_reg <= N66;
      shift_counter_r_4_sv2v_reg <= N65;
      shift_counter_r_3_sv2v_reg <= N64;
      shift_counter_r_2_sv2v_reg <= N63;
      shift_counter_r_1_sv2v_reg <= N62;
      shift_counter_r_0_sv2v_reg <= N61;
    end 
    if(reset_i) begin
      signed_opA_r_sv2v_reg <= 1'b0;
      signed_opB_r_sv2v_reg <= 1'b0;
      need_neg_result_r_sv2v_reg <= 1'b0;
      gets_high_part_r_sv2v_reg <= 1'b0;
    end else if(latch_input) begin
      signed_opA_r_sv2v_reg <= signed_opA;
      signed_opB_r_sv2v_reg <= signed_opB;
      need_neg_result_r_sv2v_reg <= N266;
      gets_high_part_r_sv2v_reg <= gets_high_part_i;
    end 
    if(reset_i) begin
      opA_r_63_sv2v_reg <= 1'b0;
      opA_r_62_sv2v_reg <= 1'b0;
      opA_r_61_sv2v_reg <= 1'b0;
      opA_r_60_sv2v_reg <= 1'b0;
      opA_r_59_sv2v_reg <= 1'b0;
      opA_r_58_sv2v_reg <= 1'b0;
      opA_r_57_sv2v_reg <= 1'b0;
      opA_r_56_sv2v_reg <= 1'b0;
      opA_r_55_sv2v_reg <= 1'b0;
      opA_r_54_sv2v_reg <= 1'b0;
      opA_r_53_sv2v_reg <= 1'b0;
      opA_r_52_sv2v_reg <= 1'b0;
      opA_r_51_sv2v_reg <= 1'b0;
      opA_r_50_sv2v_reg <= 1'b0;
      opA_r_49_sv2v_reg <= 1'b0;
      opA_r_48_sv2v_reg <= 1'b0;
      opA_r_47_sv2v_reg <= 1'b0;
      opA_r_46_sv2v_reg <= 1'b0;
      opA_r_45_sv2v_reg <= 1'b0;
      opA_r_44_sv2v_reg <= 1'b0;
      opA_r_43_sv2v_reg <= 1'b0;
      opA_r_42_sv2v_reg <= 1'b0;
      opA_r_41_sv2v_reg <= 1'b0;
      opA_r_40_sv2v_reg <= 1'b0;
      opA_r_39_sv2v_reg <= 1'b0;
      opA_r_38_sv2v_reg <= 1'b0;
      opA_r_37_sv2v_reg <= 1'b0;
      opA_r_36_sv2v_reg <= 1'b0;
      opA_r_35_sv2v_reg <= 1'b0;
      opA_r_34_sv2v_reg <= 1'b0;
      opA_r_33_sv2v_reg <= 1'b0;
      opA_r_32_sv2v_reg <= 1'b0;
      opA_r_31_sv2v_reg <= 1'b0;
      opA_r_30_sv2v_reg <= 1'b0;
      opA_r_29_sv2v_reg <= 1'b0;
      opA_r_28_sv2v_reg <= 1'b0;
      opA_r_27_sv2v_reg <= 1'b0;
      opA_r_26_sv2v_reg <= 1'b0;
      opA_r_25_sv2v_reg <= 1'b0;
      opA_r_24_sv2v_reg <= 1'b0;
      opA_r_23_sv2v_reg <= 1'b0;
      opA_r_22_sv2v_reg <= 1'b0;
      opA_r_21_sv2v_reg <= 1'b0;
      opA_r_20_sv2v_reg <= 1'b0;
      opA_r_19_sv2v_reg <= 1'b0;
      opA_r_18_sv2v_reg <= 1'b0;
      opA_r_17_sv2v_reg <= 1'b0;
      opA_r_16_sv2v_reg <= 1'b0;
      opA_r_15_sv2v_reg <= 1'b0;
      opA_r_14_sv2v_reg <= 1'b0;
      opA_r_13_sv2v_reg <= 1'b0;
      opA_r_12_sv2v_reg <= 1'b0;
      opA_r_11_sv2v_reg <= 1'b0;
      opA_r_10_sv2v_reg <= 1'b0;
      opA_r_9_sv2v_reg <= 1'b0;
      opA_r_8_sv2v_reg <= 1'b0;
      opA_r_7_sv2v_reg <= 1'b0;
      opA_r_6_sv2v_reg <= 1'b0;
      opA_r_5_sv2v_reg <= 1'b0;
      opA_r_4_sv2v_reg <= 1'b0;
      opA_r_3_sv2v_reg <= 1'b0;
      opA_r_2_sv2v_reg <= 1'b0;
      opA_r_1_sv2v_reg <= 1'b0;
      opA_r_0_sv2v_reg <= 1'b0;
    end else if(N337) begin
      opA_r_63_sv2v_reg <= N401;
      opA_r_62_sv2v_reg <= N400;
      opA_r_61_sv2v_reg <= N399;
      opA_r_60_sv2v_reg <= N398;
      opA_r_59_sv2v_reg <= N397;
      opA_r_58_sv2v_reg <= N396;
      opA_r_57_sv2v_reg <= N395;
      opA_r_56_sv2v_reg <= N394;
      opA_r_55_sv2v_reg <= N393;
      opA_r_54_sv2v_reg <= N392;
      opA_r_53_sv2v_reg <= N391;
      opA_r_52_sv2v_reg <= N390;
      opA_r_51_sv2v_reg <= N389;
      opA_r_50_sv2v_reg <= N388;
      opA_r_49_sv2v_reg <= N387;
      opA_r_48_sv2v_reg <= N386;
      opA_r_47_sv2v_reg <= N385;
      opA_r_46_sv2v_reg <= N384;
      opA_r_45_sv2v_reg <= N383;
      opA_r_44_sv2v_reg <= N382;
      opA_r_43_sv2v_reg <= N381;
      opA_r_42_sv2v_reg <= N380;
      opA_r_41_sv2v_reg <= N379;
      opA_r_40_sv2v_reg <= N378;
      opA_r_39_sv2v_reg <= N377;
      opA_r_38_sv2v_reg <= N376;
      opA_r_37_sv2v_reg <= N375;
      opA_r_36_sv2v_reg <= N374;
      opA_r_35_sv2v_reg <= N373;
      opA_r_34_sv2v_reg <= N372;
      opA_r_33_sv2v_reg <= N371;
      opA_r_32_sv2v_reg <= N370;
      opA_r_31_sv2v_reg <= N369;
      opA_r_30_sv2v_reg <= N368;
      opA_r_29_sv2v_reg <= N367;
      opA_r_28_sv2v_reg <= N366;
      opA_r_27_sv2v_reg <= N365;
      opA_r_26_sv2v_reg <= N364;
      opA_r_25_sv2v_reg <= N363;
      opA_r_24_sv2v_reg <= N362;
      opA_r_23_sv2v_reg <= N361;
      opA_r_22_sv2v_reg <= N360;
      opA_r_21_sv2v_reg <= N359;
      opA_r_20_sv2v_reg <= N358;
      opA_r_19_sv2v_reg <= N357;
      opA_r_18_sv2v_reg <= N356;
      opA_r_17_sv2v_reg <= N355;
      opA_r_16_sv2v_reg <= N354;
      opA_r_15_sv2v_reg <= N353;
      opA_r_14_sv2v_reg <= N352;
      opA_r_13_sv2v_reg <= N351;
      opA_r_12_sv2v_reg <= N350;
      opA_r_11_sv2v_reg <= N349;
      opA_r_10_sv2v_reg <= N348;
      opA_r_9_sv2v_reg <= N347;
      opA_r_8_sv2v_reg <= N346;
      opA_r_7_sv2v_reg <= N345;
      opA_r_6_sv2v_reg <= N344;
      opA_r_5_sv2v_reg <= N343;
      opA_r_4_sv2v_reg <= N342;
      opA_r_3_sv2v_reg <= N341;
      opA_r_2_sv2v_reg <= N340;
      opA_r_1_sv2v_reg <= N339;
      opA_r_0_sv2v_reg <= N338;
    end 
    if(reset_i) begin
      opB_r_63_sv2v_reg <= 1'b0;
      opB_r_62_sv2v_reg <= 1'b0;
      opB_r_61_sv2v_reg <= 1'b0;
      opB_r_60_sv2v_reg <= 1'b0;
      opB_r_59_sv2v_reg <= 1'b0;
      opB_r_58_sv2v_reg <= 1'b0;
      opB_r_57_sv2v_reg <= 1'b0;
      opB_r_56_sv2v_reg <= 1'b0;
      opB_r_55_sv2v_reg <= 1'b0;
      opB_r_54_sv2v_reg <= 1'b0;
      opB_r_53_sv2v_reg <= 1'b0;
      opB_r_52_sv2v_reg <= 1'b0;
      opB_r_51_sv2v_reg <= 1'b0;
      opB_r_50_sv2v_reg <= 1'b0;
      opB_r_49_sv2v_reg <= 1'b0;
      opB_r_48_sv2v_reg <= 1'b0;
      opB_r_47_sv2v_reg <= 1'b0;
      opB_r_46_sv2v_reg <= 1'b0;
      opB_r_45_sv2v_reg <= 1'b0;
      opB_r_44_sv2v_reg <= 1'b0;
      opB_r_43_sv2v_reg <= 1'b0;
      opB_r_42_sv2v_reg <= 1'b0;
      opB_r_41_sv2v_reg <= 1'b0;
      opB_r_40_sv2v_reg <= 1'b0;
      opB_r_39_sv2v_reg <= 1'b0;
      opB_r_38_sv2v_reg <= 1'b0;
      opB_r_37_sv2v_reg <= 1'b0;
      opB_r_36_sv2v_reg <= 1'b0;
      opB_r_35_sv2v_reg <= 1'b0;
      opB_r_34_sv2v_reg <= 1'b0;
      opB_r_33_sv2v_reg <= 1'b0;
      opB_r_32_sv2v_reg <= 1'b0;
      opB_r_31_sv2v_reg <= 1'b0;
      opB_r_30_sv2v_reg <= 1'b0;
      opB_r_29_sv2v_reg <= 1'b0;
      opB_r_28_sv2v_reg <= 1'b0;
      opB_r_27_sv2v_reg <= 1'b0;
      opB_r_26_sv2v_reg <= 1'b0;
      opB_r_25_sv2v_reg <= 1'b0;
      opB_r_24_sv2v_reg <= 1'b0;
      opB_r_23_sv2v_reg <= 1'b0;
      opB_r_22_sv2v_reg <= 1'b0;
      opB_r_21_sv2v_reg <= 1'b0;
      opB_r_20_sv2v_reg <= 1'b0;
      opB_r_19_sv2v_reg <= 1'b0;
      opB_r_18_sv2v_reg <= 1'b0;
      opB_r_17_sv2v_reg <= 1'b0;
      opB_r_16_sv2v_reg <= 1'b0;
      opB_r_15_sv2v_reg <= 1'b0;
      opB_r_14_sv2v_reg <= 1'b0;
      opB_r_13_sv2v_reg <= 1'b0;
      opB_r_12_sv2v_reg <= 1'b0;
      opB_r_11_sv2v_reg <= 1'b0;
      opB_r_10_sv2v_reg <= 1'b0;
      opB_r_9_sv2v_reg <= 1'b0;
      opB_r_8_sv2v_reg <= 1'b0;
      opB_r_7_sv2v_reg <= 1'b0;
      opB_r_6_sv2v_reg <= 1'b0;
      opB_r_5_sv2v_reg <= 1'b0;
      opB_r_4_sv2v_reg <= 1'b0;
      opB_r_3_sv2v_reg <= 1'b0;
      opB_r_2_sv2v_reg <= 1'b0;
      opB_r_1_sv2v_reg <= 1'b0;
      opB_r_0_sv2v_reg <= 1'b0;
    end else if(N470) begin
      opB_r_63_sv2v_reg <= N534;
      opB_r_62_sv2v_reg <= N533;
      opB_r_61_sv2v_reg <= N532;
      opB_r_60_sv2v_reg <= N531;
      opB_r_59_sv2v_reg <= N530;
      opB_r_58_sv2v_reg <= N529;
      opB_r_57_sv2v_reg <= N528;
      opB_r_56_sv2v_reg <= N527;
      opB_r_55_sv2v_reg <= N526;
      opB_r_54_sv2v_reg <= N525;
      opB_r_53_sv2v_reg <= N524;
      opB_r_52_sv2v_reg <= N523;
      opB_r_51_sv2v_reg <= N522;
      opB_r_50_sv2v_reg <= N521;
      opB_r_49_sv2v_reg <= N520;
      opB_r_48_sv2v_reg <= N519;
      opB_r_47_sv2v_reg <= N518;
      opB_r_46_sv2v_reg <= N517;
      opB_r_45_sv2v_reg <= N516;
      opB_r_44_sv2v_reg <= N515;
      opB_r_43_sv2v_reg <= N514;
      opB_r_42_sv2v_reg <= N513;
      opB_r_41_sv2v_reg <= N512;
      opB_r_40_sv2v_reg <= N511;
      opB_r_39_sv2v_reg <= N510;
      opB_r_38_sv2v_reg <= N509;
      opB_r_37_sv2v_reg <= N508;
      opB_r_36_sv2v_reg <= N507;
      opB_r_35_sv2v_reg <= N506;
      opB_r_34_sv2v_reg <= N505;
      opB_r_33_sv2v_reg <= N504;
      opB_r_32_sv2v_reg <= N503;
      opB_r_31_sv2v_reg <= N502;
      opB_r_30_sv2v_reg <= N501;
      opB_r_29_sv2v_reg <= N500;
      opB_r_28_sv2v_reg <= N499;
      opB_r_27_sv2v_reg <= N498;
      opB_r_26_sv2v_reg <= N497;
      opB_r_25_sv2v_reg <= N496;
      opB_r_24_sv2v_reg <= N495;
      opB_r_23_sv2v_reg <= N494;
      opB_r_22_sv2v_reg <= N493;
      opB_r_21_sv2v_reg <= N492;
      opB_r_20_sv2v_reg <= N491;
      opB_r_19_sv2v_reg <= N490;
      opB_r_18_sv2v_reg <= N489;
      opB_r_17_sv2v_reg <= N488;
      opB_r_16_sv2v_reg <= N487;
      opB_r_15_sv2v_reg <= N486;
      opB_r_14_sv2v_reg <= N485;
      opB_r_13_sv2v_reg <= N484;
      opB_r_12_sv2v_reg <= N483;
      opB_r_11_sv2v_reg <= N482;
      opB_r_10_sv2v_reg <= N481;
      opB_r_9_sv2v_reg <= N480;
      opB_r_8_sv2v_reg <= N479;
      opB_r_7_sv2v_reg <= N478;
      opB_r_6_sv2v_reg <= N477;
      opB_r_5_sv2v_reg <= N476;
      opB_r_4_sv2v_reg <= N475;
      opB_r_3_sv2v_reg <= N474;
      opB_r_2_sv2v_reg <= N473;
      opB_r_1_sv2v_reg <= N472;
      opB_r_0_sv2v_reg <= N471;
    end 
    if(reset_i) begin
      all_sh_lsb_zero_r_sv2v_reg <= 1'b0;
    end else if(latch_input) begin
      all_sh_lsb_zero_r_sv2v_reg <= 1'b1;
    end else if(N810) begin
      all_sh_lsb_zero_r_sv2v_reg <= N536;
    end 
    if(N738) begin
      result_o_63_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_63_sv2v_reg <= N737;
    end 
    if(N801) begin
      result_o_62_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_62_sv2v_reg <= N736;
    end 
    if(N800) begin
      result_o_61_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_61_sv2v_reg <= N735;
    end 
    if(N799) begin
      result_o_60_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_60_sv2v_reg <= N734;
    end 
    if(N798) begin
      result_o_59_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_59_sv2v_reg <= N733;
    end 
    if(N797) begin
      result_o_58_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_58_sv2v_reg <= N732;
    end 
    if(N796) begin
      result_o_57_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_57_sv2v_reg <= N731;
    end 
    if(N795) begin
      result_o_56_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_56_sv2v_reg <= N730;
    end 
    if(N794) begin
      result_o_55_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_55_sv2v_reg <= N729;
    end 
    if(N793) begin
      result_o_54_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_54_sv2v_reg <= N728;
    end 
    if(N792) begin
      result_o_53_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_53_sv2v_reg <= N727;
    end 
    if(N791) begin
      result_o_52_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_52_sv2v_reg <= N726;
    end 
    if(N790) begin
      result_o_51_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_51_sv2v_reg <= N725;
    end 
    if(N789) begin
      result_o_50_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_50_sv2v_reg <= N724;
    end 
    if(N788) begin
      result_o_49_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_49_sv2v_reg <= N723;
    end 
    if(N787) begin
      result_o_48_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_48_sv2v_reg <= N722;
    end 
    if(N786) begin
      result_o_47_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_47_sv2v_reg <= N721;
    end 
    if(N785) begin
      result_o_46_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_46_sv2v_reg <= N720;
    end 
    if(N784) begin
      result_o_45_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_45_sv2v_reg <= N719;
    end 
    if(N783) begin
      result_o_44_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_44_sv2v_reg <= N718;
    end 
    if(N782) begin
      result_o_43_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_43_sv2v_reg <= N717;
    end 
    if(N781) begin
      result_o_42_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_42_sv2v_reg <= N716;
    end 
    if(N780) begin
      result_o_41_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_41_sv2v_reg <= N715;
    end 
    if(N779) begin
      result_o_40_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_40_sv2v_reg <= N714;
    end 
    if(N778) begin
      result_o_39_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_39_sv2v_reg <= N713;
    end 
    if(N777) begin
      result_o_38_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_38_sv2v_reg <= N712;
    end 
    if(N776) begin
      result_o_37_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_37_sv2v_reg <= N711;
    end 
    if(N775) begin
      result_o_36_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_36_sv2v_reg <= N710;
    end 
    if(N774) begin
      result_o_35_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_35_sv2v_reg <= N709;
    end 
    if(N773) begin
      result_o_34_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_34_sv2v_reg <= N708;
    end 
    if(N772) begin
      result_o_33_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_33_sv2v_reg <= N707;
    end 
    if(N771) begin
      result_o_32_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_32_sv2v_reg <= N706;
    end 
    if(N770) begin
      result_o_31_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_31_sv2v_reg <= N705;
    end 
    if(N769) begin
      result_o_30_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_30_sv2v_reg <= N704;
    end 
    if(N768) begin
      result_o_29_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_29_sv2v_reg <= N703;
    end 
    if(N767) begin
      result_o_28_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_28_sv2v_reg <= N702;
    end 
    if(N766) begin
      result_o_27_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_27_sv2v_reg <= N701;
    end 
    if(N765) begin
      result_o_26_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_26_sv2v_reg <= N700;
    end 
    if(N764) begin
      result_o_25_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_25_sv2v_reg <= N699;
    end 
    if(N763) begin
      result_o_24_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_24_sv2v_reg <= N698;
    end 
    if(N762) begin
      result_o_23_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_23_sv2v_reg <= N697;
    end 
    if(N761) begin
      result_o_22_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_22_sv2v_reg <= N696;
    end 
    if(N760) begin
      result_o_21_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_21_sv2v_reg <= N695;
    end 
    if(N759) begin
      result_o_20_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_20_sv2v_reg <= N694;
    end 
    if(N758) begin
      result_o_19_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_19_sv2v_reg <= N693;
    end 
    if(N757) begin
      result_o_18_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_18_sv2v_reg <= N692;
    end 
    if(N756) begin
      result_o_17_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_17_sv2v_reg <= N691;
    end 
    if(N755) begin
      result_o_16_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_16_sv2v_reg <= N690;
    end 
    if(N754) begin
      result_o_15_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_15_sv2v_reg <= N689;
    end 
    if(N753) begin
      result_o_14_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_14_sv2v_reg <= N688;
    end 
    if(N752) begin
      result_o_13_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_13_sv2v_reg <= N687;
    end 
    if(N751) begin
      result_o_12_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_12_sv2v_reg <= N686;
    end 
    if(N750) begin
      result_o_11_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_11_sv2v_reg <= N685;
    end 
    if(N749) begin
      result_o_10_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_10_sv2v_reg <= N684;
    end 
    if(N748) begin
      result_o_9_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_9_sv2v_reg <= N683;
    end 
    if(N747) begin
      result_o_8_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_8_sv2v_reg <= N682;
    end 
    if(N746) begin
      result_o_7_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_7_sv2v_reg <= N681;
    end 
    if(N745) begin
      result_o_6_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_6_sv2v_reg <= N680;
    end 
    if(N744) begin
      result_o_5_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_5_sv2v_reg <= N679;
    end 
    if(N743) begin
      result_o_4_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_4_sv2v_reg <= N678;
    end 
    if(N742) begin
      result_o_3_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_3_sv2v_reg <= N677;
    end 
    if(N741) begin
      result_o_2_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_2_sv2v_reg <= N676;
    end 
    if(N740) begin
      result_o_1_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_1_sv2v_reg <= N675;
    end 
    if(N739) begin
      result_o_0_sv2v_reg <= 1'b0;
    end else if(N673) begin
      result_o_0_sv2v_reg <= N674;
    end 
  end


endmodule



module bsg_dff_en_width_p1
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  input en_i;
  wire [0:0] data_o;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mux_one_hot_width_p65_els_p2
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [129:0] data_i;
  input [1:0] sel_one_hot_i;
  output [64:0] data_o;
  wire [64:0] data_o;
  wire [129:0] data_masked;
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[1];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[1];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[1];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[1];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[1];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_o[0] = data_masked[65] | data_masked[0];
  assign data_o[1] = data_masked[66] | data_masked[1];
  assign data_o[2] = data_masked[67] | data_masked[2];
  assign data_o[3] = data_masked[68] | data_masked[3];
  assign data_o[4] = data_masked[69] | data_masked[4];
  assign data_o[5] = data_masked[70] | data_masked[5];
  assign data_o[6] = data_masked[71] | data_masked[6];
  assign data_o[7] = data_masked[72] | data_masked[7];
  assign data_o[8] = data_masked[73] | data_masked[8];
  assign data_o[9] = data_masked[74] | data_masked[9];
  assign data_o[10] = data_masked[75] | data_masked[10];
  assign data_o[11] = data_masked[76] | data_masked[11];
  assign data_o[12] = data_masked[77] | data_masked[12];
  assign data_o[13] = data_masked[78] | data_masked[13];
  assign data_o[14] = data_masked[79] | data_masked[14];
  assign data_o[15] = data_masked[80] | data_masked[15];
  assign data_o[16] = data_masked[81] | data_masked[16];
  assign data_o[17] = data_masked[82] | data_masked[17];
  assign data_o[18] = data_masked[83] | data_masked[18];
  assign data_o[19] = data_masked[84] | data_masked[19];
  assign data_o[20] = data_masked[85] | data_masked[20];
  assign data_o[21] = data_masked[86] | data_masked[21];
  assign data_o[22] = data_masked[87] | data_masked[22];
  assign data_o[23] = data_masked[88] | data_masked[23];
  assign data_o[24] = data_masked[89] | data_masked[24];
  assign data_o[25] = data_masked[90] | data_masked[25];
  assign data_o[26] = data_masked[91] | data_masked[26];
  assign data_o[27] = data_masked[92] | data_masked[27];
  assign data_o[28] = data_masked[93] | data_masked[28];
  assign data_o[29] = data_masked[94] | data_masked[29];
  assign data_o[30] = data_masked[95] | data_masked[30];
  assign data_o[31] = data_masked[96] | data_masked[31];
  assign data_o[32] = data_masked[97] | data_masked[32];
  assign data_o[33] = data_masked[98] | data_masked[33];
  assign data_o[34] = data_masked[99] | data_masked[34];
  assign data_o[35] = data_masked[100] | data_masked[35];
  assign data_o[36] = data_masked[101] | data_masked[36];
  assign data_o[37] = data_masked[102] | data_masked[37];
  assign data_o[38] = data_masked[103] | data_masked[38];
  assign data_o[39] = data_masked[104] | data_masked[39];
  assign data_o[40] = data_masked[105] | data_masked[40];
  assign data_o[41] = data_masked[106] | data_masked[41];
  assign data_o[42] = data_masked[107] | data_masked[42];
  assign data_o[43] = data_masked[108] | data_masked[43];
  assign data_o[44] = data_masked[109] | data_masked[44];
  assign data_o[45] = data_masked[110] | data_masked[45];
  assign data_o[46] = data_masked[111] | data_masked[46];
  assign data_o[47] = data_masked[112] | data_masked[47];
  assign data_o[48] = data_masked[113] | data_masked[48];
  assign data_o[49] = data_masked[114] | data_masked[49];
  assign data_o[50] = data_masked[115] | data_masked[50];
  assign data_o[51] = data_masked[116] | data_masked[51];
  assign data_o[52] = data_masked[117] | data_masked[52];
  assign data_o[53] = data_masked[118] | data_masked[53];
  assign data_o[54] = data_masked[119] | data_masked[54];
  assign data_o[55] = data_masked[120] | data_masked[55];
  assign data_o[56] = data_masked[121] | data_masked[56];
  assign data_o[57] = data_masked[122] | data_masked[57];
  assign data_o[58] = data_masked[123] | data_masked[58];
  assign data_o[59] = data_masked[124] | data_masked[59];
  assign data_o[60] = data_masked[125] | data_masked[60];
  assign data_o[61] = data_masked[126] | data_masked[61];
  assign data_o[62] = data_masked[127] | data_masked[62];
  assign data_o[63] = data_masked[128] | data_masked[63];
  assign data_o[64] = data_masked[129] | data_masked[64];

endmodule



module bsg_mux_one_hot_width_p65_els_p4
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [259:0] data_i;
  input [3:0] sel_one_hot_i;
  output [64:0] data_o;
  wire [64:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129;
  wire [259:0] data_masked;
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[1];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[1];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[1];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[1];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[1];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[2];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[2];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[2];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[2];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[2];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[2];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[2];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[2];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[2];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[2];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[2];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[2];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[2];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[2];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[2];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[2];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[2];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[2];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[2];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[2];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[2];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[2];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[2];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[2];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[2];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[2];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[2];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[2];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[2];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[2];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[2];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[2];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[2];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[2];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[2];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[2];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[2];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[2];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[2];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[2];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[2];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[2];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[2];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[2];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[2];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[2];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[2];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[2];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[2];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[2];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[2];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[2];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[2];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[2];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[2];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[2];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[2];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[2];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[2];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[2];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[2];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[2];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[2];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[2];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[2];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[3];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[3];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[3];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[3];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[3];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[3];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[3];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[3];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[3];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[3];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[3];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[3];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[3];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[3];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[3];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[3];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[3];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[3];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[3];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[3];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[3];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[3];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[3];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[3];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[3];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[3];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[3];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[3];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[3];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[3];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[3];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[3];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[3];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[3];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[3];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[3];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[3];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[3];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[3];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[3];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[3];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[3];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[3];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[3];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[3];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[3];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[3];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[3];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[3];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[3];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[3];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[3];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[3];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[3];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[3];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[3];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[3];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[3];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[3];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[3];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[3];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[3];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[3];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[3];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[3];
  assign data_o[0] = N1 | data_masked[0];
  assign N1 = N0 | data_masked[65];
  assign N0 = data_masked[195] | data_masked[130];
  assign data_o[1] = N3 | data_masked[1];
  assign N3 = N2 | data_masked[66];
  assign N2 = data_masked[196] | data_masked[131];
  assign data_o[2] = N5 | data_masked[2];
  assign N5 = N4 | data_masked[67];
  assign N4 = data_masked[197] | data_masked[132];
  assign data_o[3] = N7 | data_masked[3];
  assign N7 = N6 | data_masked[68];
  assign N6 = data_masked[198] | data_masked[133];
  assign data_o[4] = N9 | data_masked[4];
  assign N9 = N8 | data_masked[69];
  assign N8 = data_masked[199] | data_masked[134];
  assign data_o[5] = N11 | data_masked[5];
  assign N11 = N10 | data_masked[70];
  assign N10 = data_masked[200] | data_masked[135];
  assign data_o[6] = N13 | data_masked[6];
  assign N13 = N12 | data_masked[71];
  assign N12 = data_masked[201] | data_masked[136];
  assign data_o[7] = N15 | data_masked[7];
  assign N15 = N14 | data_masked[72];
  assign N14 = data_masked[202] | data_masked[137];
  assign data_o[8] = N17 | data_masked[8];
  assign N17 = N16 | data_masked[73];
  assign N16 = data_masked[203] | data_masked[138];
  assign data_o[9] = N19 | data_masked[9];
  assign N19 = N18 | data_masked[74];
  assign N18 = data_masked[204] | data_masked[139];
  assign data_o[10] = N21 | data_masked[10];
  assign N21 = N20 | data_masked[75];
  assign N20 = data_masked[205] | data_masked[140];
  assign data_o[11] = N23 | data_masked[11];
  assign N23 = N22 | data_masked[76];
  assign N22 = data_masked[206] | data_masked[141];
  assign data_o[12] = N25 | data_masked[12];
  assign N25 = N24 | data_masked[77];
  assign N24 = data_masked[207] | data_masked[142];
  assign data_o[13] = N27 | data_masked[13];
  assign N27 = N26 | data_masked[78];
  assign N26 = data_masked[208] | data_masked[143];
  assign data_o[14] = N29 | data_masked[14];
  assign N29 = N28 | data_masked[79];
  assign N28 = data_masked[209] | data_masked[144];
  assign data_o[15] = N31 | data_masked[15];
  assign N31 = N30 | data_masked[80];
  assign N30 = data_masked[210] | data_masked[145];
  assign data_o[16] = N33 | data_masked[16];
  assign N33 = N32 | data_masked[81];
  assign N32 = data_masked[211] | data_masked[146];
  assign data_o[17] = N35 | data_masked[17];
  assign N35 = N34 | data_masked[82];
  assign N34 = data_masked[212] | data_masked[147];
  assign data_o[18] = N37 | data_masked[18];
  assign N37 = N36 | data_masked[83];
  assign N36 = data_masked[213] | data_masked[148];
  assign data_o[19] = N39 | data_masked[19];
  assign N39 = N38 | data_masked[84];
  assign N38 = data_masked[214] | data_masked[149];
  assign data_o[20] = N41 | data_masked[20];
  assign N41 = N40 | data_masked[85];
  assign N40 = data_masked[215] | data_masked[150];
  assign data_o[21] = N43 | data_masked[21];
  assign N43 = N42 | data_masked[86];
  assign N42 = data_masked[216] | data_masked[151];
  assign data_o[22] = N45 | data_masked[22];
  assign N45 = N44 | data_masked[87];
  assign N44 = data_masked[217] | data_masked[152];
  assign data_o[23] = N47 | data_masked[23];
  assign N47 = N46 | data_masked[88];
  assign N46 = data_masked[218] | data_masked[153];
  assign data_o[24] = N49 | data_masked[24];
  assign N49 = N48 | data_masked[89];
  assign N48 = data_masked[219] | data_masked[154];
  assign data_o[25] = N51 | data_masked[25];
  assign N51 = N50 | data_masked[90];
  assign N50 = data_masked[220] | data_masked[155];
  assign data_o[26] = N53 | data_masked[26];
  assign N53 = N52 | data_masked[91];
  assign N52 = data_masked[221] | data_masked[156];
  assign data_o[27] = N55 | data_masked[27];
  assign N55 = N54 | data_masked[92];
  assign N54 = data_masked[222] | data_masked[157];
  assign data_o[28] = N57 | data_masked[28];
  assign N57 = N56 | data_masked[93];
  assign N56 = data_masked[223] | data_masked[158];
  assign data_o[29] = N59 | data_masked[29];
  assign N59 = N58 | data_masked[94];
  assign N58 = data_masked[224] | data_masked[159];
  assign data_o[30] = N61 | data_masked[30];
  assign N61 = N60 | data_masked[95];
  assign N60 = data_masked[225] | data_masked[160];
  assign data_o[31] = N63 | data_masked[31];
  assign N63 = N62 | data_masked[96];
  assign N62 = data_masked[226] | data_masked[161];
  assign data_o[32] = N65 | data_masked[32];
  assign N65 = N64 | data_masked[97];
  assign N64 = data_masked[227] | data_masked[162];
  assign data_o[33] = N67 | data_masked[33];
  assign N67 = N66 | data_masked[98];
  assign N66 = data_masked[228] | data_masked[163];
  assign data_o[34] = N69 | data_masked[34];
  assign N69 = N68 | data_masked[99];
  assign N68 = data_masked[229] | data_masked[164];
  assign data_o[35] = N71 | data_masked[35];
  assign N71 = N70 | data_masked[100];
  assign N70 = data_masked[230] | data_masked[165];
  assign data_o[36] = N73 | data_masked[36];
  assign N73 = N72 | data_masked[101];
  assign N72 = data_masked[231] | data_masked[166];
  assign data_o[37] = N75 | data_masked[37];
  assign N75 = N74 | data_masked[102];
  assign N74 = data_masked[232] | data_masked[167];
  assign data_o[38] = N77 | data_masked[38];
  assign N77 = N76 | data_masked[103];
  assign N76 = data_masked[233] | data_masked[168];
  assign data_o[39] = N79 | data_masked[39];
  assign N79 = N78 | data_masked[104];
  assign N78 = data_masked[234] | data_masked[169];
  assign data_o[40] = N81 | data_masked[40];
  assign N81 = N80 | data_masked[105];
  assign N80 = data_masked[235] | data_masked[170];
  assign data_o[41] = N83 | data_masked[41];
  assign N83 = N82 | data_masked[106];
  assign N82 = data_masked[236] | data_masked[171];
  assign data_o[42] = N85 | data_masked[42];
  assign N85 = N84 | data_masked[107];
  assign N84 = data_masked[237] | data_masked[172];
  assign data_o[43] = N87 | data_masked[43];
  assign N87 = N86 | data_masked[108];
  assign N86 = data_masked[238] | data_masked[173];
  assign data_o[44] = N89 | data_masked[44];
  assign N89 = N88 | data_masked[109];
  assign N88 = data_masked[239] | data_masked[174];
  assign data_o[45] = N91 | data_masked[45];
  assign N91 = N90 | data_masked[110];
  assign N90 = data_masked[240] | data_masked[175];
  assign data_o[46] = N93 | data_masked[46];
  assign N93 = N92 | data_masked[111];
  assign N92 = data_masked[241] | data_masked[176];
  assign data_o[47] = N95 | data_masked[47];
  assign N95 = N94 | data_masked[112];
  assign N94 = data_masked[242] | data_masked[177];
  assign data_o[48] = N97 | data_masked[48];
  assign N97 = N96 | data_masked[113];
  assign N96 = data_masked[243] | data_masked[178];
  assign data_o[49] = N99 | data_masked[49];
  assign N99 = N98 | data_masked[114];
  assign N98 = data_masked[244] | data_masked[179];
  assign data_o[50] = N101 | data_masked[50];
  assign N101 = N100 | data_masked[115];
  assign N100 = data_masked[245] | data_masked[180];
  assign data_o[51] = N103 | data_masked[51];
  assign N103 = N102 | data_masked[116];
  assign N102 = data_masked[246] | data_masked[181];
  assign data_o[52] = N105 | data_masked[52];
  assign N105 = N104 | data_masked[117];
  assign N104 = data_masked[247] | data_masked[182];
  assign data_o[53] = N107 | data_masked[53];
  assign N107 = N106 | data_masked[118];
  assign N106 = data_masked[248] | data_masked[183];
  assign data_o[54] = N109 | data_masked[54];
  assign N109 = N108 | data_masked[119];
  assign N108 = data_masked[249] | data_masked[184];
  assign data_o[55] = N111 | data_masked[55];
  assign N111 = N110 | data_masked[120];
  assign N110 = data_masked[250] | data_masked[185];
  assign data_o[56] = N113 | data_masked[56];
  assign N113 = N112 | data_masked[121];
  assign N112 = data_masked[251] | data_masked[186];
  assign data_o[57] = N115 | data_masked[57];
  assign N115 = N114 | data_masked[122];
  assign N114 = data_masked[252] | data_masked[187];
  assign data_o[58] = N117 | data_masked[58];
  assign N117 = N116 | data_masked[123];
  assign N116 = data_masked[253] | data_masked[188];
  assign data_o[59] = N119 | data_masked[59];
  assign N119 = N118 | data_masked[124];
  assign N118 = data_masked[254] | data_masked[189];
  assign data_o[60] = N121 | data_masked[60];
  assign N121 = N120 | data_masked[125];
  assign N120 = data_masked[255] | data_masked[190];
  assign data_o[61] = N123 | data_masked[61];
  assign N123 = N122 | data_masked[126];
  assign N122 = data_masked[256] | data_masked[191];
  assign data_o[62] = N125 | data_masked[62];
  assign N125 = N124 | data_masked[127];
  assign N124 = data_masked[257] | data_masked[192];
  assign data_o[63] = N127 | data_masked[63];
  assign N127 = N126 | data_masked[128];
  assign N126 = data_masked[258] | data_masked[193];
  assign data_o[64] = N129 | data_masked[64];
  assign N129 = N128 | data_masked[129];
  assign N128 = data_masked[259] | data_masked[194];

endmodule



module bsg_dff_en_width_p65
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [64:0] data_i;
  output [64:0] data_o;
  input clk_i;
  input en_i;
  wire [64:0] data_o;
  reg data_o_64_sv2v_reg,data_o_63_sv2v_reg,data_o_62_sv2v_reg,data_o_61_sv2v_reg,
  data_o_60_sv2v_reg,data_o_59_sv2v_reg,data_o_58_sv2v_reg,data_o_57_sv2v_reg,
  data_o_56_sv2v_reg,data_o_55_sv2v_reg,data_o_54_sv2v_reg,data_o_53_sv2v_reg,
  data_o_52_sv2v_reg,data_o_51_sv2v_reg,data_o_50_sv2v_reg,data_o_49_sv2v_reg,
  data_o_48_sv2v_reg,data_o_47_sv2v_reg,data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,
  data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,
  data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,
  data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,
  data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,
  data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,
  data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,
  data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,
  data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_adder_cin_width_p65
(
  a_i,
  b_i,
  cin_i,
  o
);

  input [64:0] a_i;
  input [64:0] b_i;
  output [64:0] o;
  input cin_i;
  wire [64:0] o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64;
  assign { N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0 } = a_i + b_i;
  assign o = { N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0 } + cin_i;

endmodule



module bsg_counter_clear_up_00000020_0_1
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [5:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire [5:0] count_o;
  wire N0,N1,N4,N5,N6,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N2,N3,N7,N30,N19;
  reg count_o_5_sv2v_reg,count_o_4_sv2v_reg,count_o_3_sv2v_reg,count_o_2_sv2v_reg,
  count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[5] = count_o_5_sv2v_reg;
  assign count_o[4] = count_o_4_sv2v_reg;
  assign count_o[3] = count_o_3_sv2v_reg;
  assign count_o[2] = count_o_2_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign N19 = reset_i | clear_i;
  assign { N11, N10, N9, N8, N6, N5 } = count_o + 1'b1;
  assign N12 = (N0)? 1'b1 : 
               (N7)? 1'b1 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = clear_i;
  assign N14 = (N1)? 1'b1 : 
               (N30)? 1'b0 : 1'b0;
  assign N1 = up_i;
  assign N13 = (N0)? up_i : 
               (N7)? N5 : 1'b0;
  assign N4 = N18;
  assign N15 = ~reset_i;
  assign N16 = ~clear_i;
  assign N17 = N15 & N16;
  assign N18 = up_i & N17;
  assign N2 = up_i | clear_i;
  assign N3 = ~N2;
  assign N7 = up_i & N16;
  assign N30 = ~up_i;

  always @(posedge clk_i) begin
    if(N19) begin
      count_o_5_sv2v_reg <= 1'b0;
      count_o_4_sv2v_reg <= 1'b0;
      count_o_3_sv2v_reg <= 1'b0;
      count_o_2_sv2v_reg <= 1'b0;
      count_o_1_sv2v_reg <= 1'b0;
    end else if(N14) begin
      count_o_5_sv2v_reg <= N11;
      count_o_4_sv2v_reg <= N10;
      count_o_3_sv2v_reg <= N9;
      count_o_2_sv2v_reg <= N8;
      count_o_1_sv2v_reg <= N6;
    end 
    if(reset_i) begin
      count_o_0_sv2v_reg <= 1'b0;
    end else if(N12) begin
      count_o_0_sv2v_reg <= N13;
    end 
  end


endmodule



module bsg_idiv_iterative_controller_64_2
(
  clk_i,
  reset_i,
  v_i,
  ready_and_o,
  zero_divisor_i,
  signed_div_r_i,
  adder1_result_is_neg_i,
  adder2_result_is_neg_i,
  opA_is_neg_i,
  opC_is_neg_i,
  opA_sel_o,
  opA_ld_o,
  opA_inv_o,
  opA_clr_l_o,
  opB_sel_o,
  opB_ld_o,
  opB_inv_o,
  opB_clr_l_o,
  opC_sel_o,
  opC_ld_o,
  latch_signed_div_o,
  adder1_cin_o,
  v_o,
  yumi_i
);

  output [1:0] opA_sel_o;
  output [3:0] opB_sel_o;
  output [3:0] opC_sel_o;
  input clk_i;
  input reset_i;
  input v_i;
  input zero_divisor_i;
  input signed_div_r_i;
  input adder1_result_is_neg_i;
  input adder2_result_is_neg_i;
  input opA_is_neg_i;
  input opC_is_neg_i;
  input yumi_i;
  output ready_and_o;
  output opA_ld_o;
  output opA_inv_o;
  output opA_clr_l_o;
  output opB_ld_o;
  output opB_inv_o;
  output opB_clr_l_o;
  output opC_ld_o;
  output latch_signed_div_o;
  output adder1_cin_o;
  output v_o;
  wire [1:0] opA_sel_o;
  wire [3:0] opB_sel_o,opC_sel_o,next_state;
  wire ready_and_o,opA_ld_o,opA_inv_o,opA_clr_l_o,opB_ld_o,opB_inv_o,opB_clr_l_o,
  opC_ld_o,latch_signed_div_o,adder1_cin_o,v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,
  N12,N13,add1_neg_last_r,add2_neg_last_r,neg_ld,N14,q_neg_r,N15,r_neg_r,calc_up_li,
  N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,
  N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,
  N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,
  N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,
  N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N110,N111,N112,N113,
  N114,N115,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138;
  wire [5:0] state,calc_cnt;
  reg add1_neg_last_r_sv2v_reg,add2_neg_last_r_sv2v_reg,r_neg_r_sv2v_reg,
  q_neg_r_sv2v_reg,state_5_sv2v_reg,state_4_sv2v_reg,state_3_sv2v_reg,state_2_sv2v_reg,
  state_1_sv2v_reg,state_0_sv2v_reg;
  assign add1_neg_last_r = add1_neg_last_r_sv2v_reg;
  assign add2_neg_last_r = add2_neg_last_r_sv2v_reg;
  assign r_neg_r = r_neg_r_sv2v_reg;
  assign q_neg_r = q_neg_r_sv2v_reg;
  assign state[5] = state_5_sv2v_reg;
  assign state[4] = state_4_sv2v_reg;
  assign state[3] = state_3_sv2v_reg;
  assign state[2] = state_2_sv2v_reg;
  assign state[1] = state_1_sv2v_reg;
  assign state[0] = state_0_sv2v_reg;

  bsg_counter_clear_up_00000020_0_1
  calc_counter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(N136),
    .up_i(calc_up_li),
    .count_o(calc_cnt)
  );

  assign N19 = N17 & N18;
  assign N22 = N110 & N117;
  assign N23 = N20 & N21;
  assign N24 = N22 & N23;
  assign N25 = state[3] | state[2];
  assign N26 = state[1] | N21;
  assign N27 = N25 | N26;
  assign N29 = state[3] | state[2];
  assign N30 = N20 | state[0];
  assign N31 = N29 | N30;
  assign N33 = state[3] | state[2];
  assign N34 = N20 | N21;
  assign N35 = N33 | N34;
  assign N37 = state[3] | N117;
  assign N38 = state[1] | state[0];
  assign N39 = N37 | N38;
  assign N41 = state[3] | N117;
  assign N42 = state[1] | N21;
  assign N43 = N41 | N42;
  assign N45 = state[3] | N117;
  assign N46 = N20 | state[0];
  assign N47 = N45 | N46;
  assign N49 = state[3] | N117;
  assign N50 = N20 | N21;
  assign N51 = N49 | N50;
  assign N53 = N110 | state[2];
  assign N54 = state[1] | state[0];
  assign N55 = N53 | N54;
  assign N104 = state[4] | state[5];
  assign N105 = state[3] | N104;
  assign N106 = state[2] | N105;
  assign N107 = state[1] | N106;
  assign N108 = state[0] | N107;
  assign ready_and_o = ~N108;
  assign N110 = ~state[3];
  assign N111 = state[4] | state[5];
  assign N112 = N110 | N111;
  assign N113 = state[2] | N112;
  assign N114 = state[1] | N113;
  assign N115 = state[0] | N114;
  assign v_o = ~N115;
  assign N117 = ~state[2];
  assign N118 = state[4] | state[5];
  assign N119 = state[3] | N118;
  assign N120 = N117 | N119;
  assign N121 = state[1] | N120;
  assign N122 = state[0] | N121;
  assign N123 = ~N122;
  assign N124 = calc_cnt[4] | calc_cnt[5];
  assign N125 = calc_cnt[3] | N124;
  assign N126 = calc_cnt[2] | N125;
  assign N127 = calc_cnt[1] | N126;
  assign N128 = calc_cnt[0] | N127;
  assign N129 = ~N128;
  assign N130 = ~calc_cnt[5];
  assign N131 = calc_cnt[4] | N130;
  assign N132 = calc_cnt[3] | N131;
  assign N133 = calc_cnt[2] | N132;
  assign N134 = calc_cnt[1] | N133;
  assign N135 = calc_cnt[0] | N134;
  assign N136 = ~N135;
  assign N58 = ~N15;
  assign N63 = (N0)? N62 : 
               (N1)? N16 : 1'b0;
  assign N0 = N129;
  assign N1 = N128;
  assign N64 = (N0)? N62 : 
               (N1)? N16 : 1'b0;
  assign { N67, N66 } = (N2)? { N65, adder1_result_is_neg_i } : 
                        (N3)? { 1'b0, 1'b0 } : 1'b0;
  assign N2 = N61;
  assign N3 = N60;
  assign N69 = ~N68;
  assign { N82, N81, N80 } = (N4)? { 1'b0, 1'b0, N57 } : 
                             (N5)? { 1'b0, 1'b0, 1'b1 } : 
                             (N6)? { 1'b1, 1'b0, 1'b0 } : 
                             (N7)? { 1'b0, 1'b1, 1'b0 } : 
                             (N8)? { 1'b0, N61, N60 } : 
                             (N9)? { 1'b0, 1'b0, 1'b1 } : 
                             (N10)? { 1'b0, 1'b0, 1'b1 } : 
                             (N11)? { 1'b1, 1'b0, 1'b0 } : 
                             (N12)? { 1'b0, 1'b0, 1'b1 } : 
                             (N79)? { 1'b0, 1'b0, 1'b1 } : 1'b0;
  assign N4 = N24;
  assign N5 = N28;
  assign N6 = N32;
  assign N7 = N36;
  assign N8 = N40;
  assign N9 = N44;
  assign N10 = N48;
  assign N11 = N52;
  assign N12 = N56;
  assign N85 = (N4)? v_i : 
               (N84)? 1'b0 : 1'b0;
  assign N86 = (N4)? v_i : 
               (N5)? N59 : 
               (N6)? 1'b0 : 
               (N7)? 1'b0 : 
               (N8)? 1'b0 : 
               (N9)? 1'b0 : 
               (N10)? 1'b1 : 
               (N11)? 1'b0 : 
               (N12)? 1'b0 : 
               (N79)? 1'b0 : 1'b0;
  assign N87 = (N4)? v_i : 
               (N5)? 1'b0 : 
               (N6)? 1'b1 : 
               (N7)? 1'b1 : 
               (N8)? 1'b1 : 
               (N9)? 1'b0 : 
               (N10)? 1'b0 : 
               (N11)? 1'b1 : 
               (N12)? 1'b0 : 
               (N79)? 1'b0 : 1'b0;
  assign N88 = (N4)? v_i : 
               (N5)? 1'b0 : 
               (N6)? 1'b0 : 
               (N7)? 1'b0 : 
               (N8)? 1'b0 : 
               (N9)? 1'b0 : 
               (N10)? 1'b0 : 
               (N11)? 1'b0 : 
               (N12)? 1'b0 : 
               (N79)? 1'b0 : 1'b0;
  assign { N92, N91, N90, N89 } = (N4)? { 1'b0, 1'b0, 1'b0, v_i } : 
                                  (N5)? { 1'b0, 1'b0, 1'b1, N58 } : 
                                  (N6)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                  (N7)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                  (N8)? { 1'b0, 1'b1, N67, N66 } : 
                                  (N9)? { 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                  (N10)? { N68, N69, N69, N69 } : 
                                  (N11)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                  (N12)? { N70, 1'b0, 1'b0, 1'b0 } : 
                                  (N79)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N93 = (N4)? 1'b0 : 
               (N5)? 1'b1 : 
               (N6)? 1'b0 : 
               (N7)? 1'b0 : 
               (N8)? 1'b0 : 
               (N9)? 1'b0 : 
               (N10)? 1'b1 : 
               (N11)? 1'b0 : 
               (N12)? 1'b0 : 
               (N79)? 1'b0 : 1'b0;
  assign N94 = (N4)? N16 : 
               (N5)? 1'b1 : 
               (N6)? N16 : 
               (N7)? N16 : 
               (N8)? N63 : 
               (N9)? 1'b0 : 
               (N10)? N16 : 
               (N11)? N16 : 
               (N12)? N16 : 
               (N79)? N16 : 1'b0;
  assign N95 = (N4)? 1'b1 : 
               (N5)? 1'b0 : 
               (N6)? 1'b1 : 
               (N7)? 1'b0 : 
               (N8)? 1'b1 : 
               (N9)? 1'b1 : 
               (N10)? 1'b1 : 
               (N11)? 1'b1 : 
               (N12)? 1'b1 : 
               (N79)? 1'b1 : 1'b0;
  assign N96 = (N4)? 1'b0 : 
               (N5)? 1'b1 : 
               (N6)? 1'b0 : 
               (N7)? 1'b1 : 
               (N8)? 1'b1 : 
               (N9)? 1'b1 : 
               (N10)? 1'b1 : 
               (N11)? 1'b0 : 
               (N12)? 1'b0 : 
               (N79)? 1'b0 : 1'b0;
  assign N97 = (N4)? 1'b0 : 
               (N5)? 1'b1 : 
               (N6)? 1'b0 : 
               (N7)? 1'b0 : 
               (N8)? 1'b0 : 
               (N9)? 1'b0 : 
               (N10)? 1'b0 : 
               (N11)? 1'b0 : 
               (N12)? 1'b0 : 
               (N79)? 1'b0 : 1'b0;
  assign N98 = (N4)? N16 : 
               (N5)? 1'b1 : 
               (N6)? 1'b1 : 
               (N7)? 1'b0 : 
               (N8)? N64 : 
               (N9)? 1'b0 : 
               (N10)? r_neg_r : 
               (N11)? 1'b1 : 
               (N12)? N16 : 
               (N79)? N16 : 1'b0;
  assign { N100, N99 } = (N4)? { 1'b0, 1'b1 } : 
                         (N5)? { 1'b0, 1'b0 } : 
                         (N6)? { 1'b0, 1'b1 } : 
                         (N7)? { 1'b0, 1'b0 } : 
                         (N8)? { N61, N60 } : 
                         (N9)? { 1'b1, 1'b0 } : 
                         (N10)? { 1'b0, 1'b0 } : 
                         (N11)? { 1'b0, 1'b1 } : 
                         (N12)? { 1'b0, 1'b1 } : 
                         (N79)? { 1'b0, 1'b1 } : 1'b0;
  assign N101 = (N4)? 1'b1 : 
                (N5)? 1'b1 : 
                (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N8)? 1'b1 : 
                (N9)? 1'b1 : 
                (N10)? 1'b0 : 
                (N11)? 1'b0 : 
                (N12)? 1'b1 : 
                (N79)? 1'b1 : 1'b0;
  assign N102 = (N4)? 1'b0 : 
                (N5)? 1'b0 : 
                (N6)? 1'b1 : 
                (N7)? 1'b0 : 
                (N8)? 1'b0 : 
                (N9)? 1'b0 : 
                (N10)? r_neg_r : 
                (N11)? 1'b1 : 
                (N12)? 1'b0 : 
                (N79)? 1'b0 : 1'b0;
  assign opA_clr_l_o = (N13)? N101 : 
                       (N103)? 1'b1 : 1'b0;
  assign N13 = N19;
  assign opB_inv_o = (N13)? N102 : 
                     (N103)? 1'b0 : 1'b0;
  assign opC_sel_o = (N13)? { N85, N82, N81, N80 } : 
                     (N103)? { 1'b0, 1'b0, 1'b0, 1'b1 } : 1'b0;
  assign opA_ld_o = (N13)? N86 : 
                    (N103)? 1'b0 : 1'b0;
  assign opC_ld_o = (N13)? N87 : 
                    (N103)? 1'b0 : 1'b0;
  assign latch_signed_div_o = (N13)? N88 : 
                              (N103)? 1'b0 : 1'b0;
  assign next_state = (N13)? { N92, N91, N90, N89 } : 
                      (N103)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign opA_sel_o = (N13)? { N85, N93 } : 
                     (N103)? { 1'b0, 1'b0 } : 1'b0;
  assign opA_inv_o = (N13)? N94 : 
                     (N103)? N16 : 1'b0;
  assign opB_clr_l_o = (N13)? N95 : 
                       (N103)? 1'b1 : 1'b0;
  assign opB_ld_o = (N13)? N96 : 
                    (N103)? 1'b0 : 1'b0;
  assign neg_ld = (N13)? N97 : 
                  (N103)? 1'b0 : 1'b0;
  assign adder1_cin_o = (N13)? N98 : 
                        (N103)? N16 : 1'b0;
  assign opB_sel_o = (N13)? { N93, N100, N36, N99 } : 
                     (N103)? { 1'b0, 1'b0, 1'b0, 1'b1 } : 1'b0;
  assign N14 = N137 & signed_div_r_i;
  assign N137 = opA_is_neg_i ^ opC_is_neg_i;
  assign N15 = opC_is_neg_i & signed_div_r_i;
  assign calc_up_li = N123 & N130;
  assign N16 = ~add2_neg_last_r;
  assign N17 = ~state[5];
  assign N18 = ~state[4];
  assign N20 = ~state[1];
  assign N21 = ~state[0];
  assign N28 = ~N27;
  assign N32 = ~N31;
  assign N36 = ~N35;
  assign N40 = ~N39;
  assign N44 = ~N43;
  assign N48 = ~N47;
  assign N52 = ~N51;
  assign N56 = ~N55;
  assign N57 = ~v_i;
  assign N59 = opA_is_neg_i & signed_div_r_i;
  assign N60 = ~N136;
  assign N61 = N136;
  assign N62 = ~add1_neg_last_r;
  assign N65 = ~adder1_result_is_neg_i;
  assign N68 = zero_divisor_i | N138;
  assign N138 = ~q_neg_r;
  assign N70 = ~yumi_i;
  assign N71 = N28 | N24;
  assign N72 = N32 | N71;
  assign N73 = N36 | N72;
  assign N74 = N40 | N73;
  assign N75 = N44 | N74;
  assign N76 = N48 | N75;
  assign N77 = N52 | N76;
  assign N78 = N56 | N77;
  assign N79 = ~N78;
  assign N83 = ~N24;
  assign N84 = N83;
  assign N103 = ~N19;

  always @(posedge clk_i) begin
    if(1'b1) begin
      add1_neg_last_r_sv2v_reg <= adder1_result_is_neg_i;
      add2_neg_last_r_sv2v_reg <= adder2_result_is_neg_i;
    end 
    if(neg_ld) begin
      r_neg_r_sv2v_reg <= N15;
      q_neg_r_sv2v_reg <= N14;
    end 
    if(reset_i) begin
      state_5_sv2v_reg <= 1'b0;
      state_4_sv2v_reg <= 1'b0;
      state_3_sv2v_reg <= 1'b0;
      state_2_sv2v_reg <= 1'b0;
      state_1_sv2v_reg <= 1'b0;
      state_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      state_5_sv2v_reg <= 1'b0;
      state_4_sv2v_reg <= 1'b0;
      state_3_sv2v_reg <= next_state[3];
      state_2_sv2v_reg <= next_state[2];
      state_1_sv2v_reg <= next_state[1];
      state_0_sv2v_reg <= next_state[0];
    end 
  end


endmodule



module bsg_idiv_iterative_64_2
(
  clk_i,
  reset_i,
  v_i,
  ready_and_o,
  dividend_i,
  divisor_i,
  signed_div_i,
  v_o,
  quotient_o,
  remainder_o,
  yumi_i
);

  input [63:0] dividend_i;
  input [63:0] divisor_i;
  output [63:0] quotient_o;
  output [63:0] remainder_o;
  input clk_i;
  input reset_i;
  input v_i;
  input signed_div_i;
  input yumi_i;
  output ready_and_o;
  output v_o;
  wire [63:0] quotient_o,remainder_o;
  wire ready_and_o,v_o,divisor_msb,dividend_msb,signed_div_r,latch_signed_div_lo,
  zero_divisor_li,_2_net__65_,_2_net__1_,_2_net__0_,opA_ld_lo,opB_ld_lo,opC_ld_lo,
  opA_inv_lo,opA_clr_lo,opB_inv_lo,opB_clr_lo,adder1_cin_lo,\genblk3.adder2_cin ,N0,N1,
  N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,
  N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,
  N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,
  N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,
  N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,
  N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,
  N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,
  N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,
  N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,
  N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,
  N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,
  N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,
  N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,
  N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,
  N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258;
  wire [64:64] opA_r,opC_r,add1_out;
  wire [64:0] opA_mux,opB_mux,add2_out,opC_mux,opB_r,add1_in0,add1_in1,add2_in0;
  wire [1:0] opA_sel_lo;
  wire [3:0] opB_sel_lo,opC_sel_lo;
  wire [64:1] add2_in1;

  bsg_dff_en_width_p1
  req_reg
  (
    .clk_i(clk_i),
    .data_i(signed_div_i),
    .en_i(latch_signed_div_lo),
    .data_o(signed_div_r)
  );


  bsg_mux_one_hot_width_p65_els_p2
  muxA
  (
    .data_i({ divisor_msb, divisor_i, add1_out[64:64], add2_in1 }),
    .sel_one_hot_i(opA_sel_lo),
    .data_o(opA_mux)
  );


  bsg_mux_one_hot_width_p65_els_p4
  \genblk1.muxB 
  (
    .data_i({ opC_r[64:64], quotient_o, add1_out[64:64], add2_in1, add2_in1, opC_r[64:64], add2_out[63:0], quotient_o[63:63] }),
    .sel_one_hot_i(opB_sel_lo),
    .data_o(opB_mux)
  );


  bsg_mux_one_hot_width_p65_els_p4
  \genblk1.muxC 
  (
    .data_i({ dividend_msb, dividend_i, add1_out[64:64], add2_in1, quotient_o, _2_net__65_, quotient_o[62:0], _2_net__1_, _2_net__0_ }),
    .sel_one_hot_i(opC_sel_lo),
    .data_o(opC_mux)
  );


  bsg_dff_en_width_p65
  opA_reg
  (
    .clk_i(clk_i),
    .data_i(opA_mux),
    .en_i(opA_ld_lo),
    .data_o({ opA_r[64:64], remainder_o })
  );


  bsg_dff_en_width_p65
  opB_reg
  (
    .clk_i(clk_i),
    .data_i(opB_mux),
    .en_i(opB_ld_lo),
    .data_o(opB_r)
  );


  bsg_dff_en_width_p65
  opC_reg
  (
    .clk_i(clk_i),
    .data_i(opC_mux),
    .en_i(opC_ld_lo),
    .data_o({ opC_r[64:64], quotient_o })
  );


  bsg_adder_cin_width_p65
  adder1
  (
    .a_i(add1_in0),
    .b_i(add1_in1),
    .cin_i(adder1_cin_lo),
    .o({ add1_out[64:64], add2_in1 })
  );


  bsg_adder_cin_width_p65
  \genblk3.adder2 
  (
    .a_i(add2_in0),
    .b_i({ add2_in1, opC_r[64:64] }),
    .cin_i(\genblk3.adder2_cin ),
    .o(add2_out)
  );


  bsg_idiv_iterative_controller_64_2
  control
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_and_o(ready_and_o),
    .zero_divisor_i(zero_divisor_li),
    .signed_div_r_i(signed_div_r),
    .adder1_result_is_neg_i(add1_out[64]),
    .adder2_result_is_neg_i(add2_out[64]),
    .opA_is_neg_i(opA_r[64]),
    .opC_is_neg_i(opC_r[64]),
    .opA_sel_o(opA_sel_lo),
    .opA_ld_o(opA_ld_lo),
    .opA_inv_o(opA_inv_lo),
    .opA_clr_l_o(opA_clr_lo),
    .opB_sel_o(opB_sel_lo),
    .opB_ld_o(opB_ld_lo),
    .opB_inv_o(opB_inv_lo),
    .opB_clr_l_o(opB_clr_lo),
    .opC_sel_o(opC_sel_lo),
    .opC_ld_o(opC_ld_lo),
    .latch_signed_div_o(latch_signed_div_lo),
    .adder1_cin_o(adder1_cin_lo),
    .v_o(v_o),
    .yumi_i(yumi_i)
  );

  assign divisor_msb = signed_div_i & divisor_i[63];
  assign dividend_msb = signed_div_i & dividend_i[63];
  assign zero_divisor_li = ~N63;
  assign N63 = N62 | remainder_o[0];
  assign N62 = N61 | remainder_o[1];
  assign N61 = N60 | remainder_o[2];
  assign N60 = N59 | remainder_o[3];
  assign N59 = N58 | remainder_o[4];
  assign N58 = N57 | remainder_o[5];
  assign N57 = N56 | remainder_o[6];
  assign N56 = N55 | remainder_o[7];
  assign N55 = N54 | remainder_o[8];
  assign N54 = N53 | remainder_o[9];
  assign N53 = N52 | remainder_o[10];
  assign N52 = N51 | remainder_o[11];
  assign N51 = N50 | remainder_o[12];
  assign N50 = N49 | remainder_o[13];
  assign N49 = N48 | remainder_o[14];
  assign N48 = N47 | remainder_o[15];
  assign N47 = N46 | remainder_o[16];
  assign N46 = N45 | remainder_o[17];
  assign N45 = N44 | remainder_o[18];
  assign N44 = N43 | remainder_o[19];
  assign N43 = N42 | remainder_o[20];
  assign N42 = N41 | remainder_o[21];
  assign N41 = N40 | remainder_o[22];
  assign N40 = N39 | remainder_o[23];
  assign N39 = N38 | remainder_o[24];
  assign N38 = N37 | remainder_o[25];
  assign N37 = N36 | remainder_o[26];
  assign N36 = N35 | remainder_o[27];
  assign N35 = N34 | remainder_o[28];
  assign N34 = N33 | remainder_o[29];
  assign N33 = N32 | remainder_o[30];
  assign N32 = N31 | remainder_o[31];
  assign N31 = N30 | remainder_o[32];
  assign N30 = N29 | remainder_o[33];
  assign N29 = N28 | remainder_o[34];
  assign N28 = N27 | remainder_o[35];
  assign N27 = N26 | remainder_o[36];
  assign N26 = N25 | remainder_o[37];
  assign N25 = N24 | remainder_o[38];
  assign N24 = N23 | remainder_o[39];
  assign N23 = N22 | remainder_o[40];
  assign N22 = N21 | remainder_o[41];
  assign N21 = N20 | remainder_o[42];
  assign N20 = N19 | remainder_o[43];
  assign N19 = N18 | remainder_o[44];
  assign N18 = N17 | remainder_o[45];
  assign N17 = N16 | remainder_o[46];
  assign N16 = N15 | remainder_o[47];
  assign N15 = N14 | remainder_o[48];
  assign N14 = N13 | remainder_o[49];
  assign N13 = N12 | remainder_o[50];
  assign N12 = N11 | remainder_o[51];
  assign N11 = N10 | remainder_o[52];
  assign N10 = N9 | remainder_o[53];
  assign N9 = N8 | remainder_o[54];
  assign N8 = N7 | remainder_o[55];
  assign N7 = N6 | remainder_o[56];
  assign N6 = N5 | remainder_o[57];
  assign N5 = N4 | remainder_o[58];
  assign N4 = N3 | remainder_o[59];
  assign N3 = N2 | remainder_o[60];
  assign N2 = N1 | remainder_o[61];
  assign N1 = N0 | remainder_o[62];
  assign N0 = opA_r[64] | remainder_o[63];
  assign _2_net__65_ = ~add1_out[64];
  assign _2_net__1_ = ~add1_out[64];
  assign _2_net__0_ = ~add2_out[64];
  assign add1_in0[64] = N64 & opA_clr_lo;
  assign N64 = opA_r[64] ^ opA_inv_lo;
  assign add1_in0[63] = N65 & opA_clr_lo;
  assign N65 = remainder_o[63] ^ opA_inv_lo;
  assign add1_in0[62] = N66 & opA_clr_lo;
  assign N66 = remainder_o[62] ^ opA_inv_lo;
  assign add1_in0[61] = N67 & opA_clr_lo;
  assign N67 = remainder_o[61] ^ opA_inv_lo;
  assign add1_in0[60] = N68 & opA_clr_lo;
  assign N68 = remainder_o[60] ^ opA_inv_lo;
  assign add1_in0[59] = N69 & opA_clr_lo;
  assign N69 = remainder_o[59] ^ opA_inv_lo;
  assign add1_in0[58] = N70 & opA_clr_lo;
  assign N70 = remainder_o[58] ^ opA_inv_lo;
  assign add1_in0[57] = N71 & opA_clr_lo;
  assign N71 = remainder_o[57] ^ opA_inv_lo;
  assign add1_in0[56] = N72 & opA_clr_lo;
  assign N72 = remainder_o[56] ^ opA_inv_lo;
  assign add1_in0[55] = N73 & opA_clr_lo;
  assign N73 = remainder_o[55] ^ opA_inv_lo;
  assign add1_in0[54] = N74 & opA_clr_lo;
  assign N74 = remainder_o[54] ^ opA_inv_lo;
  assign add1_in0[53] = N75 & opA_clr_lo;
  assign N75 = remainder_o[53] ^ opA_inv_lo;
  assign add1_in0[52] = N76 & opA_clr_lo;
  assign N76 = remainder_o[52] ^ opA_inv_lo;
  assign add1_in0[51] = N77 & opA_clr_lo;
  assign N77 = remainder_o[51] ^ opA_inv_lo;
  assign add1_in0[50] = N78 & opA_clr_lo;
  assign N78 = remainder_o[50] ^ opA_inv_lo;
  assign add1_in0[49] = N79 & opA_clr_lo;
  assign N79 = remainder_o[49] ^ opA_inv_lo;
  assign add1_in0[48] = N80 & opA_clr_lo;
  assign N80 = remainder_o[48] ^ opA_inv_lo;
  assign add1_in0[47] = N81 & opA_clr_lo;
  assign N81 = remainder_o[47] ^ opA_inv_lo;
  assign add1_in0[46] = N82 & opA_clr_lo;
  assign N82 = remainder_o[46] ^ opA_inv_lo;
  assign add1_in0[45] = N83 & opA_clr_lo;
  assign N83 = remainder_o[45] ^ opA_inv_lo;
  assign add1_in0[44] = N84 & opA_clr_lo;
  assign N84 = remainder_o[44] ^ opA_inv_lo;
  assign add1_in0[43] = N85 & opA_clr_lo;
  assign N85 = remainder_o[43] ^ opA_inv_lo;
  assign add1_in0[42] = N86 & opA_clr_lo;
  assign N86 = remainder_o[42] ^ opA_inv_lo;
  assign add1_in0[41] = N87 & opA_clr_lo;
  assign N87 = remainder_o[41] ^ opA_inv_lo;
  assign add1_in0[40] = N88 & opA_clr_lo;
  assign N88 = remainder_o[40] ^ opA_inv_lo;
  assign add1_in0[39] = N89 & opA_clr_lo;
  assign N89 = remainder_o[39] ^ opA_inv_lo;
  assign add1_in0[38] = N90 & opA_clr_lo;
  assign N90 = remainder_o[38] ^ opA_inv_lo;
  assign add1_in0[37] = N91 & opA_clr_lo;
  assign N91 = remainder_o[37] ^ opA_inv_lo;
  assign add1_in0[36] = N92 & opA_clr_lo;
  assign N92 = remainder_o[36] ^ opA_inv_lo;
  assign add1_in0[35] = N93 & opA_clr_lo;
  assign N93 = remainder_o[35] ^ opA_inv_lo;
  assign add1_in0[34] = N94 & opA_clr_lo;
  assign N94 = remainder_o[34] ^ opA_inv_lo;
  assign add1_in0[33] = N95 & opA_clr_lo;
  assign N95 = remainder_o[33] ^ opA_inv_lo;
  assign add1_in0[32] = N96 & opA_clr_lo;
  assign N96 = remainder_o[32] ^ opA_inv_lo;
  assign add1_in0[31] = N97 & opA_clr_lo;
  assign N97 = remainder_o[31] ^ opA_inv_lo;
  assign add1_in0[30] = N98 & opA_clr_lo;
  assign N98 = remainder_o[30] ^ opA_inv_lo;
  assign add1_in0[29] = N99 & opA_clr_lo;
  assign N99 = remainder_o[29] ^ opA_inv_lo;
  assign add1_in0[28] = N100 & opA_clr_lo;
  assign N100 = remainder_o[28] ^ opA_inv_lo;
  assign add1_in0[27] = N101 & opA_clr_lo;
  assign N101 = remainder_o[27] ^ opA_inv_lo;
  assign add1_in0[26] = N102 & opA_clr_lo;
  assign N102 = remainder_o[26] ^ opA_inv_lo;
  assign add1_in0[25] = N103 & opA_clr_lo;
  assign N103 = remainder_o[25] ^ opA_inv_lo;
  assign add1_in0[24] = N104 & opA_clr_lo;
  assign N104 = remainder_o[24] ^ opA_inv_lo;
  assign add1_in0[23] = N105 & opA_clr_lo;
  assign N105 = remainder_o[23] ^ opA_inv_lo;
  assign add1_in0[22] = N106 & opA_clr_lo;
  assign N106 = remainder_o[22] ^ opA_inv_lo;
  assign add1_in0[21] = N107 & opA_clr_lo;
  assign N107 = remainder_o[21] ^ opA_inv_lo;
  assign add1_in0[20] = N108 & opA_clr_lo;
  assign N108 = remainder_o[20] ^ opA_inv_lo;
  assign add1_in0[19] = N109 & opA_clr_lo;
  assign N109 = remainder_o[19] ^ opA_inv_lo;
  assign add1_in0[18] = N110 & opA_clr_lo;
  assign N110 = remainder_o[18] ^ opA_inv_lo;
  assign add1_in0[17] = N111 & opA_clr_lo;
  assign N111 = remainder_o[17] ^ opA_inv_lo;
  assign add1_in0[16] = N112 & opA_clr_lo;
  assign N112 = remainder_o[16] ^ opA_inv_lo;
  assign add1_in0[15] = N113 & opA_clr_lo;
  assign N113 = remainder_o[15] ^ opA_inv_lo;
  assign add1_in0[14] = N114 & opA_clr_lo;
  assign N114 = remainder_o[14] ^ opA_inv_lo;
  assign add1_in0[13] = N115 & opA_clr_lo;
  assign N115 = remainder_o[13] ^ opA_inv_lo;
  assign add1_in0[12] = N116 & opA_clr_lo;
  assign N116 = remainder_o[12] ^ opA_inv_lo;
  assign add1_in0[11] = N117 & opA_clr_lo;
  assign N117 = remainder_o[11] ^ opA_inv_lo;
  assign add1_in0[10] = N118 & opA_clr_lo;
  assign N118 = remainder_o[10] ^ opA_inv_lo;
  assign add1_in0[9] = N119 & opA_clr_lo;
  assign N119 = remainder_o[9] ^ opA_inv_lo;
  assign add1_in0[8] = N120 & opA_clr_lo;
  assign N120 = remainder_o[8] ^ opA_inv_lo;
  assign add1_in0[7] = N121 & opA_clr_lo;
  assign N121 = remainder_o[7] ^ opA_inv_lo;
  assign add1_in0[6] = N122 & opA_clr_lo;
  assign N122 = remainder_o[6] ^ opA_inv_lo;
  assign add1_in0[5] = N123 & opA_clr_lo;
  assign N123 = remainder_o[5] ^ opA_inv_lo;
  assign add1_in0[4] = N124 & opA_clr_lo;
  assign N124 = remainder_o[4] ^ opA_inv_lo;
  assign add1_in0[3] = N125 & opA_clr_lo;
  assign N125 = remainder_o[3] ^ opA_inv_lo;
  assign add1_in0[2] = N126 & opA_clr_lo;
  assign N126 = remainder_o[2] ^ opA_inv_lo;
  assign add1_in0[1] = N127 & opA_clr_lo;
  assign N127 = remainder_o[1] ^ opA_inv_lo;
  assign add1_in0[0] = N128 & opA_clr_lo;
  assign N128 = remainder_o[0] ^ opA_inv_lo;
  assign add1_in1[64] = N129 & opB_clr_lo;
  assign N129 = opB_r[64] ^ opB_inv_lo;
  assign add1_in1[63] = N130 & opB_clr_lo;
  assign N130 = opB_r[63] ^ opB_inv_lo;
  assign add1_in1[62] = N131 & opB_clr_lo;
  assign N131 = opB_r[62] ^ opB_inv_lo;
  assign add1_in1[61] = N132 & opB_clr_lo;
  assign N132 = opB_r[61] ^ opB_inv_lo;
  assign add1_in1[60] = N133 & opB_clr_lo;
  assign N133 = opB_r[60] ^ opB_inv_lo;
  assign add1_in1[59] = N134 & opB_clr_lo;
  assign N134 = opB_r[59] ^ opB_inv_lo;
  assign add1_in1[58] = N135 & opB_clr_lo;
  assign N135 = opB_r[58] ^ opB_inv_lo;
  assign add1_in1[57] = N136 & opB_clr_lo;
  assign N136 = opB_r[57] ^ opB_inv_lo;
  assign add1_in1[56] = N137 & opB_clr_lo;
  assign N137 = opB_r[56] ^ opB_inv_lo;
  assign add1_in1[55] = N138 & opB_clr_lo;
  assign N138 = opB_r[55] ^ opB_inv_lo;
  assign add1_in1[54] = N139 & opB_clr_lo;
  assign N139 = opB_r[54] ^ opB_inv_lo;
  assign add1_in1[53] = N140 & opB_clr_lo;
  assign N140 = opB_r[53] ^ opB_inv_lo;
  assign add1_in1[52] = N141 & opB_clr_lo;
  assign N141 = opB_r[52] ^ opB_inv_lo;
  assign add1_in1[51] = N142 & opB_clr_lo;
  assign N142 = opB_r[51] ^ opB_inv_lo;
  assign add1_in1[50] = N143 & opB_clr_lo;
  assign N143 = opB_r[50] ^ opB_inv_lo;
  assign add1_in1[49] = N144 & opB_clr_lo;
  assign N144 = opB_r[49] ^ opB_inv_lo;
  assign add1_in1[48] = N145 & opB_clr_lo;
  assign N145 = opB_r[48] ^ opB_inv_lo;
  assign add1_in1[47] = N146 & opB_clr_lo;
  assign N146 = opB_r[47] ^ opB_inv_lo;
  assign add1_in1[46] = N147 & opB_clr_lo;
  assign N147 = opB_r[46] ^ opB_inv_lo;
  assign add1_in1[45] = N148 & opB_clr_lo;
  assign N148 = opB_r[45] ^ opB_inv_lo;
  assign add1_in1[44] = N149 & opB_clr_lo;
  assign N149 = opB_r[44] ^ opB_inv_lo;
  assign add1_in1[43] = N150 & opB_clr_lo;
  assign N150 = opB_r[43] ^ opB_inv_lo;
  assign add1_in1[42] = N151 & opB_clr_lo;
  assign N151 = opB_r[42] ^ opB_inv_lo;
  assign add1_in1[41] = N152 & opB_clr_lo;
  assign N152 = opB_r[41] ^ opB_inv_lo;
  assign add1_in1[40] = N153 & opB_clr_lo;
  assign N153 = opB_r[40] ^ opB_inv_lo;
  assign add1_in1[39] = N154 & opB_clr_lo;
  assign N154 = opB_r[39] ^ opB_inv_lo;
  assign add1_in1[38] = N155 & opB_clr_lo;
  assign N155 = opB_r[38] ^ opB_inv_lo;
  assign add1_in1[37] = N156 & opB_clr_lo;
  assign N156 = opB_r[37] ^ opB_inv_lo;
  assign add1_in1[36] = N157 & opB_clr_lo;
  assign N157 = opB_r[36] ^ opB_inv_lo;
  assign add1_in1[35] = N158 & opB_clr_lo;
  assign N158 = opB_r[35] ^ opB_inv_lo;
  assign add1_in1[34] = N159 & opB_clr_lo;
  assign N159 = opB_r[34] ^ opB_inv_lo;
  assign add1_in1[33] = N160 & opB_clr_lo;
  assign N160 = opB_r[33] ^ opB_inv_lo;
  assign add1_in1[32] = N161 & opB_clr_lo;
  assign N161 = opB_r[32] ^ opB_inv_lo;
  assign add1_in1[31] = N162 & opB_clr_lo;
  assign N162 = opB_r[31] ^ opB_inv_lo;
  assign add1_in1[30] = N163 & opB_clr_lo;
  assign N163 = opB_r[30] ^ opB_inv_lo;
  assign add1_in1[29] = N164 & opB_clr_lo;
  assign N164 = opB_r[29] ^ opB_inv_lo;
  assign add1_in1[28] = N165 & opB_clr_lo;
  assign N165 = opB_r[28] ^ opB_inv_lo;
  assign add1_in1[27] = N166 & opB_clr_lo;
  assign N166 = opB_r[27] ^ opB_inv_lo;
  assign add1_in1[26] = N167 & opB_clr_lo;
  assign N167 = opB_r[26] ^ opB_inv_lo;
  assign add1_in1[25] = N168 & opB_clr_lo;
  assign N168 = opB_r[25] ^ opB_inv_lo;
  assign add1_in1[24] = N169 & opB_clr_lo;
  assign N169 = opB_r[24] ^ opB_inv_lo;
  assign add1_in1[23] = N170 & opB_clr_lo;
  assign N170 = opB_r[23] ^ opB_inv_lo;
  assign add1_in1[22] = N171 & opB_clr_lo;
  assign N171 = opB_r[22] ^ opB_inv_lo;
  assign add1_in1[21] = N172 & opB_clr_lo;
  assign N172 = opB_r[21] ^ opB_inv_lo;
  assign add1_in1[20] = N173 & opB_clr_lo;
  assign N173 = opB_r[20] ^ opB_inv_lo;
  assign add1_in1[19] = N174 & opB_clr_lo;
  assign N174 = opB_r[19] ^ opB_inv_lo;
  assign add1_in1[18] = N175 & opB_clr_lo;
  assign N175 = opB_r[18] ^ opB_inv_lo;
  assign add1_in1[17] = N176 & opB_clr_lo;
  assign N176 = opB_r[17] ^ opB_inv_lo;
  assign add1_in1[16] = N177 & opB_clr_lo;
  assign N177 = opB_r[16] ^ opB_inv_lo;
  assign add1_in1[15] = N178 & opB_clr_lo;
  assign N178 = opB_r[15] ^ opB_inv_lo;
  assign add1_in1[14] = N179 & opB_clr_lo;
  assign N179 = opB_r[14] ^ opB_inv_lo;
  assign add1_in1[13] = N180 & opB_clr_lo;
  assign N180 = opB_r[13] ^ opB_inv_lo;
  assign add1_in1[12] = N181 & opB_clr_lo;
  assign N181 = opB_r[12] ^ opB_inv_lo;
  assign add1_in1[11] = N182 & opB_clr_lo;
  assign N182 = opB_r[11] ^ opB_inv_lo;
  assign add1_in1[10] = N183 & opB_clr_lo;
  assign N183 = opB_r[10] ^ opB_inv_lo;
  assign add1_in1[9] = N184 & opB_clr_lo;
  assign N184 = opB_r[9] ^ opB_inv_lo;
  assign add1_in1[8] = N185 & opB_clr_lo;
  assign N185 = opB_r[8] ^ opB_inv_lo;
  assign add1_in1[7] = N186 & opB_clr_lo;
  assign N186 = opB_r[7] ^ opB_inv_lo;
  assign add1_in1[6] = N187 & opB_clr_lo;
  assign N187 = opB_r[6] ^ opB_inv_lo;
  assign add1_in1[5] = N188 & opB_clr_lo;
  assign N188 = opB_r[5] ^ opB_inv_lo;
  assign add1_in1[4] = N189 & opB_clr_lo;
  assign N189 = opB_r[4] ^ opB_inv_lo;
  assign add1_in1[3] = N190 & opB_clr_lo;
  assign N190 = opB_r[3] ^ opB_inv_lo;
  assign add1_in1[2] = N191 & opB_clr_lo;
  assign N191 = opB_r[2] ^ opB_inv_lo;
  assign add1_in1[1] = N192 & opB_clr_lo;
  assign N192 = opB_r[1] ^ opB_inv_lo;
  assign add1_in1[0] = N193 & opB_clr_lo;
  assign N193 = opB_r[0] ^ opB_inv_lo;
  assign add2_in0[64] = opA_r[64] ^ N194;
  assign N194 = ~add1_out[64];
  assign add2_in0[63] = remainder_o[63] ^ N195;
  assign N195 = ~add1_out[64];
  assign add2_in0[62] = remainder_o[62] ^ N196;
  assign N196 = ~add1_out[64];
  assign add2_in0[61] = remainder_o[61] ^ N197;
  assign N197 = ~add1_out[64];
  assign add2_in0[60] = remainder_o[60] ^ N198;
  assign N198 = ~add1_out[64];
  assign add2_in0[59] = remainder_o[59] ^ N199;
  assign N199 = ~add1_out[64];
  assign add2_in0[58] = remainder_o[58] ^ N200;
  assign N200 = ~add1_out[64];
  assign add2_in0[57] = remainder_o[57] ^ N201;
  assign N201 = ~add1_out[64];
  assign add2_in0[56] = remainder_o[56] ^ N202;
  assign N202 = ~add1_out[64];
  assign add2_in0[55] = remainder_o[55] ^ N203;
  assign N203 = ~add1_out[64];
  assign add2_in0[54] = remainder_o[54] ^ N204;
  assign N204 = ~add1_out[64];
  assign add2_in0[53] = remainder_o[53] ^ N205;
  assign N205 = ~add1_out[64];
  assign add2_in0[52] = remainder_o[52] ^ N206;
  assign N206 = ~add1_out[64];
  assign add2_in0[51] = remainder_o[51] ^ N207;
  assign N207 = ~add1_out[64];
  assign add2_in0[50] = remainder_o[50] ^ N208;
  assign N208 = ~add1_out[64];
  assign add2_in0[49] = remainder_o[49] ^ N209;
  assign N209 = ~add1_out[64];
  assign add2_in0[48] = remainder_o[48] ^ N210;
  assign N210 = ~add1_out[64];
  assign add2_in0[47] = remainder_o[47] ^ N211;
  assign N211 = ~add1_out[64];
  assign add2_in0[46] = remainder_o[46] ^ N212;
  assign N212 = ~add1_out[64];
  assign add2_in0[45] = remainder_o[45] ^ N213;
  assign N213 = ~add1_out[64];
  assign add2_in0[44] = remainder_o[44] ^ N214;
  assign N214 = ~add1_out[64];
  assign add2_in0[43] = remainder_o[43] ^ N215;
  assign N215 = ~add1_out[64];
  assign add2_in0[42] = remainder_o[42] ^ N216;
  assign N216 = ~add1_out[64];
  assign add2_in0[41] = remainder_o[41] ^ N217;
  assign N217 = ~add1_out[64];
  assign add2_in0[40] = remainder_o[40] ^ N218;
  assign N218 = ~add1_out[64];
  assign add2_in0[39] = remainder_o[39] ^ N219;
  assign N219 = ~add1_out[64];
  assign add2_in0[38] = remainder_o[38] ^ N220;
  assign N220 = ~add1_out[64];
  assign add2_in0[37] = remainder_o[37] ^ N221;
  assign N221 = ~add1_out[64];
  assign add2_in0[36] = remainder_o[36] ^ N222;
  assign N222 = ~add1_out[64];
  assign add2_in0[35] = remainder_o[35] ^ N223;
  assign N223 = ~add1_out[64];
  assign add2_in0[34] = remainder_o[34] ^ N224;
  assign N224 = ~add1_out[64];
  assign add2_in0[33] = remainder_o[33] ^ N225;
  assign N225 = ~add1_out[64];
  assign add2_in0[32] = remainder_o[32] ^ N226;
  assign N226 = ~add1_out[64];
  assign add2_in0[31] = remainder_o[31] ^ N227;
  assign N227 = ~add1_out[64];
  assign add2_in0[30] = remainder_o[30] ^ N228;
  assign N228 = ~add1_out[64];
  assign add2_in0[29] = remainder_o[29] ^ N229;
  assign N229 = ~add1_out[64];
  assign add2_in0[28] = remainder_o[28] ^ N230;
  assign N230 = ~add1_out[64];
  assign add2_in0[27] = remainder_o[27] ^ N231;
  assign N231 = ~add1_out[64];
  assign add2_in0[26] = remainder_o[26] ^ N232;
  assign N232 = ~add1_out[64];
  assign add2_in0[25] = remainder_o[25] ^ N233;
  assign N233 = ~add1_out[64];
  assign add2_in0[24] = remainder_o[24] ^ N234;
  assign N234 = ~add1_out[64];
  assign add2_in0[23] = remainder_o[23] ^ N235;
  assign N235 = ~add1_out[64];
  assign add2_in0[22] = remainder_o[22] ^ N236;
  assign N236 = ~add1_out[64];
  assign add2_in0[21] = remainder_o[21] ^ N237;
  assign N237 = ~add1_out[64];
  assign add2_in0[20] = remainder_o[20] ^ N238;
  assign N238 = ~add1_out[64];
  assign add2_in0[19] = remainder_o[19] ^ N239;
  assign N239 = ~add1_out[64];
  assign add2_in0[18] = remainder_o[18] ^ N240;
  assign N240 = ~add1_out[64];
  assign add2_in0[17] = remainder_o[17] ^ N241;
  assign N241 = ~add1_out[64];
  assign add2_in0[16] = remainder_o[16] ^ N242;
  assign N242 = ~add1_out[64];
  assign add2_in0[15] = remainder_o[15] ^ N243;
  assign N243 = ~add1_out[64];
  assign add2_in0[14] = remainder_o[14] ^ N244;
  assign N244 = ~add1_out[64];
  assign add2_in0[13] = remainder_o[13] ^ N245;
  assign N245 = ~add1_out[64];
  assign add2_in0[12] = remainder_o[12] ^ N246;
  assign N246 = ~add1_out[64];
  assign add2_in0[11] = remainder_o[11] ^ N247;
  assign N247 = ~add1_out[64];
  assign add2_in0[10] = remainder_o[10] ^ N248;
  assign N248 = ~add1_out[64];
  assign add2_in0[9] = remainder_o[9] ^ N249;
  assign N249 = ~add1_out[64];
  assign add2_in0[8] = remainder_o[8] ^ N250;
  assign N250 = ~add1_out[64];
  assign add2_in0[7] = remainder_o[7] ^ N251;
  assign N251 = ~add1_out[64];
  assign add2_in0[6] = remainder_o[6] ^ N252;
  assign N252 = ~add1_out[64];
  assign add2_in0[5] = remainder_o[5] ^ N253;
  assign N253 = ~add1_out[64];
  assign add2_in0[4] = remainder_o[4] ^ N254;
  assign N254 = ~add1_out[64];
  assign add2_in0[3] = remainder_o[3] ^ N255;
  assign N255 = ~add1_out[64];
  assign add2_in0[2] = remainder_o[2] ^ N256;
  assign N256 = ~add1_out[64];
  assign add2_in0[1] = remainder_o[1] ^ N257;
  assign N257 = ~add1_out[64];
  assign add2_in0[0] = remainder_o[0] ^ N258;
  assign N258 = ~add1_out[64];
  assign \genblk3.adder2_cin  = ~add1_out[64];

endmodule



module bsg_dff_en_width_p13
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [12:0] data_i;
  output [12:0] data_o;
  input clk_i;
  input en_i;
  wire [12:0] data_o;
  reg data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,
  data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,
  data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mux_one_hot_width_p55_els_p5
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [274:0] data_i;
  input [4:0] sel_one_hot_i;
  output [54:0] data_o;
  wire [54:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164;
  wire [274:0] data_masked;
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[1];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[1];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[1];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[1];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[1];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[1];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[1];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[1];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[1];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[1];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[1];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[1];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[2];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[2];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[2];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[2];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[2];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[2];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[2];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[2];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[2];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[2];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[2];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[2];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[2];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[2];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[2];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[2];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[2];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[2];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[2];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[2];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[2];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[2];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[2];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[2];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[2];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[2];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[2];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[2];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[2];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[2];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[2];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[2];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[2];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[2];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[2];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[2];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[2];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[2];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[2];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[2];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[2];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[2];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[2];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[2];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[2];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[2];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[2];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[2];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[2];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[2];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[2];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[2];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[2];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[2];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[2];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[3];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[3];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[3];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[3];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[3];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[3];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[3];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[3];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[3];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[3];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[3];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[3];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[3];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[3];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[3];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[3];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[3];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[3];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[3];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[3];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[3];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[3];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[3];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[3];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[3];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[3];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[3];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[3];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[3];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[3];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[3];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[3];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[3];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[3];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[3];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[3];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[3];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[3];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[3];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[3];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[3];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[3];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[3];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[3];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[3];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[3];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[3];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[3];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[3];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[3];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[3];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[3];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[3];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[3];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[3];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[4];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[4];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[4];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[4];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[4];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[4];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[4];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[4];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[4];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[4];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[4];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[4];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[4];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[4];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[4];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[4];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[4];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[4];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[4];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[4];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[4];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[4];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[4];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[4];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[4];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[4];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[4];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[4];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[4];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[4];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[4];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[4];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[4];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[4];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[4];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[4];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[4];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[4];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[4];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[4];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[4];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[4];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[4];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[4];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[4];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[4];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[4];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[4];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[4];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[4];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[4];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[4];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[4];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[4];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[4];
  assign data_o[0] = N2 | data_masked[0];
  assign N2 = N1 | data_masked[55];
  assign N1 = N0 | data_masked[110];
  assign N0 = data_masked[220] | data_masked[165];
  assign data_o[1] = N5 | data_masked[1];
  assign N5 = N4 | data_masked[56];
  assign N4 = N3 | data_masked[111];
  assign N3 = data_masked[221] | data_masked[166];
  assign data_o[2] = N8 | data_masked[2];
  assign N8 = N7 | data_masked[57];
  assign N7 = N6 | data_masked[112];
  assign N6 = data_masked[222] | data_masked[167];
  assign data_o[3] = N11 | data_masked[3];
  assign N11 = N10 | data_masked[58];
  assign N10 = N9 | data_masked[113];
  assign N9 = data_masked[223] | data_masked[168];
  assign data_o[4] = N14 | data_masked[4];
  assign N14 = N13 | data_masked[59];
  assign N13 = N12 | data_masked[114];
  assign N12 = data_masked[224] | data_masked[169];
  assign data_o[5] = N17 | data_masked[5];
  assign N17 = N16 | data_masked[60];
  assign N16 = N15 | data_masked[115];
  assign N15 = data_masked[225] | data_masked[170];
  assign data_o[6] = N20 | data_masked[6];
  assign N20 = N19 | data_masked[61];
  assign N19 = N18 | data_masked[116];
  assign N18 = data_masked[226] | data_masked[171];
  assign data_o[7] = N23 | data_masked[7];
  assign N23 = N22 | data_masked[62];
  assign N22 = N21 | data_masked[117];
  assign N21 = data_masked[227] | data_masked[172];
  assign data_o[8] = N26 | data_masked[8];
  assign N26 = N25 | data_masked[63];
  assign N25 = N24 | data_masked[118];
  assign N24 = data_masked[228] | data_masked[173];
  assign data_o[9] = N29 | data_masked[9];
  assign N29 = N28 | data_masked[64];
  assign N28 = N27 | data_masked[119];
  assign N27 = data_masked[229] | data_masked[174];
  assign data_o[10] = N32 | data_masked[10];
  assign N32 = N31 | data_masked[65];
  assign N31 = N30 | data_masked[120];
  assign N30 = data_masked[230] | data_masked[175];
  assign data_o[11] = N35 | data_masked[11];
  assign N35 = N34 | data_masked[66];
  assign N34 = N33 | data_masked[121];
  assign N33 = data_masked[231] | data_masked[176];
  assign data_o[12] = N38 | data_masked[12];
  assign N38 = N37 | data_masked[67];
  assign N37 = N36 | data_masked[122];
  assign N36 = data_masked[232] | data_masked[177];
  assign data_o[13] = N41 | data_masked[13];
  assign N41 = N40 | data_masked[68];
  assign N40 = N39 | data_masked[123];
  assign N39 = data_masked[233] | data_masked[178];
  assign data_o[14] = N44 | data_masked[14];
  assign N44 = N43 | data_masked[69];
  assign N43 = N42 | data_masked[124];
  assign N42 = data_masked[234] | data_masked[179];
  assign data_o[15] = N47 | data_masked[15];
  assign N47 = N46 | data_masked[70];
  assign N46 = N45 | data_masked[125];
  assign N45 = data_masked[235] | data_masked[180];
  assign data_o[16] = N50 | data_masked[16];
  assign N50 = N49 | data_masked[71];
  assign N49 = N48 | data_masked[126];
  assign N48 = data_masked[236] | data_masked[181];
  assign data_o[17] = N53 | data_masked[17];
  assign N53 = N52 | data_masked[72];
  assign N52 = N51 | data_masked[127];
  assign N51 = data_masked[237] | data_masked[182];
  assign data_o[18] = N56 | data_masked[18];
  assign N56 = N55 | data_masked[73];
  assign N55 = N54 | data_masked[128];
  assign N54 = data_masked[238] | data_masked[183];
  assign data_o[19] = N59 | data_masked[19];
  assign N59 = N58 | data_masked[74];
  assign N58 = N57 | data_masked[129];
  assign N57 = data_masked[239] | data_masked[184];
  assign data_o[20] = N62 | data_masked[20];
  assign N62 = N61 | data_masked[75];
  assign N61 = N60 | data_masked[130];
  assign N60 = data_masked[240] | data_masked[185];
  assign data_o[21] = N65 | data_masked[21];
  assign N65 = N64 | data_masked[76];
  assign N64 = N63 | data_masked[131];
  assign N63 = data_masked[241] | data_masked[186];
  assign data_o[22] = N68 | data_masked[22];
  assign N68 = N67 | data_masked[77];
  assign N67 = N66 | data_masked[132];
  assign N66 = data_masked[242] | data_masked[187];
  assign data_o[23] = N71 | data_masked[23];
  assign N71 = N70 | data_masked[78];
  assign N70 = N69 | data_masked[133];
  assign N69 = data_masked[243] | data_masked[188];
  assign data_o[24] = N74 | data_masked[24];
  assign N74 = N73 | data_masked[79];
  assign N73 = N72 | data_masked[134];
  assign N72 = data_masked[244] | data_masked[189];
  assign data_o[25] = N77 | data_masked[25];
  assign N77 = N76 | data_masked[80];
  assign N76 = N75 | data_masked[135];
  assign N75 = data_masked[245] | data_masked[190];
  assign data_o[26] = N80 | data_masked[26];
  assign N80 = N79 | data_masked[81];
  assign N79 = N78 | data_masked[136];
  assign N78 = data_masked[246] | data_masked[191];
  assign data_o[27] = N83 | data_masked[27];
  assign N83 = N82 | data_masked[82];
  assign N82 = N81 | data_masked[137];
  assign N81 = data_masked[247] | data_masked[192];
  assign data_o[28] = N86 | data_masked[28];
  assign N86 = N85 | data_masked[83];
  assign N85 = N84 | data_masked[138];
  assign N84 = data_masked[248] | data_masked[193];
  assign data_o[29] = N89 | data_masked[29];
  assign N89 = N88 | data_masked[84];
  assign N88 = N87 | data_masked[139];
  assign N87 = data_masked[249] | data_masked[194];
  assign data_o[30] = N92 | data_masked[30];
  assign N92 = N91 | data_masked[85];
  assign N91 = N90 | data_masked[140];
  assign N90 = data_masked[250] | data_masked[195];
  assign data_o[31] = N95 | data_masked[31];
  assign N95 = N94 | data_masked[86];
  assign N94 = N93 | data_masked[141];
  assign N93 = data_masked[251] | data_masked[196];
  assign data_o[32] = N98 | data_masked[32];
  assign N98 = N97 | data_masked[87];
  assign N97 = N96 | data_masked[142];
  assign N96 = data_masked[252] | data_masked[197];
  assign data_o[33] = N101 | data_masked[33];
  assign N101 = N100 | data_masked[88];
  assign N100 = N99 | data_masked[143];
  assign N99 = data_masked[253] | data_masked[198];
  assign data_o[34] = N104 | data_masked[34];
  assign N104 = N103 | data_masked[89];
  assign N103 = N102 | data_masked[144];
  assign N102 = data_masked[254] | data_masked[199];
  assign data_o[35] = N107 | data_masked[35];
  assign N107 = N106 | data_masked[90];
  assign N106 = N105 | data_masked[145];
  assign N105 = data_masked[255] | data_masked[200];
  assign data_o[36] = N110 | data_masked[36];
  assign N110 = N109 | data_masked[91];
  assign N109 = N108 | data_masked[146];
  assign N108 = data_masked[256] | data_masked[201];
  assign data_o[37] = N113 | data_masked[37];
  assign N113 = N112 | data_masked[92];
  assign N112 = N111 | data_masked[147];
  assign N111 = data_masked[257] | data_masked[202];
  assign data_o[38] = N116 | data_masked[38];
  assign N116 = N115 | data_masked[93];
  assign N115 = N114 | data_masked[148];
  assign N114 = data_masked[258] | data_masked[203];
  assign data_o[39] = N119 | data_masked[39];
  assign N119 = N118 | data_masked[94];
  assign N118 = N117 | data_masked[149];
  assign N117 = data_masked[259] | data_masked[204];
  assign data_o[40] = N122 | data_masked[40];
  assign N122 = N121 | data_masked[95];
  assign N121 = N120 | data_masked[150];
  assign N120 = data_masked[260] | data_masked[205];
  assign data_o[41] = N125 | data_masked[41];
  assign N125 = N124 | data_masked[96];
  assign N124 = N123 | data_masked[151];
  assign N123 = data_masked[261] | data_masked[206];
  assign data_o[42] = N128 | data_masked[42];
  assign N128 = N127 | data_masked[97];
  assign N127 = N126 | data_masked[152];
  assign N126 = data_masked[262] | data_masked[207];
  assign data_o[43] = N131 | data_masked[43];
  assign N131 = N130 | data_masked[98];
  assign N130 = N129 | data_masked[153];
  assign N129 = data_masked[263] | data_masked[208];
  assign data_o[44] = N134 | data_masked[44];
  assign N134 = N133 | data_masked[99];
  assign N133 = N132 | data_masked[154];
  assign N132 = data_masked[264] | data_masked[209];
  assign data_o[45] = N137 | data_masked[45];
  assign N137 = N136 | data_masked[100];
  assign N136 = N135 | data_masked[155];
  assign N135 = data_masked[265] | data_masked[210];
  assign data_o[46] = N140 | data_masked[46];
  assign N140 = N139 | data_masked[101];
  assign N139 = N138 | data_masked[156];
  assign N138 = data_masked[266] | data_masked[211];
  assign data_o[47] = N143 | data_masked[47];
  assign N143 = N142 | data_masked[102];
  assign N142 = N141 | data_masked[157];
  assign N141 = data_masked[267] | data_masked[212];
  assign data_o[48] = N146 | data_masked[48];
  assign N146 = N145 | data_masked[103];
  assign N145 = N144 | data_masked[158];
  assign N144 = data_masked[268] | data_masked[213];
  assign data_o[49] = N149 | data_masked[49];
  assign N149 = N148 | data_masked[104];
  assign N148 = N147 | data_masked[159];
  assign N147 = data_masked[269] | data_masked[214];
  assign data_o[50] = N152 | data_masked[50];
  assign N152 = N151 | data_masked[105];
  assign N151 = N150 | data_masked[160];
  assign N150 = data_masked[270] | data_masked[215];
  assign data_o[51] = N155 | data_masked[51];
  assign N155 = N154 | data_masked[106];
  assign N154 = N153 | data_masked[161];
  assign N153 = data_masked[271] | data_masked[216];
  assign data_o[52] = N158 | data_masked[52];
  assign N158 = N157 | data_masked[107];
  assign N157 = N156 | data_masked[162];
  assign N156 = data_masked[272] | data_masked[217];
  assign data_o[53] = N161 | data_masked[53];
  assign N161 = N160 | data_masked[108];
  assign N160 = N159 | data_masked[163];
  assign N159 = data_masked[273] | data_masked[218];
  assign data_o[54] = N164 | data_masked[54];
  assign N164 = N163 | data_masked[109];
  assign N163 = N162 | data_masked[164];
  assign N162 = data_masked[274] | data_masked[219];

endmodule



module bsg_mux_one_hot_width_p55_els_p4
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [219:0] data_i;
  input [3:0] sel_one_hot_i;
  output [54:0] data_o;
  wire [54:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109;
  wire [219:0] data_masked;
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[1];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[1];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[1];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[1];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[1];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[1];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[1];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[1];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[1];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[1];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[1];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[1];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[2];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[2];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[2];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[2];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[2];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[2];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[2];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[2];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[2];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[2];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[2];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[2];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[2];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[2];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[2];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[2];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[2];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[2];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[2];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[2];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[2];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[2];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[2];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[2];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[2];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[2];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[2];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[2];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[2];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[2];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[2];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[2];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[2];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[2];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[2];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[2];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[2];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[2];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[2];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[2];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[2];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[2];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[2];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[2];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[2];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[2];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[2];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[2];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[2];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[2];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[2];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[2];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[2];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[2];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[2];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[3];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[3];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[3];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[3];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[3];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[3];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[3];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[3];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[3];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[3];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[3];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[3];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[3];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[3];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[3];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[3];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[3];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[3];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[3];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[3];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[3];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[3];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[3];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[3];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[3];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[3];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[3];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[3];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[3];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[3];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[3];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[3];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[3];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[3];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[3];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[3];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[3];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[3];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[3];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[3];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[3];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[3];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[3];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[3];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[3];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[3];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[3];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[3];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[3];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[3];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[3];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[3];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[3];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[3];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[3];
  assign data_o[0] = N1 | data_masked[0];
  assign N1 = N0 | data_masked[55];
  assign N0 = data_masked[165] | data_masked[110];
  assign data_o[1] = N3 | data_masked[1];
  assign N3 = N2 | data_masked[56];
  assign N2 = data_masked[166] | data_masked[111];
  assign data_o[2] = N5 | data_masked[2];
  assign N5 = N4 | data_masked[57];
  assign N4 = data_masked[167] | data_masked[112];
  assign data_o[3] = N7 | data_masked[3];
  assign N7 = N6 | data_masked[58];
  assign N6 = data_masked[168] | data_masked[113];
  assign data_o[4] = N9 | data_masked[4];
  assign N9 = N8 | data_masked[59];
  assign N8 = data_masked[169] | data_masked[114];
  assign data_o[5] = N11 | data_masked[5];
  assign N11 = N10 | data_masked[60];
  assign N10 = data_masked[170] | data_masked[115];
  assign data_o[6] = N13 | data_masked[6];
  assign N13 = N12 | data_masked[61];
  assign N12 = data_masked[171] | data_masked[116];
  assign data_o[7] = N15 | data_masked[7];
  assign N15 = N14 | data_masked[62];
  assign N14 = data_masked[172] | data_masked[117];
  assign data_o[8] = N17 | data_masked[8];
  assign N17 = N16 | data_masked[63];
  assign N16 = data_masked[173] | data_masked[118];
  assign data_o[9] = N19 | data_masked[9];
  assign N19 = N18 | data_masked[64];
  assign N18 = data_masked[174] | data_masked[119];
  assign data_o[10] = N21 | data_masked[10];
  assign N21 = N20 | data_masked[65];
  assign N20 = data_masked[175] | data_masked[120];
  assign data_o[11] = N23 | data_masked[11];
  assign N23 = N22 | data_masked[66];
  assign N22 = data_masked[176] | data_masked[121];
  assign data_o[12] = N25 | data_masked[12];
  assign N25 = N24 | data_masked[67];
  assign N24 = data_masked[177] | data_masked[122];
  assign data_o[13] = N27 | data_masked[13];
  assign N27 = N26 | data_masked[68];
  assign N26 = data_masked[178] | data_masked[123];
  assign data_o[14] = N29 | data_masked[14];
  assign N29 = N28 | data_masked[69];
  assign N28 = data_masked[179] | data_masked[124];
  assign data_o[15] = N31 | data_masked[15];
  assign N31 = N30 | data_masked[70];
  assign N30 = data_masked[180] | data_masked[125];
  assign data_o[16] = N33 | data_masked[16];
  assign N33 = N32 | data_masked[71];
  assign N32 = data_masked[181] | data_masked[126];
  assign data_o[17] = N35 | data_masked[17];
  assign N35 = N34 | data_masked[72];
  assign N34 = data_masked[182] | data_masked[127];
  assign data_o[18] = N37 | data_masked[18];
  assign N37 = N36 | data_masked[73];
  assign N36 = data_masked[183] | data_masked[128];
  assign data_o[19] = N39 | data_masked[19];
  assign N39 = N38 | data_masked[74];
  assign N38 = data_masked[184] | data_masked[129];
  assign data_o[20] = N41 | data_masked[20];
  assign N41 = N40 | data_masked[75];
  assign N40 = data_masked[185] | data_masked[130];
  assign data_o[21] = N43 | data_masked[21];
  assign N43 = N42 | data_masked[76];
  assign N42 = data_masked[186] | data_masked[131];
  assign data_o[22] = N45 | data_masked[22];
  assign N45 = N44 | data_masked[77];
  assign N44 = data_masked[187] | data_masked[132];
  assign data_o[23] = N47 | data_masked[23];
  assign N47 = N46 | data_masked[78];
  assign N46 = data_masked[188] | data_masked[133];
  assign data_o[24] = N49 | data_masked[24];
  assign N49 = N48 | data_masked[79];
  assign N48 = data_masked[189] | data_masked[134];
  assign data_o[25] = N51 | data_masked[25];
  assign N51 = N50 | data_masked[80];
  assign N50 = data_masked[190] | data_masked[135];
  assign data_o[26] = N53 | data_masked[26];
  assign N53 = N52 | data_masked[81];
  assign N52 = data_masked[191] | data_masked[136];
  assign data_o[27] = N55 | data_masked[27];
  assign N55 = N54 | data_masked[82];
  assign N54 = data_masked[192] | data_masked[137];
  assign data_o[28] = N57 | data_masked[28];
  assign N57 = N56 | data_masked[83];
  assign N56 = data_masked[193] | data_masked[138];
  assign data_o[29] = N59 | data_masked[29];
  assign N59 = N58 | data_masked[84];
  assign N58 = data_masked[194] | data_masked[139];
  assign data_o[30] = N61 | data_masked[30];
  assign N61 = N60 | data_masked[85];
  assign N60 = data_masked[195] | data_masked[140];
  assign data_o[31] = N63 | data_masked[31];
  assign N63 = N62 | data_masked[86];
  assign N62 = data_masked[196] | data_masked[141];
  assign data_o[32] = N65 | data_masked[32];
  assign N65 = N64 | data_masked[87];
  assign N64 = data_masked[197] | data_masked[142];
  assign data_o[33] = N67 | data_masked[33];
  assign N67 = N66 | data_masked[88];
  assign N66 = data_masked[198] | data_masked[143];
  assign data_o[34] = N69 | data_masked[34];
  assign N69 = N68 | data_masked[89];
  assign N68 = data_masked[199] | data_masked[144];
  assign data_o[35] = N71 | data_masked[35];
  assign N71 = N70 | data_masked[90];
  assign N70 = data_masked[200] | data_masked[145];
  assign data_o[36] = N73 | data_masked[36];
  assign N73 = N72 | data_masked[91];
  assign N72 = data_masked[201] | data_masked[146];
  assign data_o[37] = N75 | data_masked[37];
  assign N75 = N74 | data_masked[92];
  assign N74 = data_masked[202] | data_masked[147];
  assign data_o[38] = N77 | data_masked[38];
  assign N77 = N76 | data_masked[93];
  assign N76 = data_masked[203] | data_masked[148];
  assign data_o[39] = N79 | data_masked[39];
  assign N79 = N78 | data_masked[94];
  assign N78 = data_masked[204] | data_masked[149];
  assign data_o[40] = N81 | data_masked[40];
  assign N81 = N80 | data_masked[95];
  assign N80 = data_masked[205] | data_masked[150];
  assign data_o[41] = N83 | data_masked[41];
  assign N83 = N82 | data_masked[96];
  assign N82 = data_masked[206] | data_masked[151];
  assign data_o[42] = N85 | data_masked[42];
  assign N85 = N84 | data_masked[97];
  assign N84 = data_masked[207] | data_masked[152];
  assign data_o[43] = N87 | data_masked[43];
  assign N87 = N86 | data_masked[98];
  assign N86 = data_masked[208] | data_masked[153];
  assign data_o[44] = N89 | data_masked[44];
  assign N89 = N88 | data_masked[99];
  assign N88 = data_masked[209] | data_masked[154];
  assign data_o[45] = N91 | data_masked[45];
  assign N91 = N90 | data_masked[100];
  assign N90 = data_masked[210] | data_masked[155];
  assign data_o[46] = N93 | data_masked[46];
  assign N93 = N92 | data_masked[101];
  assign N92 = data_masked[211] | data_masked[156];
  assign data_o[47] = N95 | data_masked[47];
  assign N95 = N94 | data_masked[102];
  assign N94 = data_masked[212] | data_masked[157];
  assign data_o[48] = N97 | data_masked[48];
  assign N97 = N96 | data_masked[103];
  assign N96 = data_masked[213] | data_masked[158];
  assign data_o[49] = N99 | data_masked[49];
  assign N99 = N98 | data_masked[104];
  assign N98 = data_masked[214] | data_masked[159];
  assign data_o[50] = N101 | data_masked[50];
  assign N101 = N100 | data_masked[105];
  assign N100 = data_masked[215] | data_masked[160];
  assign data_o[51] = N103 | data_masked[51];
  assign N103 = N102 | data_masked[106];
  assign N102 = data_masked[216] | data_masked[161];
  assign data_o[52] = N105 | data_masked[52];
  assign N105 = N104 | data_masked[107];
  assign N104 = data_masked[217] | data_masked[162];
  assign data_o[53] = N107 | data_masked[53];
  assign N107 = N106 | data_masked[108];
  assign N106 = data_masked[218] | data_masked[163];
  assign data_o[54] = N109 | data_masked[54];
  assign N109 = N108 | data_masked[109];
  assign N108 = data_masked[219] | data_masked[164];

endmodule



module divSqrtRecFNToRaw_medium_expWidth11_sigWidth53_options0
(
  nReset,
  clock,
  control,
  inReady,
  inValid,
  sqrtOp,
  a,
  b,
  roundingMode,
  outValid,
  sqrtOpOut,
  roundingModeOut,
  invalidExc,
  infiniteExc,
  out_isNaN,
  out_isInf,
  out_isZero,
  out_sign,
  out_sExp,
  out_sig
);

  input [0:0] control;
  input [64:0] a;
  input [64:0] b;
  input [2:0] roundingMode;
  output [2:0] roundingModeOut;
  output [12:0] out_sExp;
  output [55:0] out_sig;
  input nReset;
  input clock;
  input inValid;
  input sqrtOp;
  output inReady;
  output outValid;
  output sqrtOpOut;
  output invalidExc;
  output infiniteExc;
  output out_isNaN;
  output out_isInf;
  output out_isZero;
  output out_sign;
  wire [2:0] roundingModeOut;
  wire [12:0] out_sExp,sExpA_S,sExpB_S;
  wire [55:0] out_sig;
  wire inReady,outValid,sqrtOpOut,invalidExc,infiniteExc,out_isNaN,out_isInf,
  out_isZero,out_sign,N0,N1,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,isNaNA_S,isInfA_S,isZeroA_S,signA_S,isSigNaNA_S,isNaNB_S,isInfB_S,
  isZeroB_S,signB_S,isSigNaNB_S,notSigNaNIn_invalidExc_S_div,
  notSigNaNIn_invalidExc_S_sqrt,N24,N25,majorExc_S,N26,N27,isNaN_S,N28,isInf_S,N29,isZero_S,N30,sign_S,
  specialCaseA_S,specialCaseB_S,normalCase_S_div,normalCase_S_sqrt,normalCase_S,
  N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,evenSqrt_S,oddSqrt_S,entering,
  entering_normalCase,skipCycle2,N44,step1Case,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,
  N74,majorExc_Z,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,
  N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,
  N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,
  N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,
  N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,
  N157,N158,N159,N160,trialTermMuxIn_0__53_,trialTermMuxIn_0__52_,
  trialTermMuxIn_0__51_,trialTermMuxIn_0__50_,trialTermMuxIn_0__49_,trialTermMuxIn_0__48_,
  trialTermMuxIn_0__47_,trialTermMuxIn_0__46_,trialTermMuxIn_0__45_,trialTermMuxIn_0__44_,
  trialTermMuxIn_0__43_,trialTermMuxIn_0__42_,trialTermMuxIn_0__41_,
  trialTermMuxIn_0__40_,trialTermMuxIn_0__39_,trialTermMuxIn_0__38_,trialTermMuxIn_0__37_,
  trialTermMuxIn_0__36_,trialTermMuxIn_0__35_,trialTermMuxIn_0__34_,
  trialTermMuxIn_0__33_,trialTermMuxIn_0__32_,trialTermMuxIn_0__31_,trialTermMuxIn_0__30_,
  trialTermMuxIn_0__29_,trialTermMuxIn_0__28_,trialTermMuxIn_0__27_,trialTermMuxIn_0__26_,
  trialTermMuxIn_0__25_,trialTermMuxIn_0__24_,trialTermMuxIn_0__23_,
  trialTermMuxIn_0__22_,trialTermMuxIn_0__21_,trialTermMuxIn_0__20_,trialTermMuxIn_0__19_,
  trialTermMuxIn_0__18_,trialTermMuxIn_0__17_,trialTermMuxIn_0__16_,trialTermMuxIn_0__15_,
  trialTermMuxIn_0__14_,trialTermMuxIn_0__13_,trialTermMuxIn_0__12_,
  trialTermMuxIn_0__11_,trialTermMuxIn_0__10_,trialTermMuxIn_0__9_,trialTermMuxIn_0__8_,
  trialTermMuxIn_0__7_,trialTermMuxIn_0__6_,trialTermMuxIn_0__5_,trialTermMuxIn_0__4_,
  trialTermMuxIn_0__3_,trialTermMuxIn_0__2_,trialTermMuxIn_0__1_,N161,N162,N163,N164,
  N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,
  N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
  N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,
  N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,
  N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,
  N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,
  N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,newBit2,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,sigX_NMuxIn_3__54_,sigX_NMuxIn_0__53_,sigX_NMuxIn_0__52_,
  sigX_NMuxIn_0__51_,sigX_NMuxIn_0__50_,sigX_NMuxIn_0__49_,sigX_NMuxIn_0__48_,
  sigX_NMuxIn_0__47_,sigX_NMuxIn_0__46_,sigX_NMuxIn_0__45_,sigX_NMuxIn_0__44_,sigX_NMuxIn_0__43_,
  sigX_NMuxIn_0__42_,sigX_NMuxIn_0__41_,sigX_NMuxIn_0__40_,sigX_NMuxIn_0__39_,
  sigX_NMuxIn_0__38_,sigX_NMuxIn_0__37_,sigX_NMuxIn_0__36_,sigX_NMuxIn_0__35_,
  sigX_NMuxIn_0__34_,sigX_NMuxIn_0__33_,sigX_NMuxIn_0__32_,sigX_NMuxIn_0__31_,
  sigX_NMuxIn_0__30_,sigX_NMuxIn_0__29_,sigX_NMuxIn_0__28_,sigX_NMuxIn_0__27_,
  sigX_NMuxIn_0__26_,sigX_NMuxIn_0__25_,sigX_NMuxIn_0__24_,sigX_NMuxIn_0__23_,sigX_NMuxIn_0__22_,
  sigX_NMuxIn_0__21_,sigX_NMuxIn_0__20_,sigX_NMuxIn_0__19_,sigX_NMuxIn_0__18_,
  sigX_NMuxIn_0__17_,sigX_NMuxIn_0__16_,sigX_NMuxIn_0__15_,sigX_NMuxIn_0__14_,
  sigX_NMuxIn_0__13_,sigX_NMuxIn_0__12_,sigX_NMuxIn_0__11_,sigX_NMuxIn_0__10_,
  sigX_NMuxIn_0__9_,sigX_NMuxIn_0__8_,sigX_NMuxIn_0__7_,sigX_NMuxIn_0__6_,sigX_NMuxIn_0__5_,
  sigX_NMuxIn_0__4_,sigX_NMuxIn_0__3_,sigX_NMuxIn_0__2_,sigX_NMuxIn_0__1_,
  sigX_NMuxIn_0__0_,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,
  N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,
  N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,
  N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,
  N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,
  N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,
  N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,
  N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N2,N449,N450,N451,
  N452,N453,N454,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,
  N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,
  N485,N486,N487,N488,N489,N490,N491,N492,sv2v_dc_1,sv2v_dc_2;
  wire [53:0] sigA_S,sigB_S,bitMask,sigXNext;
  wire [13:0] sExpQuot_S_div;
  wire [12:9] sSatExpQuot_S_div;
  wire [5:0] cycleNum;
  wire [51:0] fractB_Z;
  wire [1:0] decHiSigA_S;
  wire [55:1] rem,remNext;
  wire [54:0] rem_Z,trialTerm,trialTermNext,sigX_N;
  wire [4:0] trialTermSel;
  wire [56:0] trialRem1,trialRem2;
  wire [0:0] sigX_NSel;
  reg cycleNum_5_sv2v_reg,cycleNum_4_sv2v_reg,cycleNum_3_sv2v_reg,cycleNum_2_sv2v_reg,
  cycleNum_1_sv2v_reg,cycleNum_0_sv2v_reg,fractB_Z_51_sv2v_reg,
  fractB_Z_50_sv2v_reg,fractB_Z_49_sv2v_reg,fractB_Z_48_sv2v_reg,fractB_Z_47_sv2v_reg,
  fractB_Z_46_sv2v_reg,fractB_Z_45_sv2v_reg,fractB_Z_44_sv2v_reg,fractB_Z_43_sv2v_reg,
  fractB_Z_42_sv2v_reg,fractB_Z_41_sv2v_reg,fractB_Z_40_sv2v_reg,fractB_Z_39_sv2v_reg,
  fractB_Z_38_sv2v_reg,fractB_Z_37_sv2v_reg,fractB_Z_36_sv2v_reg,fractB_Z_35_sv2v_reg,
  fractB_Z_34_sv2v_reg,fractB_Z_33_sv2v_reg,fractB_Z_32_sv2v_reg,
  fractB_Z_31_sv2v_reg,fractB_Z_30_sv2v_reg,fractB_Z_29_sv2v_reg,fractB_Z_28_sv2v_reg,
  fractB_Z_27_sv2v_reg,fractB_Z_26_sv2v_reg,fractB_Z_25_sv2v_reg,fractB_Z_24_sv2v_reg,
  fractB_Z_23_sv2v_reg,fractB_Z_22_sv2v_reg,fractB_Z_21_sv2v_reg,fractB_Z_20_sv2v_reg,
  fractB_Z_19_sv2v_reg,fractB_Z_18_sv2v_reg,fractB_Z_17_sv2v_reg,fractB_Z_16_sv2v_reg,
  fractB_Z_15_sv2v_reg,fractB_Z_14_sv2v_reg,fractB_Z_13_sv2v_reg,fractB_Z_12_sv2v_reg,
  fractB_Z_11_sv2v_reg,fractB_Z_10_sv2v_reg,fractB_Z_9_sv2v_reg,
  fractB_Z_8_sv2v_reg,fractB_Z_7_sv2v_reg,fractB_Z_6_sv2v_reg,fractB_Z_5_sv2v_reg,
  fractB_Z_4_sv2v_reg,fractB_Z_3_sv2v_reg,fractB_Z_2_sv2v_reg,fractB_Z_1_sv2v_reg,
  fractB_Z_0_sv2v_reg,sqrtOpOut_sv2v_reg,majorExc_Z_sv2v_reg,out_isNaN_sv2v_reg,out_isInf_sv2v_reg,
  out_isZero_sv2v_reg,out_sign_sv2v_reg,out_sExp_12_sv2v_reg,out_sExp_11_sv2v_reg,
  out_sExp_10_sv2v_reg,out_sExp_9_sv2v_reg,out_sExp_8_sv2v_reg,out_sExp_7_sv2v_reg,
  out_sExp_6_sv2v_reg,out_sExp_5_sv2v_reg,out_sExp_4_sv2v_reg,out_sExp_3_sv2v_reg,
  out_sExp_2_sv2v_reg,out_sExp_1_sv2v_reg,out_sExp_0_sv2v_reg,
  roundingModeOut_2_sv2v_reg,roundingModeOut_1_sv2v_reg,roundingModeOut_0_sv2v_reg,out_sig_0_sv2v_reg,
  rem_Z_54_sv2v_reg,rem_Z_53_sv2v_reg,rem_Z_52_sv2v_reg,rem_Z_51_sv2v_reg,
  rem_Z_50_sv2v_reg,rem_Z_49_sv2v_reg,rem_Z_48_sv2v_reg,rem_Z_47_sv2v_reg,
  rem_Z_46_sv2v_reg,rem_Z_45_sv2v_reg,rem_Z_44_sv2v_reg,rem_Z_43_sv2v_reg,rem_Z_42_sv2v_reg,
  rem_Z_41_sv2v_reg,rem_Z_40_sv2v_reg,rem_Z_39_sv2v_reg,rem_Z_38_sv2v_reg,
  rem_Z_37_sv2v_reg,rem_Z_36_sv2v_reg,rem_Z_35_sv2v_reg,rem_Z_34_sv2v_reg,rem_Z_33_sv2v_reg,
  rem_Z_32_sv2v_reg,rem_Z_31_sv2v_reg,rem_Z_30_sv2v_reg,rem_Z_29_sv2v_reg,
  rem_Z_28_sv2v_reg,rem_Z_27_sv2v_reg,rem_Z_26_sv2v_reg,rem_Z_25_sv2v_reg,rem_Z_24_sv2v_reg,
  rem_Z_23_sv2v_reg,rem_Z_22_sv2v_reg,rem_Z_21_sv2v_reg,rem_Z_20_sv2v_reg,
  rem_Z_19_sv2v_reg,rem_Z_18_sv2v_reg,rem_Z_17_sv2v_reg,rem_Z_16_sv2v_reg,rem_Z_15_sv2v_reg,
  rem_Z_14_sv2v_reg,rem_Z_13_sv2v_reg,rem_Z_12_sv2v_reg,rem_Z_11_sv2v_reg,
  rem_Z_10_sv2v_reg,rem_Z_9_sv2v_reg,rem_Z_8_sv2v_reg,rem_Z_7_sv2v_reg,rem_Z_6_sv2v_reg,
  rem_Z_5_sv2v_reg,rem_Z_4_sv2v_reg,rem_Z_3_sv2v_reg,rem_Z_2_sv2v_reg,
  rem_Z_1_sv2v_reg,rem_Z_0_sv2v_reg,out_sig_55_sv2v_reg,out_sig_54_sv2v_reg,out_sig_53_sv2v_reg,
  out_sig_52_sv2v_reg,out_sig_51_sv2v_reg,out_sig_50_sv2v_reg,out_sig_49_sv2v_reg,
  out_sig_48_sv2v_reg,out_sig_47_sv2v_reg,out_sig_46_sv2v_reg,out_sig_45_sv2v_reg,
  out_sig_44_sv2v_reg,out_sig_43_sv2v_reg,out_sig_42_sv2v_reg,out_sig_41_sv2v_reg,
  out_sig_40_sv2v_reg,out_sig_39_sv2v_reg,out_sig_38_sv2v_reg,out_sig_37_sv2v_reg,
  out_sig_36_sv2v_reg,out_sig_35_sv2v_reg,out_sig_34_sv2v_reg,out_sig_33_sv2v_reg,
  out_sig_32_sv2v_reg,out_sig_31_sv2v_reg,out_sig_30_sv2v_reg,out_sig_29_sv2v_reg,
  out_sig_28_sv2v_reg,out_sig_27_sv2v_reg,out_sig_26_sv2v_reg,out_sig_25_sv2v_reg,
  out_sig_24_sv2v_reg,out_sig_23_sv2v_reg,out_sig_22_sv2v_reg,out_sig_21_sv2v_reg,
  out_sig_20_sv2v_reg,out_sig_19_sv2v_reg,out_sig_18_sv2v_reg,out_sig_17_sv2v_reg,
  out_sig_16_sv2v_reg,out_sig_15_sv2v_reg,out_sig_14_sv2v_reg,out_sig_13_sv2v_reg,
  out_sig_12_sv2v_reg,out_sig_11_sv2v_reg,out_sig_10_sv2v_reg,out_sig_9_sv2v_reg,
  out_sig_8_sv2v_reg,out_sig_7_sv2v_reg,out_sig_6_sv2v_reg,out_sig_5_sv2v_reg,
  out_sig_4_sv2v_reg,out_sig_3_sv2v_reg,out_sig_2_sv2v_reg,out_sig_1_sv2v_reg;
  assign cycleNum[5] = cycleNum_5_sv2v_reg;
  assign cycleNum[4] = cycleNum_4_sv2v_reg;
  assign cycleNum[3] = cycleNum_3_sv2v_reg;
  assign cycleNum[2] = cycleNum_2_sv2v_reg;
  assign cycleNum[1] = cycleNum_1_sv2v_reg;
  assign cycleNum[0] = cycleNum_0_sv2v_reg;
  assign fractB_Z[51] = fractB_Z_51_sv2v_reg;
  assign fractB_Z[50] = fractB_Z_50_sv2v_reg;
  assign fractB_Z[49] = fractB_Z_49_sv2v_reg;
  assign fractB_Z[48] = fractB_Z_48_sv2v_reg;
  assign fractB_Z[47] = fractB_Z_47_sv2v_reg;
  assign fractB_Z[46] = fractB_Z_46_sv2v_reg;
  assign fractB_Z[45] = fractB_Z_45_sv2v_reg;
  assign fractB_Z[44] = fractB_Z_44_sv2v_reg;
  assign fractB_Z[43] = fractB_Z_43_sv2v_reg;
  assign fractB_Z[42] = fractB_Z_42_sv2v_reg;
  assign fractB_Z[41] = fractB_Z_41_sv2v_reg;
  assign fractB_Z[40] = fractB_Z_40_sv2v_reg;
  assign fractB_Z[39] = fractB_Z_39_sv2v_reg;
  assign fractB_Z[38] = fractB_Z_38_sv2v_reg;
  assign fractB_Z[37] = fractB_Z_37_sv2v_reg;
  assign fractB_Z[36] = fractB_Z_36_sv2v_reg;
  assign fractB_Z[35] = fractB_Z_35_sv2v_reg;
  assign fractB_Z[34] = fractB_Z_34_sv2v_reg;
  assign fractB_Z[33] = fractB_Z_33_sv2v_reg;
  assign fractB_Z[32] = fractB_Z_32_sv2v_reg;
  assign fractB_Z[31] = fractB_Z_31_sv2v_reg;
  assign fractB_Z[30] = fractB_Z_30_sv2v_reg;
  assign fractB_Z[29] = fractB_Z_29_sv2v_reg;
  assign fractB_Z[28] = fractB_Z_28_sv2v_reg;
  assign fractB_Z[27] = fractB_Z_27_sv2v_reg;
  assign fractB_Z[26] = fractB_Z_26_sv2v_reg;
  assign fractB_Z[25] = fractB_Z_25_sv2v_reg;
  assign fractB_Z[24] = fractB_Z_24_sv2v_reg;
  assign fractB_Z[23] = fractB_Z_23_sv2v_reg;
  assign fractB_Z[22] = fractB_Z_22_sv2v_reg;
  assign fractB_Z[21] = fractB_Z_21_sv2v_reg;
  assign fractB_Z[20] = fractB_Z_20_sv2v_reg;
  assign fractB_Z[19] = fractB_Z_19_sv2v_reg;
  assign fractB_Z[18] = fractB_Z_18_sv2v_reg;
  assign fractB_Z[17] = fractB_Z_17_sv2v_reg;
  assign fractB_Z[16] = fractB_Z_16_sv2v_reg;
  assign fractB_Z[15] = fractB_Z_15_sv2v_reg;
  assign fractB_Z[14] = fractB_Z_14_sv2v_reg;
  assign fractB_Z[13] = fractB_Z_13_sv2v_reg;
  assign fractB_Z[12] = fractB_Z_12_sv2v_reg;
  assign fractB_Z[11] = fractB_Z_11_sv2v_reg;
  assign fractB_Z[10] = fractB_Z_10_sv2v_reg;
  assign fractB_Z[9] = fractB_Z_9_sv2v_reg;
  assign fractB_Z[8] = fractB_Z_8_sv2v_reg;
  assign fractB_Z[7] = fractB_Z_7_sv2v_reg;
  assign fractB_Z[6] = fractB_Z_6_sv2v_reg;
  assign fractB_Z[5] = fractB_Z_5_sv2v_reg;
  assign fractB_Z[4] = fractB_Z_4_sv2v_reg;
  assign fractB_Z[3] = fractB_Z_3_sv2v_reg;
  assign fractB_Z[2] = fractB_Z_2_sv2v_reg;
  assign fractB_Z[1] = fractB_Z_1_sv2v_reg;
  assign fractB_Z[0] = fractB_Z_0_sv2v_reg;
  assign sqrtOpOut = sqrtOpOut_sv2v_reg;
  assign majorExc_Z = majorExc_Z_sv2v_reg;
  assign out_isNaN = out_isNaN_sv2v_reg;
  assign out_isInf = out_isInf_sv2v_reg;
  assign out_isZero = out_isZero_sv2v_reg;
  assign out_sign = out_sign_sv2v_reg;
  assign out_sExp[12] = out_sExp_12_sv2v_reg;
  assign out_sExp[11] = out_sExp_11_sv2v_reg;
  assign out_sExp[10] = out_sExp_10_sv2v_reg;
  assign out_sExp[9] = out_sExp_9_sv2v_reg;
  assign out_sExp[8] = out_sExp_8_sv2v_reg;
  assign out_sExp[7] = out_sExp_7_sv2v_reg;
  assign out_sExp[6] = out_sExp_6_sv2v_reg;
  assign out_sExp[5] = out_sExp_5_sv2v_reg;
  assign out_sExp[4] = out_sExp_4_sv2v_reg;
  assign out_sExp[3] = out_sExp_3_sv2v_reg;
  assign out_sExp[2] = out_sExp_2_sv2v_reg;
  assign out_sExp[1] = out_sExp_1_sv2v_reg;
  assign out_sExp[0] = out_sExp_0_sv2v_reg;
  assign roundingModeOut[2] = roundingModeOut_2_sv2v_reg;
  assign roundingModeOut[1] = roundingModeOut_1_sv2v_reg;
  assign roundingModeOut[0] = roundingModeOut_0_sv2v_reg;
  assign out_sig[0] = out_sig_0_sv2v_reg;
  assign rem_Z[54] = rem_Z_54_sv2v_reg;
  assign rem_Z[53] = rem_Z_53_sv2v_reg;
  assign rem_Z[52] = rem_Z_52_sv2v_reg;
  assign rem_Z[51] = rem_Z_51_sv2v_reg;
  assign rem_Z[50] = rem_Z_50_sv2v_reg;
  assign rem_Z[49] = rem_Z_49_sv2v_reg;
  assign rem_Z[48] = rem_Z_48_sv2v_reg;
  assign rem_Z[47] = rem_Z_47_sv2v_reg;
  assign rem_Z[46] = rem_Z_46_sv2v_reg;
  assign rem_Z[45] = rem_Z_45_sv2v_reg;
  assign rem_Z[44] = rem_Z_44_sv2v_reg;
  assign rem_Z[43] = rem_Z_43_sv2v_reg;
  assign rem_Z[42] = rem_Z_42_sv2v_reg;
  assign rem_Z[41] = rem_Z_41_sv2v_reg;
  assign rem_Z[40] = rem_Z_40_sv2v_reg;
  assign rem_Z[39] = rem_Z_39_sv2v_reg;
  assign rem_Z[38] = rem_Z_38_sv2v_reg;
  assign rem_Z[37] = rem_Z_37_sv2v_reg;
  assign rem_Z[36] = rem_Z_36_sv2v_reg;
  assign rem_Z[35] = rem_Z_35_sv2v_reg;
  assign rem_Z[34] = rem_Z_34_sv2v_reg;
  assign rem_Z[33] = rem_Z_33_sv2v_reg;
  assign rem_Z[32] = rem_Z_32_sv2v_reg;
  assign rem_Z[31] = rem_Z_31_sv2v_reg;
  assign rem_Z[30] = rem_Z_30_sv2v_reg;
  assign rem_Z[29] = rem_Z_29_sv2v_reg;
  assign rem_Z[28] = rem_Z_28_sv2v_reg;
  assign rem_Z[27] = rem_Z_27_sv2v_reg;
  assign rem_Z[26] = rem_Z_26_sv2v_reg;
  assign rem_Z[25] = rem_Z_25_sv2v_reg;
  assign rem_Z[24] = rem_Z_24_sv2v_reg;
  assign rem_Z[23] = rem_Z_23_sv2v_reg;
  assign rem_Z[22] = rem_Z_22_sv2v_reg;
  assign rem_Z[21] = rem_Z_21_sv2v_reg;
  assign rem_Z[20] = rem_Z_20_sv2v_reg;
  assign rem_Z[19] = rem_Z_19_sv2v_reg;
  assign rem_Z[18] = rem_Z_18_sv2v_reg;
  assign rem_Z[17] = rem_Z_17_sv2v_reg;
  assign rem_Z[16] = rem_Z_16_sv2v_reg;
  assign rem_Z[15] = rem_Z_15_sv2v_reg;
  assign rem_Z[14] = rem_Z_14_sv2v_reg;
  assign rem_Z[13] = rem_Z_13_sv2v_reg;
  assign rem_Z[12] = rem_Z_12_sv2v_reg;
  assign rem_Z[11] = rem_Z_11_sv2v_reg;
  assign rem_Z[10] = rem_Z_10_sv2v_reg;
  assign rem_Z[9] = rem_Z_9_sv2v_reg;
  assign rem_Z[8] = rem_Z_8_sv2v_reg;
  assign rem_Z[7] = rem_Z_7_sv2v_reg;
  assign rem_Z[6] = rem_Z_6_sv2v_reg;
  assign rem_Z[5] = rem_Z_5_sv2v_reg;
  assign rem_Z[4] = rem_Z_4_sv2v_reg;
  assign rem_Z[3] = rem_Z_3_sv2v_reg;
  assign rem_Z[2] = rem_Z_2_sv2v_reg;
  assign rem_Z[1] = rem_Z_1_sv2v_reg;
  assign rem_Z[0] = rem_Z_0_sv2v_reg;
  assign out_sig[55] = out_sig_55_sv2v_reg;
  assign out_sig[54] = out_sig_54_sv2v_reg;
  assign out_sig[53] = out_sig_53_sv2v_reg;
  assign out_sig[52] = out_sig_52_sv2v_reg;
  assign out_sig[51] = out_sig_51_sv2v_reg;
  assign out_sig[50] = out_sig_50_sv2v_reg;
  assign out_sig[49] = out_sig_49_sv2v_reg;
  assign out_sig[48] = out_sig_48_sv2v_reg;
  assign out_sig[47] = out_sig_47_sv2v_reg;
  assign out_sig[46] = out_sig_46_sv2v_reg;
  assign out_sig[45] = out_sig_45_sv2v_reg;
  assign out_sig[44] = out_sig_44_sv2v_reg;
  assign out_sig[43] = out_sig_43_sv2v_reg;
  assign out_sig[42] = out_sig_42_sv2v_reg;
  assign out_sig[41] = out_sig_41_sv2v_reg;
  assign out_sig[40] = out_sig_40_sv2v_reg;
  assign out_sig[39] = out_sig_39_sv2v_reg;
  assign out_sig[38] = out_sig_38_sv2v_reg;
  assign out_sig[37] = out_sig_37_sv2v_reg;
  assign out_sig[36] = out_sig_36_sv2v_reg;
  assign out_sig[35] = out_sig_35_sv2v_reg;
  assign out_sig[34] = out_sig_34_sv2v_reg;
  assign out_sig[33] = out_sig_33_sv2v_reg;
  assign out_sig[32] = out_sig_32_sv2v_reg;
  assign out_sig[31] = out_sig_31_sv2v_reg;
  assign out_sig[30] = out_sig_30_sv2v_reg;
  assign out_sig[29] = out_sig_29_sv2v_reg;
  assign out_sig[28] = out_sig_28_sv2v_reg;
  assign out_sig[27] = out_sig_27_sv2v_reg;
  assign out_sig[26] = out_sig_26_sv2v_reg;
  assign out_sig[25] = out_sig_25_sv2v_reg;
  assign out_sig[24] = out_sig_24_sv2v_reg;
  assign out_sig[23] = out_sig_23_sv2v_reg;
  assign out_sig[22] = out_sig_22_sv2v_reg;
  assign out_sig[21] = out_sig_21_sv2v_reg;
  assign out_sig[20] = out_sig_20_sv2v_reg;
  assign out_sig[19] = out_sig_19_sv2v_reg;
  assign out_sig[18] = out_sig_18_sv2v_reg;
  assign out_sig[17] = out_sig_17_sv2v_reg;
  assign out_sig[16] = out_sig_16_sv2v_reg;
  assign out_sig[15] = out_sig_15_sv2v_reg;
  assign out_sig[14] = out_sig_14_sv2v_reg;
  assign out_sig[13] = out_sig_13_sv2v_reg;
  assign out_sig[12] = out_sig_12_sv2v_reg;
  assign out_sig[11] = out_sig_11_sv2v_reg;
  assign out_sig[10] = out_sig_10_sv2v_reg;
  assign out_sig[9] = out_sig_9_sv2v_reg;
  assign out_sig[8] = out_sig_8_sv2v_reg;
  assign out_sig[7] = out_sig_7_sv2v_reg;
  assign out_sig[6] = out_sig_6_sv2v_reg;
  assign out_sig[5] = out_sig_5_sv2v_reg;
  assign out_sig[4] = out_sig_4_sv2v_reg;
  assign out_sig[3] = out_sig_3_sv2v_reg;
  assign out_sig[2] = out_sig_2_sv2v_reg;
  assign out_sig[1] = out_sig_1_sv2v_reg;

  recFNToRawFN_expWidth11_sigWidth53
  recFNToRawFN_a
  (
    .in(a),
    .isNaN(isNaNA_S),
    .isInf(isInfA_S),
    .isZero(isZeroA_S),
    .sign(signA_S),
    .sExp(sExpA_S),
    .sig(sigA_S)
  );


  isSigNaNRecFN_expWidth11_sigWidth53
  isSigNaN_a
  (
    .in(a),
    .isSigNaN(isSigNaNA_S)
  );


  recFNToRawFN_expWidth11_sigWidth53
  recFNToRawFN_b
  (
    .in(b),
    .isNaN(isNaNB_S),
    .isInf(isInfB_S),
    .isZero(isZeroB_S),
    .sign(signB_S),
    .sExp(sExpB_S),
    .sig(sigB_S)
  );


  isSigNaNRecFN_expWidth11_sigWidth53
  isSigNaN_b
  (
    .in(b),
    .isSigNaN(isSigNaNB_S)
  );

  assign N42 = $signed({ 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) <= $signed(sExpQuot_S_div);
  assign inReady = cycleNum <= 1'b1;
  assign N44 = cycleNum <= { 1'b1, 1'b0 };
  assign { bitMask, sv2v_dc_1, sv2v_dc_2 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << cycleNum;

  bsg_mux_one_hot_width_p55_els_p5
  trialTerm_mux
  (
    .data_i({ sigB_S, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, fractB_Z, 1'b0, out_sig[54:54], trialTermMuxIn_0__53_, trialTermMuxIn_0__52_, trialTermMuxIn_0__51_, trialTermMuxIn_0__50_, trialTermMuxIn_0__49_, trialTermMuxIn_0__48_, trialTermMuxIn_0__47_, trialTermMuxIn_0__46_, trialTermMuxIn_0__45_, trialTermMuxIn_0__44_, trialTermMuxIn_0__43_, trialTermMuxIn_0__42_, trialTermMuxIn_0__41_, trialTermMuxIn_0__40_, trialTermMuxIn_0__39_, trialTermMuxIn_0__38_, trialTermMuxIn_0__37_, trialTermMuxIn_0__36_, trialTermMuxIn_0__35_, trialTermMuxIn_0__34_, trialTermMuxIn_0__33_, trialTermMuxIn_0__32_, trialTermMuxIn_0__31_, trialTermMuxIn_0__30_, trialTermMuxIn_0__29_, trialTermMuxIn_0__28_, trialTermMuxIn_0__27_, trialTermMuxIn_0__26_, trialTermMuxIn_0__25_, trialTermMuxIn_0__24_, trialTermMuxIn_0__23_, trialTermMuxIn_0__22_, trialTermMuxIn_0__21_, trialTermMuxIn_0__20_, trialTermMuxIn_0__19_, trialTermMuxIn_0__18_, trialTermMuxIn_0__17_, trialTermMuxIn_0__16_, trialTermMuxIn_0__15_, trialTermMuxIn_0__14_, trialTermMuxIn_0__13_, trialTermMuxIn_0__12_, trialTermMuxIn_0__11_, trialTermMuxIn_0__10_, trialTermMuxIn_0__9_, trialTermMuxIn_0__8_, trialTermMuxIn_0__7_, trialTermMuxIn_0__6_, trialTermMuxIn_0__5_, trialTermMuxIn_0__4_, trialTermMuxIn_0__3_, trialTermMuxIn_0__2_, trialTermMuxIn_0__1_, bitMask[0:0] }),
    .sel_one_hot_i(trialTermSel),
    .data_o(trialTerm)
  );

  assign sigX_NMuxIn_3__54_ = $signed(1'b0) <= $signed(trialRem1);
  assign newBit2 = $signed(1'b0) <= $signed(trialRem2);

  bsg_mux_one_hot_width_p55_els_p4
  sigX_N_mux
  (
    .data_i({ sigX_NMuxIn_3__54_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, sigX_NMuxIn_3__54_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, out_sig[55:55], sigX_NMuxIn_0__53_, sigX_NMuxIn_0__52_, sigX_NMuxIn_0__51_, sigX_NMuxIn_0__50_, sigX_NMuxIn_0__49_, sigX_NMuxIn_0__48_, sigX_NMuxIn_0__47_, sigX_NMuxIn_0__46_, sigX_NMuxIn_0__45_, sigX_NMuxIn_0__44_, sigX_NMuxIn_0__43_, sigX_NMuxIn_0__42_, sigX_NMuxIn_0__41_, sigX_NMuxIn_0__40_, sigX_NMuxIn_0__39_, sigX_NMuxIn_0__38_, sigX_NMuxIn_0__37_, sigX_NMuxIn_0__36_, sigX_NMuxIn_0__35_, sigX_NMuxIn_0__34_, sigX_NMuxIn_0__33_, sigX_NMuxIn_0__32_, sigX_NMuxIn_0__31_, sigX_NMuxIn_0__30_, sigX_NMuxIn_0__29_, sigX_NMuxIn_0__28_, sigX_NMuxIn_0__27_, sigX_NMuxIn_0__26_, sigX_NMuxIn_0__25_, sigX_NMuxIn_0__24_, sigX_NMuxIn_0__23_, sigX_NMuxIn_0__22_, sigX_NMuxIn_0__21_, sigX_NMuxIn_0__20_, sigX_NMuxIn_0__19_, sigX_NMuxIn_0__18_, sigX_NMuxIn_0__17_, sigX_NMuxIn_0__16_, sigX_NMuxIn_0__15_, sigX_NMuxIn_0__14_, sigX_NMuxIn_0__13_, sigX_NMuxIn_0__12_, sigX_NMuxIn_0__11_, sigX_NMuxIn_0__10_, sigX_NMuxIn_0__9_, sigX_NMuxIn_0__8_, sigX_NMuxIn_0__7_, sigX_NMuxIn_0__6_, sigX_NMuxIn_0__5_, sigX_NMuxIn_0__4_, sigX_NMuxIn_0__3_, sigX_NMuxIn_0__2_, sigX_NMuxIn_0__1_, sigX_NMuxIn_0__0_ }),
    .sel_one_hot_i({ trialTermSel[4:2], sigX_NSel[0:0] }),
    .data_o(sigX_N)
  );

  assign N326 = cycleNum > { 1'b1, 1'b0 };
  assign N444 = $signed(trialRem1) != $signed(1'b0);
  assign N445 = $signed(trialRem2) != $signed(1'b0);
  assign N449 = ~cycleNum[0];
  assign N450 = cycleNum[4] | cycleNum[5];
  assign N451 = cycleNum[3] | N450;
  assign N452 = cycleNum[2] | N451;
  assign N453 = cycleNum[1] | N452;
  assign N454 = N449 | N453;
  assign outValid = ~N454;
  assign N456 = ~cycleNum[2];
  assign N457 = cycleNum[4] | cycleNum[5];
  assign N458 = cycleNum[3] | N457;
  assign N459 = N456 | N458;
  assign N460 = cycleNum[1] | N459;
  assign N461 = cycleNum[0] | N460;
  assign N462 = ~N461;
  assign N463 = cycleNum[4] | cycleNum[5];
  assign N464 = cycleNum[3] | N463;
  assign N465 = cycleNum[2] | N464;
  assign N466 = cycleNum[1] | N465;
  assign N467 = cycleNum[0] | N466;
  assign N468 = ~N467;
  assign sExpQuot_S_div = sExpA_S + { sExpB_S[11:11], sExpB_S[11:11], sExpB_S[11:11], N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41 };
  assign decHiSigA_S = sigA_S[52:51] - 1'b1;
  assign trialRem1 = { rem, 1'b0 } - trialTerm;
  assign { N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77 } = $signed(sExpA_S[12:1]) + $signed({ 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 });
  assign { N61, N60, N59, N58, N57, N56 } = cycleNum - { N55, step1Case };
  assign trialRem2 = { remNext, 1'b0 } - trialTermNext;
  assign majorExc_S = (N0)? N25 : 
                      (N1)? N26 : 1'b0;
  assign N0 = sqrtOp;
  assign N1 = N24;
  assign isNaN_S = (N0)? N27 : 
                   (N1)? N28 : 1'b0;
  assign isInf_S = (N0)? isInfA_S : 
                   (N1)? N29 : 1'b0;
  assign isZero_S = (N0)? isZeroA_S : 
                    (N1)? N30 : 1'b0;
  assign normalCase_S = (N0)? normalCase_S_sqrt : 
                        (N1)? normalCase_S_div : 1'b0;
  assign sSatExpQuot_S_div = (N3)? { 1'b0, 1'b1, 1'b1, 1'b0 } : 
                             (N43)? sExpQuot_S_div[12:9] : 1'b0;
  assign N3 = N42;
  assign N50 = ~sExpA_S[0];
  assign { N52, N51 } = (N0)? { N50, sExpA_S[0:0] } : 
                        (N1)? { 1'b1, 1'b1 } : 1'b0;
  assign { N54, N53 } = (N4)? { N52, N51 } : 
                        (N5)? { 1'b0, 1'b0 } : 1'b0;
  assign N4 = entering_normalCase;
  assign N5 = N49;
  assign { N67, N66, N65, N64, N63, N62 } = (N6)? { N61, N60, N59, N58, N57, N56 } : 
                                            (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N6 = N467;
  assign N7 = N468;
  assign N73 = (N8)? 1'b1 : 
               (N2)? 1'b0 : 1'b0;
  assign N8 = N46;
  assign { N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90 } = (N0)? { N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77 } : 
                                                                                  (N1)? { sSatExpQuot_S_div, sExpQuot_S_div[8:0] } : 1'b0;
  assign { N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106 } = (N9)? { decHiSigA_S, sigA_S[50:0], 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                        (N10)? { 1'b0, sigA_S } : 1'b0;
  assign N9 = oddSqrt_S;
  assign N10 = N105;
  assign rem = (N11)? { N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106 } : 
               (N12)? rem_Z : 1'b0;
  assign N11 = inReady;
  assign N12 = N104;
  assign { N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163 } = (N13)? bitMask : 
                                                                                                                                                                                                                                                                                                                                                  (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = N162;
  assign N14 = N161;
  assign trialTermNext = (N15)? { sigXNext[53:53], N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, bitMask[1:1] } : 
                         (N16)? trialTerm : 1'b0;
  assign N15 = sqrtOpOut;
  assign N16 = N489;
  assign remNext = (N17)? trialRem1[54:0] : 
                   (N18)? { rem[54:1], 1'b0 } : 1'b0;
  assign N17 = N271;
  assign N18 = N270;
  assign { N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273 } = (N19)? bitMask[53:1] : 
                                                                                                                                                                                                                                                                                                                                            (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N19 = newBit2;
  assign N20 = N272;
  assign { N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333 } = (N21)? trialRem1[54:0] : 
                                                                                                                                                                                                                                                                                                                                                        (N22)? { rem[54:1], 1'b0 } : 1'b0;
  assign N21 = N332;
  assign N22 = N331;
  assign { N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388 } = (N23)? { N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333 } : 
                                                                                                                                                                                                                                                                                                                                                        (N448)? trialRem2[54:0] : 
                                                                                                                                                                                                                                                                                                                                                        (N330)? { remNext[54:1], 1'b0 } : 1'b0;
  assign N23 = N328;
  assign notSigNaNIn_invalidExc_S_div = N469 | N470;
  assign N469 = isZeroA_S & isZeroB_S;
  assign N470 = isInfA_S & isInfB_S;
  assign notSigNaNIn_invalidExc_S_sqrt = N473 & signA_S;
  assign N473 = N471 & N472;
  assign N471 = ~isNaNA_S;
  assign N472 = ~isZeroA_S;
  assign N24 = ~sqrtOp;
  assign N25 = isSigNaNA_S | notSigNaNIn_invalidExc_S_sqrt;
  assign N26 = N475 | N478;
  assign N475 = N474 | notSigNaNIn_invalidExc_S_div;
  assign N474 = isSigNaNA_S | isSigNaNB_S;
  assign N478 = N477 & isZeroB_S;
  assign N477 = N471 & N476;
  assign N476 = ~isInfA_S;
  assign N27 = isNaNA_S | notSigNaNIn_invalidExc_S_sqrt;
  assign N28 = N479 | notSigNaNIn_invalidExc_S_div;
  assign N479 = isNaNA_S | isNaNB_S;
  assign N29 = isInfA_S | isZeroB_S;
  assign N30 = isZeroA_S | isInfB_S;
  assign sign_S = signA_S ^ N480;
  assign N480 = N24 & signB_S;
  assign specialCaseA_S = N481 | isZeroA_S;
  assign N481 = isNaNA_S | isInfA_S;
  assign specialCaseB_S = N482 | isZeroB_S;
  assign N482 = isNaNB_S | isInfB_S;
  assign normalCase_S_div = N483 & N484;
  assign N483 = ~specialCaseA_S;
  assign N484 = ~specialCaseB_S;
  assign normalCase_S_sqrt = N483 & N485;
  assign N485 = ~signA_S;
  assign N31 = ~sExpB_S[10];
  assign N32 = ~sExpB_S[9];
  assign N33 = ~sExpB_S[8];
  assign N34 = ~sExpB_S[7];
  assign N35 = ~sExpB_S[6];
  assign N36 = ~sExpB_S[5];
  assign N37 = ~sExpB_S[4];
  assign N38 = ~sExpB_S[3];
  assign N39 = ~sExpB_S[2];
  assign N40 = ~sExpB_S[1];
  assign N41 = ~sExpB_S[0];
  assign N43 = ~N42;
  assign evenSqrt_S = sqrtOp & N486;
  assign N486 = ~sExpA_S[0];
  assign oddSqrt_S = sqrtOp & sExpA_S[0];
  assign entering = inReady & inValid;
  assign entering_normalCase = entering & normalCase_S;
  assign skipCycle2 = N462 & out_sig[55];
  assign step1Case = skipCycle2 | N44;
  assign N45 = ~nReset;
  assign N46 = inValid | N467;
  assign N47 = N74;
  assign N48 = entering & N487;
  assign N487 = ~normalCase_S;
  assign N49 = ~entering_normalCase;
  assign N55 = ~step1Case;
  assign N68 = entering_normalCase | N67;
  assign N69 = entering_normalCase | N66;
  assign N70 = entering_normalCase | N64;
  assign N71 = N54 | N63;
  assign N72 = N488 | N62;
  assign N488 = N48 | N53;
  assign N74 = N46 & nReset;
  assign N75 = nReset;
  assign N76 = N75 & entering_normalCase;
  assign N103 = entering_normalCase & N24;
  assign N104 = ~inReady;
  assign N105 = ~oddSqrt_S;
  assign trialTermSel[4] = inReady & N24;
  assign trialTermSel[3] = inReady & evenSqrt_S;
  assign trialTermSel[2] = inReady & oddSqrt_S;
  assign sigX_NSel[0] = ~inReady;
  assign trialTermSel[1] = sigX_NSel[0] & N489;
  assign N489 = ~sqrtOpOut;
  assign trialTermSel[0] = sigX_NSel[0] & sqrtOpOut;
  assign trialTermMuxIn_0__53_ = out_sig[53] | bitMask[53];
  assign trialTermMuxIn_0__52_ = out_sig[52] | bitMask[52];
  assign trialTermMuxIn_0__51_ = out_sig[51] | bitMask[51];
  assign trialTermMuxIn_0__50_ = out_sig[50] | bitMask[50];
  assign trialTermMuxIn_0__49_ = out_sig[49] | bitMask[49];
  assign trialTermMuxIn_0__48_ = out_sig[48] | bitMask[48];
  assign trialTermMuxIn_0__47_ = out_sig[47] | bitMask[47];
  assign trialTermMuxIn_0__46_ = out_sig[46] | bitMask[46];
  assign trialTermMuxIn_0__45_ = out_sig[45] | bitMask[45];
  assign trialTermMuxIn_0__44_ = out_sig[44] | bitMask[44];
  assign trialTermMuxIn_0__43_ = out_sig[43] | bitMask[43];
  assign trialTermMuxIn_0__42_ = out_sig[42] | bitMask[42];
  assign trialTermMuxIn_0__41_ = out_sig[41] | bitMask[41];
  assign trialTermMuxIn_0__40_ = out_sig[40] | bitMask[40];
  assign trialTermMuxIn_0__39_ = out_sig[39] | bitMask[39];
  assign trialTermMuxIn_0__38_ = out_sig[38] | bitMask[38];
  assign trialTermMuxIn_0__37_ = out_sig[37] | bitMask[37];
  assign trialTermMuxIn_0__36_ = out_sig[36] | bitMask[36];
  assign trialTermMuxIn_0__35_ = out_sig[35] | bitMask[35];
  assign trialTermMuxIn_0__34_ = out_sig[34] | bitMask[34];
  assign trialTermMuxIn_0__33_ = out_sig[33] | bitMask[33];
  assign trialTermMuxIn_0__32_ = out_sig[32] | bitMask[32];
  assign trialTermMuxIn_0__31_ = out_sig[31] | bitMask[31];
  assign trialTermMuxIn_0__30_ = out_sig[30] | bitMask[30];
  assign trialTermMuxIn_0__29_ = out_sig[29] | bitMask[29];
  assign trialTermMuxIn_0__28_ = out_sig[28] | bitMask[28];
  assign trialTermMuxIn_0__27_ = out_sig[27] | bitMask[27];
  assign trialTermMuxIn_0__26_ = out_sig[26] | bitMask[26];
  assign trialTermMuxIn_0__25_ = out_sig[25] | bitMask[25];
  assign trialTermMuxIn_0__24_ = out_sig[24] | bitMask[24];
  assign trialTermMuxIn_0__23_ = out_sig[23] | bitMask[23];
  assign trialTermMuxIn_0__22_ = out_sig[22] | bitMask[22];
  assign trialTermMuxIn_0__21_ = out_sig[21] | bitMask[21];
  assign trialTermMuxIn_0__20_ = out_sig[20] | bitMask[20];
  assign trialTermMuxIn_0__19_ = out_sig[19] | bitMask[19];
  assign trialTermMuxIn_0__18_ = out_sig[18] | bitMask[18];
  assign trialTermMuxIn_0__17_ = out_sig[17] | bitMask[17];
  assign trialTermMuxIn_0__16_ = out_sig[16] | bitMask[16];
  assign trialTermMuxIn_0__15_ = out_sig[15] | bitMask[15];
  assign trialTermMuxIn_0__14_ = out_sig[14] | bitMask[14];
  assign trialTermMuxIn_0__13_ = out_sig[13] | bitMask[13];
  assign trialTermMuxIn_0__12_ = out_sig[12] | bitMask[12];
  assign trialTermMuxIn_0__11_ = out_sig[11] | bitMask[11];
  assign trialTermMuxIn_0__10_ = out_sig[10] | bitMask[10];
  assign trialTermMuxIn_0__9_ = out_sig[9] | bitMask[9];
  assign trialTermMuxIn_0__8_ = out_sig[8] | bitMask[8];
  assign trialTermMuxIn_0__7_ = out_sig[7] | bitMask[7];
  assign trialTermMuxIn_0__6_ = out_sig[6] | bitMask[6];
  assign trialTermMuxIn_0__5_ = out_sig[5] | bitMask[5];
  assign trialTermMuxIn_0__4_ = out_sig[4] | bitMask[4];
  assign trialTermMuxIn_0__3_ = out_sig[3] | bitMask[3];
  assign trialTermMuxIn_0__2_ = out_sig[2] | bitMask[2];
  assign trialTermMuxIn_0__1_ = out_sig[1] | bitMask[1];
  assign N161 = ~sigX_NMuxIn_3__54_;
  assign N162 = sigX_NMuxIn_3__54_;
  assign sigXNext[53] = out_sig[54] | N216;
  assign sigXNext[52] = out_sig[53] | N215;
  assign sigXNext[51] = out_sig[52] | N214;
  assign sigXNext[50] = out_sig[51] | N213;
  assign sigXNext[49] = out_sig[50] | N212;
  assign sigXNext[48] = out_sig[49] | N211;
  assign sigXNext[47] = out_sig[48] | N210;
  assign sigXNext[46] = out_sig[47] | N209;
  assign sigXNext[45] = out_sig[46] | N208;
  assign sigXNext[44] = out_sig[45] | N207;
  assign sigXNext[43] = out_sig[44] | N206;
  assign sigXNext[42] = out_sig[43] | N205;
  assign sigXNext[41] = out_sig[42] | N204;
  assign sigXNext[40] = out_sig[41] | N203;
  assign sigXNext[39] = out_sig[40] | N202;
  assign sigXNext[38] = out_sig[39] | N201;
  assign sigXNext[37] = out_sig[38] | N200;
  assign sigXNext[36] = out_sig[37] | N199;
  assign sigXNext[35] = out_sig[36] | N198;
  assign sigXNext[34] = out_sig[35] | N197;
  assign sigXNext[33] = out_sig[34] | N196;
  assign sigXNext[32] = out_sig[33] | N195;
  assign sigXNext[31] = out_sig[32] | N194;
  assign sigXNext[30] = out_sig[31] | N193;
  assign sigXNext[29] = out_sig[30] | N192;
  assign sigXNext[28] = out_sig[29] | N191;
  assign sigXNext[27] = out_sig[28] | N190;
  assign sigXNext[26] = out_sig[27] | N189;
  assign sigXNext[25] = out_sig[26] | N188;
  assign sigXNext[24] = out_sig[25] | N187;
  assign sigXNext[23] = out_sig[24] | N186;
  assign sigXNext[22] = out_sig[23] | N185;
  assign sigXNext[21] = out_sig[22] | N184;
  assign sigXNext[20] = out_sig[21] | N183;
  assign sigXNext[19] = out_sig[20] | N182;
  assign sigXNext[18] = out_sig[19] | N181;
  assign sigXNext[17] = out_sig[18] | N180;
  assign sigXNext[16] = out_sig[17] | N179;
  assign sigXNext[15] = out_sig[16] | N178;
  assign sigXNext[14] = out_sig[15] | N177;
  assign sigXNext[13] = out_sig[14] | N176;
  assign sigXNext[12] = out_sig[13] | N175;
  assign sigXNext[11] = out_sig[12] | N174;
  assign sigXNext[10] = out_sig[11] | N173;
  assign sigXNext[9] = out_sig[10] | N172;
  assign sigXNext[8] = out_sig[9] | N171;
  assign sigXNext[7] = out_sig[8] | N170;
  assign sigXNext[6] = out_sig[7] | N169;
  assign sigXNext[5] = out_sig[6] | N168;
  assign sigXNext[4] = out_sig[5] | N167;
  assign sigXNext[3] = out_sig[4] | N166;
  assign sigXNext[2] = out_sig[3] | N165;
  assign sigXNext[1] = out_sig[2] | N164;
  assign sigXNext[0] = out_sig[1] | N163;
  assign N217 = sigXNext[52] | 1'b0;
  assign N218 = sigXNext[51] | bitMask[53];
  assign N219 = sigXNext[50] | bitMask[52];
  assign N220 = sigXNext[49] | bitMask[51];
  assign N221 = sigXNext[48] | bitMask[50];
  assign N222 = sigXNext[47] | bitMask[49];
  assign N223 = sigXNext[46] | bitMask[48];
  assign N224 = sigXNext[45] | bitMask[47];
  assign N225 = sigXNext[44] | bitMask[46];
  assign N226 = sigXNext[43] | bitMask[45];
  assign N227 = sigXNext[42] | bitMask[44];
  assign N228 = sigXNext[41] | bitMask[43];
  assign N229 = sigXNext[40] | bitMask[42];
  assign N230 = sigXNext[39] | bitMask[41];
  assign N231 = sigXNext[38] | bitMask[40];
  assign N232 = sigXNext[37] | bitMask[39];
  assign N233 = sigXNext[36] | bitMask[38];
  assign N234 = sigXNext[35] | bitMask[37];
  assign N235 = sigXNext[34] | bitMask[36];
  assign N236 = sigXNext[33] | bitMask[35];
  assign N237 = sigXNext[32] | bitMask[34];
  assign N238 = sigXNext[31] | bitMask[33];
  assign N239 = sigXNext[30] | bitMask[32];
  assign N240 = sigXNext[29] | bitMask[31];
  assign N241 = sigXNext[28] | bitMask[30];
  assign N242 = sigXNext[27] | bitMask[29];
  assign N243 = sigXNext[26] | bitMask[28];
  assign N244 = sigXNext[25] | bitMask[27];
  assign N245 = sigXNext[24] | bitMask[26];
  assign N246 = sigXNext[23] | bitMask[25];
  assign N247 = sigXNext[22] | bitMask[24];
  assign N248 = sigXNext[21] | bitMask[23];
  assign N249 = sigXNext[20] | bitMask[22];
  assign N250 = sigXNext[19] | bitMask[21];
  assign N251 = sigXNext[18] | bitMask[20];
  assign N252 = sigXNext[17] | bitMask[19];
  assign N253 = sigXNext[16] | bitMask[18];
  assign N254 = sigXNext[15] | bitMask[17];
  assign N255 = sigXNext[14] | bitMask[16];
  assign N256 = sigXNext[13] | bitMask[15];
  assign N257 = sigXNext[12] | bitMask[14];
  assign N258 = sigXNext[11] | bitMask[13];
  assign N259 = sigXNext[10] | bitMask[12];
  assign N260 = sigXNext[9] | bitMask[11];
  assign N261 = sigXNext[8] | bitMask[10];
  assign N262 = sigXNext[7] | bitMask[9];
  assign N263 = sigXNext[6] | bitMask[8];
  assign N264 = sigXNext[5] | bitMask[7];
  assign N265 = sigXNext[4] | bitMask[6];
  assign N266 = sigXNext[3] | bitMask[5];
  assign N267 = sigXNext[2] | bitMask[4];
  assign N268 = sigXNext[1] | bitMask[3];
  assign N269 = sigXNext[0] | bitMask[2];
  assign N270 = ~sigX_NMuxIn_3__54_;
  assign N271 = sigX_NMuxIn_3__54_;
  assign N272 = ~newBit2;
  assign sigX_NMuxIn_0__53_ = sigXNext[53] | 1'b0;
  assign sigX_NMuxIn_0__52_ = sigXNext[52] | N325;
  assign sigX_NMuxIn_0__51_ = sigXNext[51] | N324;
  assign sigX_NMuxIn_0__50_ = sigXNext[50] | N323;
  assign sigX_NMuxIn_0__49_ = sigXNext[49] | N322;
  assign sigX_NMuxIn_0__48_ = sigXNext[48] | N321;
  assign sigX_NMuxIn_0__47_ = sigXNext[47] | N320;
  assign sigX_NMuxIn_0__46_ = sigXNext[46] | N319;
  assign sigX_NMuxIn_0__45_ = sigXNext[45] | N318;
  assign sigX_NMuxIn_0__44_ = sigXNext[44] | N317;
  assign sigX_NMuxIn_0__43_ = sigXNext[43] | N316;
  assign sigX_NMuxIn_0__42_ = sigXNext[42] | N315;
  assign sigX_NMuxIn_0__41_ = sigXNext[41] | N314;
  assign sigX_NMuxIn_0__40_ = sigXNext[40] | N313;
  assign sigX_NMuxIn_0__39_ = sigXNext[39] | N312;
  assign sigX_NMuxIn_0__38_ = sigXNext[38] | N311;
  assign sigX_NMuxIn_0__37_ = sigXNext[37] | N310;
  assign sigX_NMuxIn_0__36_ = sigXNext[36] | N309;
  assign sigX_NMuxIn_0__35_ = sigXNext[35] | N308;
  assign sigX_NMuxIn_0__34_ = sigXNext[34] | N307;
  assign sigX_NMuxIn_0__33_ = sigXNext[33] | N306;
  assign sigX_NMuxIn_0__32_ = sigXNext[32] | N305;
  assign sigX_NMuxIn_0__31_ = sigXNext[31] | N304;
  assign sigX_NMuxIn_0__30_ = sigXNext[30] | N303;
  assign sigX_NMuxIn_0__29_ = sigXNext[29] | N302;
  assign sigX_NMuxIn_0__28_ = sigXNext[28] | N301;
  assign sigX_NMuxIn_0__27_ = sigXNext[27] | N300;
  assign sigX_NMuxIn_0__26_ = sigXNext[26] | N299;
  assign sigX_NMuxIn_0__25_ = sigXNext[25] | N298;
  assign sigX_NMuxIn_0__24_ = sigXNext[24] | N297;
  assign sigX_NMuxIn_0__23_ = sigXNext[23] | N296;
  assign sigX_NMuxIn_0__22_ = sigXNext[22] | N295;
  assign sigX_NMuxIn_0__21_ = sigXNext[21] | N294;
  assign sigX_NMuxIn_0__20_ = sigXNext[20] | N293;
  assign sigX_NMuxIn_0__19_ = sigXNext[19] | N292;
  assign sigX_NMuxIn_0__18_ = sigXNext[18] | N291;
  assign sigX_NMuxIn_0__17_ = sigXNext[17] | N290;
  assign sigX_NMuxIn_0__16_ = sigXNext[16] | N289;
  assign sigX_NMuxIn_0__15_ = sigXNext[15] | N288;
  assign sigX_NMuxIn_0__14_ = sigXNext[14] | N287;
  assign sigX_NMuxIn_0__13_ = sigXNext[13] | N286;
  assign sigX_NMuxIn_0__12_ = sigXNext[12] | N285;
  assign sigX_NMuxIn_0__11_ = sigXNext[11] | N284;
  assign sigX_NMuxIn_0__10_ = sigXNext[10] | N283;
  assign sigX_NMuxIn_0__9_ = sigXNext[9] | N282;
  assign sigX_NMuxIn_0__8_ = sigXNext[8] | N281;
  assign sigX_NMuxIn_0__7_ = sigXNext[7] | N280;
  assign sigX_NMuxIn_0__6_ = sigXNext[6] | N279;
  assign sigX_NMuxIn_0__5_ = sigXNext[5] | N278;
  assign sigX_NMuxIn_0__4_ = sigXNext[4] | N277;
  assign sigX_NMuxIn_0__3_ = sigXNext[3] | N276;
  assign sigX_NMuxIn_0__2_ = sigXNext[2] | N275;
  assign sigX_NMuxIn_0__1_ = sigXNext[1] | N274;
  assign sigX_NMuxIn_0__0_ = sigXNext[0] | N273;
  assign N327 = entering_normalCase | N326;
  assign N328 = inReady | skipCycle2;
  assign N329 = newBit2 | N328;
  assign N330 = ~N329;
  assign N331 = ~sigX_NMuxIn_3__54_;
  assign N332 = sigX_NMuxIn_3__54_;
  assign N443 = entering_normalCase | N491;
  assign N491 = N104 & N490;
  assign N490 = sigX_NMuxIn_3__54_ | newBit2;
  assign N446 = N444 & N445;
  assign N447 = ~N328;
  assign N448 = newBit2 & N447;
  assign invalidExc = majorExc_Z & out_isNaN;
  assign infiniteExc = majorExc_Z & N492;
  assign N492 = ~out_isNaN;
  assign N2 = ~N46;

  always @(posedge clock) begin
    if(N45) begin
      cycleNum_5_sv2v_reg <= 1'b0;
      cycleNum_4_sv2v_reg <= 1'b0;
      cycleNum_3_sv2v_reg <= 1'b0;
      cycleNum_2_sv2v_reg <= 1'b0;
      cycleNum_1_sv2v_reg <= 1'b0;
      cycleNum_0_sv2v_reg <= 1'b0;
    end else if(N73) begin
      cycleNum_5_sv2v_reg <= N68;
      cycleNum_4_sv2v_reg <= N69;
      cycleNum_3_sv2v_reg <= N65;
      cycleNum_2_sv2v_reg <= N70;
      cycleNum_1_sv2v_reg <= N71;
      cycleNum_0_sv2v_reg <= N72;
    end 
    if(N45) begin
      fractB_Z_51_sv2v_reg <= 1'b0;
      fractB_Z_50_sv2v_reg <= 1'b0;
      fractB_Z_49_sv2v_reg <= 1'b0;
      fractB_Z_48_sv2v_reg <= 1'b0;
      fractB_Z_47_sv2v_reg <= 1'b0;
      fractB_Z_46_sv2v_reg <= 1'b0;
      fractB_Z_45_sv2v_reg <= 1'b0;
      fractB_Z_44_sv2v_reg <= 1'b0;
      fractB_Z_43_sv2v_reg <= 1'b0;
      fractB_Z_42_sv2v_reg <= 1'b0;
      fractB_Z_41_sv2v_reg <= 1'b0;
      fractB_Z_40_sv2v_reg <= 1'b0;
      fractB_Z_39_sv2v_reg <= 1'b0;
      fractB_Z_38_sv2v_reg <= 1'b0;
      fractB_Z_37_sv2v_reg <= 1'b0;
      fractB_Z_36_sv2v_reg <= 1'b0;
      fractB_Z_35_sv2v_reg <= 1'b0;
      fractB_Z_34_sv2v_reg <= 1'b0;
      fractB_Z_33_sv2v_reg <= 1'b0;
      fractB_Z_32_sv2v_reg <= 1'b0;
      fractB_Z_31_sv2v_reg <= 1'b0;
      fractB_Z_30_sv2v_reg <= 1'b0;
      fractB_Z_29_sv2v_reg <= 1'b0;
      fractB_Z_28_sv2v_reg <= 1'b0;
      fractB_Z_27_sv2v_reg <= 1'b0;
      fractB_Z_26_sv2v_reg <= 1'b0;
      fractB_Z_25_sv2v_reg <= 1'b0;
      fractB_Z_24_sv2v_reg <= 1'b0;
      fractB_Z_23_sv2v_reg <= 1'b0;
      fractB_Z_22_sv2v_reg <= 1'b0;
      fractB_Z_21_sv2v_reg <= 1'b0;
      fractB_Z_20_sv2v_reg <= 1'b0;
      fractB_Z_19_sv2v_reg <= 1'b0;
      fractB_Z_18_sv2v_reg <= 1'b0;
      fractB_Z_17_sv2v_reg <= 1'b0;
      fractB_Z_16_sv2v_reg <= 1'b0;
      fractB_Z_15_sv2v_reg <= 1'b0;
      fractB_Z_14_sv2v_reg <= 1'b0;
      fractB_Z_13_sv2v_reg <= 1'b0;
      fractB_Z_12_sv2v_reg <= 1'b0;
      fractB_Z_11_sv2v_reg <= 1'b0;
      fractB_Z_10_sv2v_reg <= 1'b0;
      fractB_Z_9_sv2v_reg <= 1'b0;
      fractB_Z_8_sv2v_reg <= 1'b0;
      fractB_Z_7_sv2v_reg <= 1'b0;
      fractB_Z_6_sv2v_reg <= 1'b0;
      fractB_Z_5_sv2v_reg <= 1'b0;
      fractB_Z_4_sv2v_reg <= 1'b0;
      fractB_Z_3_sv2v_reg <= 1'b0;
      fractB_Z_2_sv2v_reg <= 1'b0;
      fractB_Z_1_sv2v_reg <= 1'b0;
      fractB_Z_0_sv2v_reg <= 1'b0;
    end else if(N103) begin
      fractB_Z_51_sv2v_reg <= sigB_S[51];
      fractB_Z_50_sv2v_reg <= sigB_S[50];
      fractB_Z_49_sv2v_reg <= sigB_S[49];
      fractB_Z_48_sv2v_reg <= sigB_S[48];
      fractB_Z_47_sv2v_reg <= sigB_S[47];
      fractB_Z_46_sv2v_reg <= sigB_S[46];
      fractB_Z_45_sv2v_reg <= sigB_S[45];
      fractB_Z_44_sv2v_reg <= sigB_S[44];
      fractB_Z_43_sv2v_reg <= sigB_S[43];
      fractB_Z_42_sv2v_reg <= sigB_S[42];
      fractB_Z_41_sv2v_reg <= sigB_S[41];
      fractB_Z_40_sv2v_reg <= sigB_S[40];
      fractB_Z_39_sv2v_reg <= sigB_S[39];
      fractB_Z_38_sv2v_reg <= sigB_S[38];
      fractB_Z_37_sv2v_reg <= sigB_S[37];
      fractB_Z_36_sv2v_reg <= sigB_S[36];
      fractB_Z_35_sv2v_reg <= sigB_S[35];
      fractB_Z_34_sv2v_reg <= sigB_S[34];
      fractB_Z_33_sv2v_reg <= sigB_S[33];
      fractB_Z_32_sv2v_reg <= sigB_S[32];
      fractB_Z_31_sv2v_reg <= sigB_S[31];
      fractB_Z_30_sv2v_reg <= sigB_S[30];
      fractB_Z_29_sv2v_reg <= sigB_S[29];
      fractB_Z_28_sv2v_reg <= sigB_S[28];
      fractB_Z_27_sv2v_reg <= sigB_S[27];
      fractB_Z_26_sv2v_reg <= sigB_S[26];
      fractB_Z_25_sv2v_reg <= sigB_S[25];
      fractB_Z_24_sv2v_reg <= sigB_S[24];
      fractB_Z_23_sv2v_reg <= sigB_S[23];
      fractB_Z_22_sv2v_reg <= sigB_S[22];
      fractB_Z_21_sv2v_reg <= sigB_S[21];
      fractB_Z_20_sv2v_reg <= sigB_S[20];
      fractB_Z_19_sv2v_reg <= sigB_S[19];
      fractB_Z_18_sv2v_reg <= sigB_S[18];
      fractB_Z_17_sv2v_reg <= sigB_S[17];
      fractB_Z_16_sv2v_reg <= sigB_S[16];
      fractB_Z_15_sv2v_reg <= sigB_S[15];
      fractB_Z_14_sv2v_reg <= sigB_S[14];
      fractB_Z_13_sv2v_reg <= sigB_S[13];
      fractB_Z_12_sv2v_reg <= sigB_S[12];
      fractB_Z_11_sv2v_reg <= sigB_S[11];
      fractB_Z_10_sv2v_reg <= sigB_S[10];
      fractB_Z_9_sv2v_reg <= sigB_S[9];
      fractB_Z_8_sv2v_reg <= sigB_S[8];
      fractB_Z_7_sv2v_reg <= sigB_S[7];
      fractB_Z_6_sv2v_reg <= sigB_S[6];
      fractB_Z_5_sv2v_reg <= sigB_S[5];
      fractB_Z_4_sv2v_reg <= sigB_S[4];
      fractB_Z_3_sv2v_reg <= sigB_S[3];
      fractB_Z_2_sv2v_reg <= sigB_S[2];
      fractB_Z_1_sv2v_reg <= sigB_S[1];
      fractB_Z_0_sv2v_reg <= sigB_S[0];
    end 
    if(N45) begin
      sqrtOpOut_sv2v_reg <= 1'b0;
      majorExc_Z_sv2v_reg <= 1'b0;
      out_isNaN_sv2v_reg <= 1'b0;
      out_isInf_sv2v_reg <= 1'b0;
      out_isZero_sv2v_reg <= 1'b0;
      out_sign_sv2v_reg <= 1'b0;
    end else if(entering) begin
      sqrtOpOut_sv2v_reg <= sqrtOp;
      majorExc_Z_sv2v_reg <= majorExc_S;
      out_isNaN_sv2v_reg <= isNaN_S;
      out_isInf_sv2v_reg <= isInf_S;
      out_isZero_sv2v_reg <= isZero_S;
      out_sign_sv2v_reg <= sign_S;
    end 
    if(N45) begin
      out_sExp_12_sv2v_reg <= 1'b0;
      out_sExp_11_sv2v_reg <= 1'b0;
      out_sExp_10_sv2v_reg <= 1'b0;
      out_sExp_9_sv2v_reg <= 1'b0;
      out_sExp_8_sv2v_reg <= 1'b0;
      out_sExp_7_sv2v_reg <= 1'b0;
      out_sExp_6_sv2v_reg <= 1'b0;
      out_sExp_5_sv2v_reg <= 1'b0;
      out_sExp_4_sv2v_reg <= 1'b0;
      out_sExp_3_sv2v_reg <= 1'b0;
      out_sExp_2_sv2v_reg <= 1'b0;
      out_sExp_1_sv2v_reg <= 1'b0;
      out_sExp_0_sv2v_reg <= 1'b0;
      roundingModeOut_2_sv2v_reg <= 1'b0;
      roundingModeOut_1_sv2v_reg <= 1'b0;
      roundingModeOut_0_sv2v_reg <= 1'b0;
    end else if(entering_normalCase) begin
      out_sExp_12_sv2v_reg <= N102;
      out_sExp_11_sv2v_reg <= N101;
      out_sExp_10_sv2v_reg <= N100;
      out_sExp_9_sv2v_reg <= N99;
      out_sExp_8_sv2v_reg <= N98;
      out_sExp_7_sv2v_reg <= N97;
      out_sExp_6_sv2v_reg <= N96;
      out_sExp_5_sv2v_reg <= N95;
      out_sExp_4_sv2v_reg <= N94;
      out_sExp_3_sv2v_reg <= N93;
      out_sExp_2_sv2v_reg <= N92;
      out_sExp_1_sv2v_reg <= N91;
      out_sExp_0_sv2v_reg <= N90;
      roundingModeOut_2_sv2v_reg <= roundingMode[2];
      roundingModeOut_1_sv2v_reg <= roundingMode[1];
      roundingModeOut_0_sv2v_reg <= roundingMode[0];
    end 
    if(N45) begin
      out_sig_0_sv2v_reg <= 1'b0;
      out_sig_55_sv2v_reg <= 1'b0;
      out_sig_54_sv2v_reg <= 1'b0;
      out_sig_53_sv2v_reg <= 1'b0;
      out_sig_52_sv2v_reg <= 1'b0;
      out_sig_51_sv2v_reg <= 1'b0;
      out_sig_50_sv2v_reg <= 1'b0;
      out_sig_49_sv2v_reg <= 1'b0;
      out_sig_48_sv2v_reg <= 1'b0;
      out_sig_47_sv2v_reg <= 1'b0;
      out_sig_46_sv2v_reg <= 1'b0;
      out_sig_45_sv2v_reg <= 1'b0;
      out_sig_44_sv2v_reg <= 1'b0;
      out_sig_43_sv2v_reg <= 1'b0;
      out_sig_42_sv2v_reg <= 1'b0;
      out_sig_41_sv2v_reg <= 1'b0;
      out_sig_40_sv2v_reg <= 1'b0;
      out_sig_39_sv2v_reg <= 1'b0;
      out_sig_38_sv2v_reg <= 1'b0;
      out_sig_37_sv2v_reg <= 1'b0;
      out_sig_36_sv2v_reg <= 1'b0;
      out_sig_35_sv2v_reg <= 1'b0;
      out_sig_34_sv2v_reg <= 1'b0;
      out_sig_33_sv2v_reg <= 1'b0;
      out_sig_32_sv2v_reg <= 1'b0;
      out_sig_31_sv2v_reg <= 1'b0;
      out_sig_30_sv2v_reg <= 1'b0;
      out_sig_29_sv2v_reg <= 1'b0;
      out_sig_28_sv2v_reg <= 1'b0;
      out_sig_27_sv2v_reg <= 1'b0;
      out_sig_26_sv2v_reg <= 1'b0;
      out_sig_25_sv2v_reg <= 1'b0;
      out_sig_24_sv2v_reg <= 1'b0;
      out_sig_23_sv2v_reg <= 1'b0;
      out_sig_22_sv2v_reg <= 1'b0;
      out_sig_21_sv2v_reg <= 1'b0;
      out_sig_20_sv2v_reg <= 1'b0;
      out_sig_19_sv2v_reg <= 1'b0;
      out_sig_18_sv2v_reg <= 1'b0;
      out_sig_17_sv2v_reg <= 1'b0;
      out_sig_16_sv2v_reg <= 1'b0;
      out_sig_15_sv2v_reg <= 1'b0;
      out_sig_14_sv2v_reg <= 1'b0;
      out_sig_13_sv2v_reg <= 1'b0;
      out_sig_12_sv2v_reg <= 1'b0;
      out_sig_11_sv2v_reg <= 1'b0;
      out_sig_10_sv2v_reg <= 1'b0;
      out_sig_9_sv2v_reg <= 1'b0;
      out_sig_8_sv2v_reg <= 1'b0;
      out_sig_7_sv2v_reg <= 1'b0;
      out_sig_6_sv2v_reg <= 1'b0;
      out_sig_5_sv2v_reg <= 1'b0;
      out_sig_4_sv2v_reg <= 1'b0;
      out_sig_3_sv2v_reg <= 1'b0;
      out_sig_2_sv2v_reg <= 1'b0;
      out_sig_1_sv2v_reg <= 1'b0;
    end else if(N443) begin
      out_sig_0_sv2v_reg <= N446;
      out_sig_55_sv2v_reg <= sigX_N[54];
      out_sig_54_sv2v_reg <= sigX_N[53];
      out_sig_53_sv2v_reg <= sigX_N[52];
      out_sig_52_sv2v_reg <= sigX_N[51];
      out_sig_51_sv2v_reg <= sigX_N[50];
      out_sig_50_sv2v_reg <= sigX_N[49];
      out_sig_49_sv2v_reg <= sigX_N[48];
      out_sig_48_sv2v_reg <= sigX_N[47];
      out_sig_47_sv2v_reg <= sigX_N[46];
      out_sig_46_sv2v_reg <= sigX_N[45];
      out_sig_45_sv2v_reg <= sigX_N[44];
      out_sig_44_sv2v_reg <= sigX_N[43];
      out_sig_43_sv2v_reg <= sigX_N[42];
      out_sig_42_sv2v_reg <= sigX_N[41];
      out_sig_41_sv2v_reg <= sigX_N[40];
      out_sig_40_sv2v_reg <= sigX_N[39];
      out_sig_39_sv2v_reg <= sigX_N[38];
      out_sig_38_sv2v_reg <= sigX_N[37];
      out_sig_37_sv2v_reg <= sigX_N[36];
      out_sig_36_sv2v_reg <= sigX_N[35];
      out_sig_35_sv2v_reg <= sigX_N[34];
      out_sig_34_sv2v_reg <= sigX_N[33];
      out_sig_33_sv2v_reg <= sigX_N[32];
      out_sig_32_sv2v_reg <= sigX_N[31];
      out_sig_31_sv2v_reg <= sigX_N[30];
      out_sig_30_sv2v_reg <= sigX_N[29];
      out_sig_29_sv2v_reg <= sigX_N[28];
      out_sig_28_sv2v_reg <= sigX_N[27];
      out_sig_27_sv2v_reg <= sigX_N[26];
      out_sig_26_sv2v_reg <= sigX_N[25];
      out_sig_25_sv2v_reg <= sigX_N[24];
      out_sig_24_sv2v_reg <= sigX_N[23];
      out_sig_23_sv2v_reg <= sigX_N[22];
      out_sig_22_sv2v_reg <= sigX_N[21];
      out_sig_21_sv2v_reg <= sigX_N[20];
      out_sig_20_sv2v_reg <= sigX_N[19];
      out_sig_19_sv2v_reg <= sigX_N[18];
      out_sig_18_sv2v_reg <= sigX_N[17];
      out_sig_17_sv2v_reg <= sigX_N[16];
      out_sig_16_sv2v_reg <= sigX_N[15];
      out_sig_15_sv2v_reg <= sigX_N[14];
      out_sig_14_sv2v_reg <= sigX_N[13];
      out_sig_13_sv2v_reg <= sigX_N[12];
      out_sig_12_sv2v_reg <= sigX_N[11];
      out_sig_11_sv2v_reg <= sigX_N[10];
      out_sig_10_sv2v_reg <= sigX_N[9];
      out_sig_9_sv2v_reg <= sigX_N[8];
      out_sig_8_sv2v_reg <= sigX_N[7];
      out_sig_7_sv2v_reg <= sigX_N[6];
      out_sig_6_sv2v_reg <= sigX_N[5];
      out_sig_5_sv2v_reg <= sigX_N[4];
      out_sig_4_sv2v_reg <= sigX_N[3];
      out_sig_3_sv2v_reg <= sigX_N[2];
      out_sig_2_sv2v_reg <= sigX_N[1];
      out_sig_1_sv2v_reg <= sigX_N[0];
    end 
    if(N45) begin
      rem_Z_54_sv2v_reg <= 1'b0;
      rem_Z_53_sv2v_reg <= 1'b0;
      rem_Z_52_sv2v_reg <= 1'b0;
      rem_Z_51_sv2v_reg <= 1'b0;
      rem_Z_50_sv2v_reg <= 1'b0;
      rem_Z_49_sv2v_reg <= 1'b0;
      rem_Z_48_sv2v_reg <= 1'b0;
      rem_Z_47_sv2v_reg <= 1'b0;
      rem_Z_46_sv2v_reg <= 1'b0;
      rem_Z_45_sv2v_reg <= 1'b0;
      rem_Z_44_sv2v_reg <= 1'b0;
      rem_Z_43_sv2v_reg <= 1'b0;
      rem_Z_42_sv2v_reg <= 1'b0;
      rem_Z_41_sv2v_reg <= 1'b0;
      rem_Z_40_sv2v_reg <= 1'b0;
      rem_Z_39_sv2v_reg <= 1'b0;
      rem_Z_38_sv2v_reg <= 1'b0;
      rem_Z_37_sv2v_reg <= 1'b0;
      rem_Z_36_sv2v_reg <= 1'b0;
      rem_Z_35_sv2v_reg <= 1'b0;
      rem_Z_34_sv2v_reg <= 1'b0;
      rem_Z_33_sv2v_reg <= 1'b0;
      rem_Z_32_sv2v_reg <= 1'b0;
      rem_Z_31_sv2v_reg <= 1'b0;
      rem_Z_30_sv2v_reg <= 1'b0;
      rem_Z_29_sv2v_reg <= 1'b0;
      rem_Z_28_sv2v_reg <= 1'b0;
      rem_Z_27_sv2v_reg <= 1'b0;
      rem_Z_26_sv2v_reg <= 1'b0;
      rem_Z_25_sv2v_reg <= 1'b0;
      rem_Z_24_sv2v_reg <= 1'b0;
      rem_Z_23_sv2v_reg <= 1'b0;
      rem_Z_22_sv2v_reg <= 1'b0;
      rem_Z_21_sv2v_reg <= 1'b0;
      rem_Z_20_sv2v_reg <= 1'b0;
      rem_Z_19_sv2v_reg <= 1'b0;
      rem_Z_18_sv2v_reg <= 1'b0;
      rem_Z_17_sv2v_reg <= 1'b0;
      rem_Z_16_sv2v_reg <= 1'b0;
      rem_Z_15_sv2v_reg <= 1'b0;
      rem_Z_14_sv2v_reg <= 1'b0;
      rem_Z_13_sv2v_reg <= 1'b0;
      rem_Z_12_sv2v_reg <= 1'b0;
      rem_Z_11_sv2v_reg <= 1'b0;
      rem_Z_10_sv2v_reg <= 1'b0;
      rem_Z_9_sv2v_reg <= 1'b0;
      rem_Z_8_sv2v_reg <= 1'b0;
      rem_Z_7_sv2v_reg <= 1'b0;
      rem_Z_6_sv2v_reg <= 1'b0;
      rem_Z_5_sv2v_reg <= 1'b0;
      rem_Z_4_sv2v_reg <= 1'b0;
      rem_Z_3_sv2v_reg <= 1'b0;
      rem_Z_2_sv2v_reg <= 1'b0;
      rem_Z_1_sv2v_reg <= 1'b0;
      rem_Z_0_sv2v_reg <= 1'b0;
    end else if(N327) begin
      rem_Z_54_sv2v_reg <= N442;
      rem_Z_53_sv2v_reg <= N441;
      rem_Z_52_sv2v_reg <= N440;
      rem_Z_51_sv2v_reg <= N439;
      rem_Z_50_sv2v_reg <= N438;
      rem_Z_49_sv2v_reg <= N437;
      rem_Z_48_sv2v_reg <= N436;
      rem_Z_47_sv2v_reg <= N435;
      rem_Z_46_sv2v_reg <= N434;
      rem_Z_45_sv2v_reg <= N433;
      rem_Z_44_sv2v_reg <= N432;
      rem_Z_43_sv2v_reg <= N431;
      rem_Z_42_sv2v_reg <= N430;
      rem_Z_41_sv2v_reg <= N429;
      rem_Z_40_sv2v_reg <= N428;
      rem_Z_39_sv2v_reg <= N427;
      rem_Z_38_sv2v_reg <= N426;
      rem_Z_37_sv2v_reg <= N425;
      rem_Z_36_sv2v_reg <= N424;
      rem_Z_35_sv2v_reg <= N423;
      rem_Z_34_sv2v_reg <= N422;
      rem_Z_33_sv2v_reg <= N421;
      rem_Z_32_sv2v_reg <= N420;
      rem_Z_31_sv2v_reg <= N419;
      rem_Z_30_sv2v_reg <= N418;
      rem_Z_29_sv2v_reg <= N417;
      rem_Z_28_sv2v_reg <= N416;
      rem_Z_27_sv2v_reg <= N415;
      rem_Z_26_sv2v_reg <= N414;
      rem_Z_25_sv2v_reg <= N413;
      rem_Z_24_sv2v_reg <= N412;
      rem_Z_23_sv2v_reg <= N411;
      rem_Z_22_sv2v_reg <= N410;
      rem_Z_21_sv2v_reg <= N409;
      rem_Z_20_sv2v_reg <= N408;
      rem_Z_19_sv2v_reg <= N407;
      rem_Z_18_sv2v_reg <= N406;
      rem_Z_17_sv2v_reg <= N405;
      rem_Z_16_sv2v_reg <= N404;
      rem_Z_15_sv2v_reg <= N403;
      rem_Z_14_sv2v_reg <= N402;
      rem_Z_13_sv2v_reg <= N401;
      rem_Z_12_sv2v_reg <= N400;
      rem_Z_11_sv2v_reg <= N399;
      rem_Z_10_sv2v_reg <= N398;
      rem_Z_9_sv2v_reg <= N397;
      rem_Z_8_sv2v_reg <= N396;
      rem_Z_7_sv2v_reg <= N395;
      rem_Z_6_sv2v_reg <= N394;
      rem_Z_5_sv2v_reg <= N393;
      rem_Z_4_sv2v_reg <= N392;
      rem_Z_3_sv2v_reg <= N391;
      rem_Z_2_sv2v_reg <= N390;
      rem_Z_1_sv2v_reg <= N389;
      rem_Z_0_sv2v_reg <= N388;
    end 
  end


endmodule



module divSqrtRecFNToRaw_11_53_2
(
  nReset,
  clock,
  control,
  inReady,
  inValid,
  sqrtOp,
  a,
  b,
  roundingMode,
  outValid,
  sqrtOpOut,
  roundingModeOut,
  invalidExc,
  infiniteExc,
  out_isNaN,
  out_isInf,
  out_isZero,
  out_sign,
  out_sExp,
  out_sig
);

  input [0:0] control;
  input [64:0] a;
  input [64:0] b;
  input [2:0] roundingMode;
  output [2:0] roundingModeOut;
  output [12:0] out_sExp;
  output [55:0] out_sig;
  input nReset;
  input clock;
  input inValid;
  input sqrtOp;
  output inReady;
  output outValid;
  output sqrtOpOut;
  output invalidExc;
  output infiniteExc;
  output out_isNaN;
  output out_isInf;
  output out_isZero;
  output out_sign;
  wire [2:0] roundingModeOut;
  wire [12:0] out_sExp;
  wire [55:0] out_sig;
  wire inReady,outValid,sqrtOpOut,invalidExc,infiniteExc,out_isNaN,out_isInf,
  out_isZero,out_sign;

  divSqrtRecFNToRaw_medium_expWidth11_sigWidth53_options0
  \divSqrtTwoBitPerIter.divSqrtRecFNToRaw 
  (
    .nReset(nReset),
    .clock(clock),
    .control(control[0]),
    .inReady(inReady),
    .inValid(inValid),
    .sqrtOp(sqrtOp),
    .a(a),
    .b(b),
    .roundingMode(roundingMode),
    .outValid(outValid),
    .sqrtOpOut(sqrtOpOut),
    .roundingModeOut(roundingModeOut),
    .invalidExc(invalidExc),
    .infiniteExc(infiniteExc),
    .out_isNaN(out_isNaN),
    .out_isInf(out_isInf),
    .out_isZero(out_isZero),
    .out_sign(out_sign),
    .out_sExp(out_sExp),
    .out_sig(out_sig)
  );


endmodule



module bsg_dff_en_width_p9
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [8:0] data_i;
  output [8:0] data_o;
  input clk_i;
  input en_i;
  wire [8:0] data_o;
  reg data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,
  data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bp_be_pipe_long_00
(
  clk_i,
  reset_i,
  reservation_i,
  ibusy_o,
  fbusy_o,
  frm_dyn_i,
  flush_i,
  iwb_pkt_o,
  iwb_v_o,
  iwb_yumi_i,
  fwb_pkt_o,
  fwb_v_o,
  fwb_yumi_i
);

  input [520:0] reservation_i;
  input [2:0] frm_dyn_i;
  output [78:0] iwb_pkt_o;
  output [78:0] fwb_pkt_o;
  input clk_i;
  input reset_i;
  input flush_i;
  input iwb_yumi_i;
  input fwb_yumi_i;
  output ibusy_o;
  output fbusy_o;
  output iwb_v_o;
  output fwb_v_o;
  wire [78:0] iwb_pkt_o,fwb_pkt_o;
  wire ibusy_o,fbusy_o,iwb_v_o,fwb_v_o,N0,N1,N2,N3,N4,iwb_pkt_o_78_,fwb_pkt_o_77_,
  int_v_li,fp_v_li,fmask_r,imask_r,flush_int_li,flush_fp_li,N5,N6,N7,N8,N9,N10,N11,N12,
  N13,N14,N15,signed_div_li,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,
  N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,signed_opA_li,N42,N43,N44,N45,
  N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,signed_opB_li,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  imulh_v_li,_2_net_,imulh_ready_lo,imulh_v_lo,_4_net_,N82,N83,N84,N85,N86,N87,N88,
  N89,N90,N91,N92,N93,idiv_v_li,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,
  N105,N106,irem_v_li,_5_net_,_6_net_,idiv_ready_and_lo,idiv_v_lo,_7_net_,_8_net_,
  N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,
  N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,
  N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,
  N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,
  N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
  N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,
  fdiv_v_li,N203,N204,N205,fsqrt_v_li,fdivsqrt_v_li,_12_net_,fdivsqrt_ready_and_lo,
  fdivsqrt_v_lo,sqrt_lo,invalid_exc,infinite_exc,_19_net_,_20_net_,_21_net_,
  fdivsqrt_pending_r,fdivsqrt_pending,frd_tag_r,fflags_lo_nv_,fflags_lo_dz_,
  fflags_lo_of_,fflags_lo_uf_,fflags_lo_nx_,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,
  N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231;
  wire [63:0] imulh_result_lo,quotient_lo,remainder_lo,iresult;
  wire [5:0] fu_op_r;
  wire [1:0] ird_tag_r;
  wire [2:0] frm_li,frm_lo,frm_r;
  wire [74:0] fdivsqrt_raw_lo;
  assign fwb_pkt_o[76] = 1'b0;
  assign fwb_pkt_o[78] = 1'b0;
  assign iwb_pkt_o[0] = 1'b0;
  assign iwb_pkt_o[1] = 1'b0;
  assign iwb_pkt_o[2] = 1'b0;
  assign iwb_pkt_o[3] = 1'b0;
  assign iwb_pkt_o[4] = 1'b0;
  assign iwb_pkt_o[76] = 1'b0;
  assign iwb_pkt_o[77] = 1'b0;
  assign iwb_v_o = iwb_pkt_o_78_;
  assign iwb_pkt_o[78] = iwb_pkt_o_78_;
  assign fwb_v_o = fwb_pkt_o_77_;
  assign fwb_pkt_o[77] = fwb_pkt_o_77_;

  bsg_dff_width_p2
  mask_reg
  (
    .clk_i(clk_i),
    .data_i({ fp_v_li, int_v_li }),
    .data_o({ fmask_r, imask_r })
  );

  assign N5 = reservation_i[407] | N197;
  assign N6 = reservation_i[406] | N5;
  assign N7 = reservation_i[405] | N6;
  assign N8 = N203 | N7;
  assign N9 = ~N8;
  assign N10 = ~reservation_i[405];
  assign N11 = reservation_i[407] | N197;
  assign N12 = reservation_i[406] | N11;
  assign N13 = N10 | N12;
  assign N14 = N203 | N13;
  assign N15 = ~N14;
  assign signed_div_li = N9 | N15;
  assign N16 = reservation_i[407] | N197;
  assign N17 = reservation_i[406] | N16;
  assign N18 = reservation_i[405] | N17;
  assign N19 = N203 | N18;
  assign N20 = ~N19;
  assign N21 = ~reservation_i[405];
  assign N22 = reservation_i[407] | N197;
  assign N23 = reservation_i[406] | N22;
  assign N24 = N21 | N23;
  assign N25 = N203 | N24;
  assign N26 = ~N25;
  assign N27 = N20 | N26;
  assign N28 = ~reservation_i[406];
  assign N29 = reservation_i[407] | N197;
  assign N30 = N28 | N29;
  assign N31 = reservation_i[405] | N30;
  assign N32 = N203 | N31;
  assign N33 = ~N32;
  assign N34 = N27 | N33;
  assign N35 = ~reservation_i[406];
  assign N36 = ~reservation_i[405];
  assign N37 = reservation_i[407] | N197;
  assign N38 = N35 | N37;
  assign N39 = N36 | N38;
  assign N40 = reservation_i[404] | N39;
  assign N41 = ~N40;
  assign signed_opA_li = N34 | N41;
  assign N42 = reservation_i[407] | N197;
  assign N43 = reservation_i[406] | N42;
  assign N44 = reservation_i[405] | N43;
  assign N45 = N203 | N44;
  assign N46 = ~N45;
  assign N47 = ~reservation_i[405];
  assign N48 = reservation_i[407] | N197;
  assign N49 = reservation_i[406] | N48;
  assign N50 = N47 | N49;
  assign N51 = N203 | N50;
  assign N52 = ~N51;
  assign N53 = N46 | N52;
  assign N54 = ~reservation_i[406];
  assign N55 = reservation_i[407] | N197;
  assign N56 = N54 | N55;
  assign N57 = reservation_i[405] | N56;
  assign N58 = N203 | N57;
  assign N59 = ~N58;
  assign signed_opB_li = N53 | N59;
  assign N60 = ~reservation_i[406];
  assign N61 = reservation_i[407] | N197;
  assign N62 = N60 | N61;
  assign N63 = reservation_i[405] | N62;
  assign N64 = N203 | N63;
  assign N65 = ~N64;
  assign N66 = ~reservation_i[406];
  assign N67 = ~reservation_i[405];
  assign N68 = reservation_i[407] | N197;
  assign N69 = N66 | N68;
  assign N70 = N67 | N69;
  assign N71 = reservation_i[404] | N70;
  assign N72 = ~N71;
  assign N73 = N65 | N72;
  assign N74 = ~reservation_i[406];
  assign N75 = ~reservation_i[405];
  assign N76 = reservation_i[407] | N197;
  assign N77 = N74 | N76;
  assign N78 = N75 | N77;
  assign N79 = N203 | N78;
  assign N80 = ~N79;
  assign N81 = N73 | N80;

  bsg_imul_iterative_width_p64
  imulh
  (
    .clk_i(clk_i),
    .reset_i(_2_net_),
    .v_i(imulh_v_li),
    .ready_and_o(imulh_ready_lo),
    .opA_i(reservation_i[388:325]),
    .signed_opA_i(signed_opA_li),
    .opB_i(reservation_i[323:260]),
    .signed_opB_i(signed_opB_li),
    .gets_high_part_i(1'b1),
    .v_o(imulh_v_lo),
    .result_o(imulh_result_lo),
    .yumi_i(_4_net_)
  );

  assign N82 = reservation_i[407] | N197;
  assign N83 = reservation_i[406] | N82;
  assign N84 = reservation_i[405] | N83;
  assign N85 = N203 | N84;
  assign N86 = ~N85;
  assign N87 = ~reservation_i[405];
  assign N88 = reservation_i[407] | N197;
  assign N89 = reservation_i[406] | N88;
  assign N90 = N87 | N89;
  assign N91 = reservation_i[404] | N90;
  assign N92 = ~N91;
  assign N93 = N86 | N92;
  assign N94 = ~reservation_i[405];
  assign N95 = reservation_i[407] | N197;
  assign N96 = reservation_i[406] | N95;
  assign N97 = N94 | N96;
  assign N98 = N203 | N97;
  assign N99 = ~N98;
  assign N100 = ~reservation_i[406];
  assign N101 = reservation_i[407] | N197;
  assign N102 = N100 | N101;
  assign N103 = reservation_i[405] | N102;
  assign N104 = reservation_i[404] | N103;
  assign N105 = ~N104;
  assign N106 = N99 | N105;

  bsg_idiv_iterative_64_2
  idiv
  (
    .clk_i(clk_i),
    .reset_i(_5_net_),
    .v_i(_6_net_),
    .ready_and_o(idiv_ready_and_lo),
    .dividend_i(reservation_i[388:325]),
    .divisor_i(reservation_i[323:260]),
    .signed_div_i(signed_div_li),
    .v_o(idiv_v_lo),
    .quotient_o(quotient_lo),
    .remainder_o(remainder_lo),
    .yumi_i(_7_net_)
  );


  bsg_dff_en_width_p13
  iwb_reg
  (
    .clk_i(clk_i),
    .data_i({ reservation_i[460:456], reservation_i[409:404], reservation_i[402:401] }),
    .en_i(_8_net_),
    .data_o({ iwb_pkt_o[75:71], fu_op_r, ird_tag_r })
  );

  assign N110 = N107 & N108;
  assign N111 = N110 & N109;
  assign N115 = fu_op_r[2] | N113;
  assign N116 = N115 | N114;
  assign N118 = N117 | fu_op_r[1];
  assign N119 = N118 | fu_op_r[0];
  assign N121 = fu_op_r[2] | fu_op_r[1];
  assign N122 = N121 | N114;
  assign N123 = fu_op_r[2] | N113;
  assign N124 = N123 | fu_op_r[0];
  assign N126 = fu_op_r[2] & fu_op_r[0];
  assign N127 = fu_op_r[2] & fu_op_r[1];
  assign N128 = N117 & N113;
  assign N129 = N128 & N114;

  bp_be_int_box_00
  ird_box
  (
    .raw_i(iresult),
    .tag_i(ird_tag_r),
    .unsigned_i(1'b0),
    .reg_o(iwb_pkt_o[70:5])
  );

  assign N196 = ~reservation_i[407];
  assign N197 = reservation_i[408] | reservation_i[409];
  assign N198 = N196 | N197;
  assign N199 = reservation_i[406] | N198;
  assign N200 = reservation_i[405] | N199;
  assign N201 = reservation_i[404] | N200;
  assign N202 = ~N201;
  assign N203 = ~reservation_i[404];
  assign N204 = N203 | N200;
  assign N205 = ~N204;

  divSqrtRecFNToRaw_11_53_2
  fdiv
  (
    .nReset(_12_net_),
    .clock(clk_i),
    .control(1'b1),
    .inReady(fdivsqrt_ready_and_lo),
    .inValid(fdivsqrt_v_li),
    .sqrtOp(fsqrt_v_li),
    .a(reservation_i[194:130]),
    .b(reservation_i[129:65]),
    .roundingMode(frm_li),
    .outValid(fdivsqrt_v_lo),
    .sqrtOpOut(sqrt_lo),
    .roundingModeOut(frm_lo),
    .invalidExc(invalid_exc),
    .infiniteExc(infinite_exc),
    .out_isNaN(fdivsqrt_raw_lo[74]),
    .out_isInf(fdivsqrt_raw_lo[73]),
    .out_isZero(fdivsqrt_raw_lo[72]),
    .out_sign(fdivsqrt_raw_lo[69]),
    .out_sExp(fdivsqrt_raw_lo[68:56]),
    .out_sig(fdivsqrt_raw_lo[55:0])
  );


  bsg_dff_reset_en_width_p1
  fdivsqrt_pending_reg
  (
    .clk_i(clk_i),
    .reset_i(_19_net_),
    .en_i(_20_net_),
    .data_i(_21_net_),
    .data_o(fdivsqrt_pending_r)
  );


  bsg_dff_en_width_p9
  fwb_reg
  (
    .clk_i(clk_i),
    .data_i({ frm_li, reservation_i[460:456], reservation_i[403:403] }),
    .en_i(fdivsqrt_v_li),
    .data_o({ frm_r, fwb_pkt_o[75:71], frd_tag_r })
  );


  bp_be_fp_rebox_00
  rebox
  (
    .raw_i(fdivsqrt_raw_lo),
    .tag_i(frd_tag_r),
    .frm_i(frm_r),
    .invalid_exc_i(invalid_exc),
    .infinite_exc_i(infinite_exc),
    .reg_o(fwb_pkt_o[70:5]),
    .fflags_o({ fflags_lo_nv_, fflags_lo_dz_, fflags_lo_of_, fflags_lo_uf_, fflags_lo_nx_ })
  );

  assign N206 = reservation_i[462] & reservation_i[463];
  assign N207 = reservation_i[461] & N206;
  assign { N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131 } = (N0)? remainder_lo : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N1)? quotient_lo : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N2)? imulh_result_lo : 1'b0;
  assign N0 = N120;
  assign N1 = N125;
  assign N2 = N130;
  assign iresult = (N3)? { N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131 } : 
                   (N112)? imulh_result_lo : 1'b0;
  assign N3 = N111;
  assign frm_li = (N4)? frm_dyn_i : 
                  (N195)? reservation_i[463:461] : 1'b0;
  assign N4 = N207;
  assign int_v_li = N208 & reservation_i[435];
  assign N208 = reservation_i[520] & reservation_i[441];
  assign fp_v_li = N209 & reservation_i[434];
  assign N209 = reservation_i[520] & reservation_i[441];
  assign flush_int_li = flush_i & N210;
  assign N210 = imask_r | int_v_li;
  assign flush_fp_li = flush_i & N211;
  assign N211 = fmask_r | fp_v_li;
  assign imulh_v_li = int_v_li & N81;
  assign _4_net_ = imulh_v_lo & iwb_yumi_i;
  assign _2_net_ = reset_i | flush_int_li;
  assign idiv_v_li = int_v_li & N93;
  assign irem_v_li = int_v_li & N106;
  assign _7_net_ = idiv_v_lo & iwb_yumi_i;
  assign _6_net_ = idiv_v_li | irem_v_li;
  assign _5_net_ = reset_i | flush_int_li;
  assign _8_net_ = N212 | irem_v_li;
  assign N212 = imulh_v_li | idiv_v_li;
  assign N107 = ~fu_op_r[5];
  assign N108 = ~fu_op_r[4];
  assign N109 = ~fu_op_r[3];
  assign N112 = ~N111;
  assign N113 = ~fu_op_r[1];
  assign N114 = ~fu_op_r[0];
  assign N117 = ~fu_op_r[2];
  assign N120 = N213 | N214;
  assign N213 = ~N116;
  assign N214 = ~N119;
  assign N125 = N215 | N216;
  assign N215 = ~N122;
  assign N216 = ~N124;
  assign N130 = N126 | N217;
  assign N217 = N127 | N129;
  assign ibusy_o = N221 | imask_r;
  assign N221 = N219 | N220;
  assign N219 = int_v_li | N218;
  assign N218 = ~imulh_ready_lo;
  assign N220 = ~idiv_ready_and_lo;
  assign iwb_pkt_o_78_ = N222 & N223;
  assign N222 = ~imask_r;
  assign N223 = imulh_v_lo | idiv_v_lo;
  assign N195 = ~N207;
  assign fdiv_v_li = fp_v_li & N202;
  assign fsqrt_v_li = fp_v_li & N205;
  assign fdivsqrt_v_li = fdiv_v_li | fsqrt_v_li;
  assign _12_net_ = N224 & N225;
  assign N224 = ~reset_i;
  assign N225 = ~flush_fp_li;
  assign _21_net_ = fdivsqrt_v_lo & N226;
  assign N226 = ~fwb_yumi_i;
  assign _20_net_ = fdivsqrt_v_lo | fwb_yumi_i;
  assign _19_net_ = reset_i | flush_fp_li;
  assign fdivsqrt_pending = fdivsqrt_v_lo | fdivsqrt_pending_r;
  assign fbusy_o = N229 | fdivsqrt_pending;
  assign N229 = N228 | fmask_r;
  assign N228 = fdivsqrt_v_li | N227;
  assign N227 = ~fdivsqrt_ready_and_lo;
  assign fwb_pkt_o_77_ = N230 & N231;
  assign N230 = ~fmask_r;
  assign N231 = fdivsqrt_v_lo | fdivsqrt_pending;
  assign fwb_pkt_o[4] = fflags_lo_nv_ & fwb_pkt_o_77_;
  assign fwb_pkt_o[3] = fflags_lo_dz_ & fwb_pkt_o_77_;
  assign fwb_pkt_o[2] = fflags_lo_of_ & fwb_pkt_o_77_;
  assign fwb_pkt_o[1] = fflags_lo_uf_ & fwb_pkt_o_77_;
  assign fwb_pkt_o[0] = fflags_lo_nx_ & fwb_pkt_o_77_;

endmodule



module bsg_scan_width_p3_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [2:0] i;
  output [2:0] o;
  wire [2:0] o;
  wire t_1__2_,t_1__1_,t_1__0_;
  assign t_1__2_ = i[0] | 1'b0;
  assign t_1__1_ = i[1] | i[0];
  assign t_1__0_ = i[2] | i[1];
  assign o[0] = t_1__2_ | 1'b0;
  assign o[1] = t_1__1_ | 1'b0;
  assign o[2] = t_1__0_ | t_1__2_;

endmodule



module bsg_priority_encode_one_hot_out_width_p3_lo_to_hi_p1
(
  i,
  o,
  v_o
);

  input [2:0] i;
  output [2:0] o;
  output v_o;
  wire [2:0] o;
  wire v_o,N0,N1;
  wire [1:1] scan_lo;

  bsg_scan_width_p3_or_p1_lo_to_hi_p1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, scan_lo[1:1], o[0:0] })
  );

  assign o[2] = v_o & N0;
  assign N0 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N1;
  assign N1 = ~o[0];

endmodule



module bsg_arb_fixed_inputs_p3_lo_to_hi_p1
(
  ready_then_i,
  reqs_i,
  grants_o
);

  input [2:0] reqs_i;
  output [2:0] grants_o;
  input ready_then_i;
  wire [2:0] grants_o,grants_unmasked_lo;

  bsg_priority_encode_one_hot_out_width_p3_lo_to_hi_p1
  enc
  (
    .i(reqs_i),
    .o(grants_unmasked_lo)
  );

  assign grants_o[2] = grants_unmasked_lo[2] & ready_then_i;
  assign grants_o[1] = grants_unmasked_lo[1] & ready_then_i;
  assign grants_o[0] = grants_unmasked_lo[0] & ready_then_i;

endmodule



module bsg_mux_one_hot_width_p79_els_p3
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [236:0] data_i;
  input [2:0] sel_one_hot_i;
  output [78:0] data_o;
  wire [78:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78;
  wire [236:0] data_masked;
  assign data_masked[78] = data_i[78] & sel_one_hot_i[0];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[0];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[0];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[0];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[0];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[0];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[0];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[0];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[0];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[0];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[0];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[1];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[1];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[1];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[1];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[1];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[1];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[1];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[1];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[1];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[1];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[1];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[1];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[1];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[1];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[1];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[1];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[1];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[1];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[1];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[1];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[1];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[1];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[1];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[1];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[1];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[1];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[1];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[1];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[1];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[1];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[2];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[2];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[2];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[2];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[2];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[2];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[2];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[2];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[2];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[2];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[2];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[2];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[2];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[2];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[2];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[2];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[2];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[2];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[2];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[2];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[2];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[2];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[2];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[2];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[2];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[2];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[2];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[2];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[2];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[2];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[2];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[2];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[2];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[2];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[2];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[2];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[2];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[2];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[2];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[2];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[2];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[2];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[2];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[2];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[2];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[2];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[2];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[2];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[2];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[2];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[2];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[2];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[2];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[2];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[2];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[2];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[2];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[2];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[2];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[2];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[2];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[2];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[2];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[2];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[2];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[2];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[2];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[2];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[2];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[2];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[2];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[2];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[2];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[2];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[2];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[2];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[2];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[2];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[2];
  assign data_o[0] = N0 | data_masked[0];
  assign N0 = data_masked[158] | data_masked[79];
  assign data_o[1] = N1 | data_masked[1];
  assign N1 = data_masked[159] | data_masked[80];
  assign data_o[2] = N2 | data_masked[2];
  assign N2 = data_masked[160] | data_masked[81];
  assign data_o[3] = N3 | data_masked[3];
  assign N3 = data_masked[161] | data_masked[82];
  assign data_o[4] = N4 | data_masked[4];
  assign N4 = data_masked[162] | data_masked[83];
  assign data_o[5] = N5 | data_masked[5];
  assign N5 = data_masked[163] | data_masked[84];
  assign data_o[6] = N6 | data_masked[6];
  assign N6 = data_masked[164] | data_masked[85];
  assign data_o[7] = N7 | data_masked[7];
  assign N7 = data_masked[165] | data_masked[86];
  assign data_o[8] = N8 | data_masked[8];
  assign N8 = data_masked[166] | data_masked[87];
  assign data_o[9] = N9 | data_masked[9];
  assign N9 = data_masked[167] | data_masked[88];
  assign data_o[10] = N10 | data_masked[10];
  assign N10 = data_masked[168] | data_masked[89];
  assign data_o[11] = N11 | data_masked[11];
  assign N11 = data_masked[169] | data_masked[90];
  assign data_o[12] = N12 | data_masked[12];
  assign N12 = data_masked[170] | data_masked[91];
  assign data_o[13] = N13 | data_masked[13];
  assign N13 = data_masked[171] | data_masked[92];
  assign data_o[14] = N14 | data_masked[14];
  assign N14 = data_masked[172] | data_masked[93];
  assign data_o[15] = N15 | data_masked[15];
  assign N15 = data_masked[173] | data_masked[94];
  assign data_o[16] = N16 | data_masked[16];
  assign N16 = data_masked[174] | data_masked[95];
  assign data_o[17] = N17 | data_masked[17];
  assign N17 = data_masked[175] | data_masked[96];
  assign data_o[18] = N18 | data_masked[18];
  assign N18 = data_masked[176] | data_masked[97];
  assign data_o[19] = N19 | data_masked[19];
  assign N19 = data_masked[177] | data_masked[98];
  assign data_o[20] = N20 | data_masked[20];
  assign N20 = data_masked[178] | data_masked[99];
  assign data_o[21] = N21 | data_masked[21];
  assign N21 = data_masked[179] | data_masked[100];
  assign data_o[22] = N22 | data_masked[22];
  assign N22 = data_masked[180] | data_masked[101];
  assign data_o[23] = N23 | data_masked[23];
  assign N23 = data_masked[181] | data_masked[102];
  assign data_o[24] = N24 | data_masked[24];
  assign N24 = data_masked[182] | data_masked[103];
  assign data_o[25] = N25 | data_masked[25];
  assign N25 = data_masked[183] | data_masked[104];
  assign data_o[26] = N26 | data_masked[26];
  assign N26 = data_masked[184] | data_masked[105];
  assign data_o[27] = N27 | data_masked[27];
  assign N27 = data_masked[185] | data_masked[106];
  assign data_o[28] = N28 | data_masked[28];
  assign N28 = data_masked[186] | data_masked[107];
  assign data_o[29] = N29 | data_masked[29];
  assign N29 = data_masked[187] | data_masked[108];
  assign data_o[30] = N30 | data_masked[30];
  assign N30 = data_masked[188] | data_masked[109];
  assign data_o[31] = N31 | data_masked[31];
  assign N31 = data_masked[189] | data_masked[110];
  assign data_o[32] = N32 | data_masked[32];
  assign N32 = data_masked[190] | data_masked[111];
  assign data_o[33] = N33 | data_masked[33];
  assign N33 = data_masked[191] | data_masked[112];
  assign data_o[34] = N34 | data_masked[34];
  assign N34 = data_masked[192] | data_masked[113];
  assign data_o[35] = N35 | data_masked[35];
  assign N35 = data_masked[193] | data_masked[114];
  assign data_o[36] = N36 | data_masked[36];
  assign N36 = data_masked[194] | data_masked[115];
  assign data_o[37] = N37 | data_masked[37];
  assign N37 = data_masked[195] | data_masked[116];
  assign data_o[38] = N38 | data_masked[38];
  assign N38 = data_masked[196] | data_masked[117];
  assign data_o[39] = N39 | data_masked[39];
  assign N39 = data_masked[197] | data_masked[118];
  assign data_o[40] = N40 | data_masked[40];
  assign N40 = data_masked[198] | data_masked[119];
  assign data_o[41] = N41 | data_masked[41];
  assign N41 = data_masked[199] | data_masked[120];
  assign data_o[42] = N42 | data_masked[42];
  assign N42 = data_masked[200] | data_masked[121];
  assign data_o[43] = N43 | data_masked[43];
  assign N43 = data_masked[201] | data_masked[122];
  assign data_o[44] = N44 | data_masked[44];
  assign N44 = data_masked[202] | data_masked[123];
  assign data_o[45] = N45 | data_masked[45];
  assign N45 = data_masked[203] | data_masked[124];
  assign data_o[46] = N46 | data_masked[46];
  assign N46 = data_masked[204] | data_masked[125];
  assign data_o[47] = N47 | data_masked[47];
  assign N47 = data_masked[205] | data_masked[126];
  assign data_o[48] = N48 | data_masked[48];
  assign N48 = data_masked[206] | data_masked[127];
  assign data_o[49] = N49 | data_masked[49];
  assign N49 = data_masked[207] | data_masked[128];
  assign data_o[50] = N50 | data_masked[50];
  assign N50 = data_masked[208] | data_masked[129];
  assign data_o[51] = N51 | data_masked[51];
  assign N51 = data_masked[209] | data_masked[130];
  assign data_o[52] = N52 | data_masked[52];
  assign N52 = data_masked[210] | data_masked[131];
  assign data_o[53] = N53 | data_masked[53];
  assign N53 = data_masked[211] | data_masked[132];
  assign data_o[54] = N54 | data_masked[54];
  assign N54 = data_masked[212] | data_masked[133];
  assign data_o[55] = N55 | data_masked[55];
  assign N55 = data_masked[213] | data_masked[134];
  assign data_o[56] = N56 | data_masked[56];
  assign N56 = data_masked[214] | data_masked[135];
  assign data_o[57] = N57 | data_masked[57];
  assign N57 = data_masked[215] | data_masked[136];
  assign data_o[58] = N58 | data_masked[58];
  assign N58 = data_masked[216] | data_masked[137];
  assign data_o[59] = N59 | data_masked[59];
  assign N59 = data_masked[217] | data_masked[138];
  assign data_o[60] = N60 | data_masked[60];
  assign N60 = data_masked[218] | data_masked[139];
  assign data_o[61] = N61 | data_masked[61];
  assign N61 = data_masked[219] | data_masked[140];
  assign data_o[62] = N62 | data_masked[62];
  assign N62 = data_masked[220] | data_masked[141];
  assign data_o[63] = N63 | data_masked[63];
  assign N63 = data_masked[221] | data_masked[142];
  assign data_o[64] = N64 | data_masked[64];
  assign N64 = data_masked[222] | data_masked[143];
  assign data_o[65] = N65 | data_masked[65];
  assign N65 = data_masked[223] | data_masked[144];
  assign data_o[66] = N66 | data_masked[66];
  assign N66 = data_masked[224] | data_masked[145];
  assign data_o[67] = N67 | data_masked[67];
  assign N67 = data_masked[225] | data_masked[146];
  assign data_o[68] = N68 | data_masked[68];
  assign N68 = data_masked[226] | data_masked[147];
  assign data_o[69] = N69 | data_masked[69];
  assign N69 = data_masked[227] | data_masked[148];
  assign data_o[70] = N70 | data_masked[70];
  assign N70 = data_masked[228] | data_masked[149];
  assign data_o[71] = N71 | data_masked[71];
  assign N71 = data_masked[229] | data_masked[150];
  assign data_o[72] = N72 | data_masked[72];
  assign N72 = data_masked[230] | data_masked[151];
  assign data_o[73] = N73 | data_masked[73];
  assign N73 = data_masked[231] | data_masked[152];
  assign data_o[74] = N74 | data_masked[74];
  assign N74 = data_masked[232] | data_masked[153];
  assign data_o[75] = N75 | data_masked[75];
  assign N75 = data_masked[233] | data_masked[154];
  assign data_o[76] = N76 | data_masked[76];
  assign N76 = data_masked[234] | data_masked[155];
  assign data_o[77] = N77 | data_masked[77];
  assign N77 = data_masked[235] | data_masked[156];
  assign data_o[78] = N78 | data_masked[78];
  assign N78 = data_masked[236] | data_masked[157];

endmodule



module bsg_dff_width_p395
(
  clk_i,
  data_i,
  data_o
);

  input [394:0] data_i;
  output [394:0] data_o;
  input clk_i;
  wire [394:0] data_o;
  reg data_o_394_sv2v_reg,data_o_393_sv2v_reg,data_o_392_sv2v_reg,data_o_391_sv2v_reg,
  data_o_390_sv2v_reg,data_o_389_sv2v_reg,data_o_388_sv2v_reg,data_o_387_sv2v_reg,
  data_o_386_sv2v_reg,data_o_385_sv2v_reg,data_o_384_sv2v_reg,data_o_383_sv2v_reg,
  data_o_382_sv2v_reg,data_o_381_sv2v_reg,data_o_380_sv2v_reg,data_o_379_sv2v_reg,
  data_o_378_sv2v_reg,data_o_377_sv2v_reg,data_o_376_sv2v_reg,data_o_375_sv2v_reg,
  data_o_374_sv2v_reg,data_o_373_sv2v_reg,data_o_372_sv2v_reg,data_o_371_sv2v_reg,
  data_o_370_sv2v_reg,data_o_369_sv2v_reg,data_o_368_sv2v_reg,data_o_367_sv2v_reg,
  data_o_366_sv2v_reg,data_o_365_sv2v_reg,data_o_364_sv2v_reg,data_o_363_sv2v_reg,
  data_o_362_sv2v_reg,data_o_361_sv2v_reg,data_o_360_sv2v_reg,data_o_359_sv2v_reg,
  data_o_358_sv2v_reg,data_o_357_sv2v_reg,data_o_356_sv2v_reg,data_o_355_sv2v_reg,
  data_o_354_sv2v_reg,data_o_353_sv2v_reg,data_o_352_sv2v_reg,data_o_351_sv2v_reg,
  data_o_350_sv2v_reg,data_o_349_sv2v_reg,data_o_348_sv2v_reg,data_o_347_sv2v_reg,
  data_o_346_sv2v_reg,data_o_345_sv2v_reg,data_o_344_sv2v_reg,data_o_343_sv2v_reg,
  data_o_342_sv2v_reg,data_o_341_sv2v_reg,data_o_340_sv2v_reg,data_o_339_sv2v_reg,
  data_o_338_sv2v_reg,data_o_337_sv2v_reg,data_o_336_sv2v_reg,data_o_335_sv2v_reg,
  data_o_334_sv2v_reg,data_o_333_sv2v_reg,data_o_332_sv2v_reg,data_o_331_sv2v_reg,
  data_o_330_sv2v_reg,data_o_329_sv2v_reg,data_o_328_sv2v_reg,data_o_327_sv2v_reg,
  data_o_326_sv2v_reg,data_o_325_sv2v_reg,data_o_324_sv2v_reg,data_o_323_sv2v_reg,
  data_o_322_sv2v_reg,data_o_321_sv2v_reg,data_o_320_sv2v_reg,data_o_319_sv2v_reg,
  data_o_318_sv2v_reg,data_o_317_sv2v_reg,data_o_316_sv2v_reg,data_o_315_sv2v_reg,
  data_o_314_sv2v_reg,data_o_313_sv2v_reg,data_o_312_sv2v_reg,data_o_311_sv2v_reg,
  data_o_310_sv2v_reg,data_o_309_sv2v_reg,data_o_308_sv2v_reg,data_o_307_sv2v_reg,
  data_o_306_sv2v_reg,data_o_305_sv2v_reg,data_o_304_sv2v_reg,data_o_303_sv2v_reg,
  data_o_302_sv2v_reg,data_o_301_sv2v_reg,data_o_300_sv2v_reg,data_o_299_sv2v_reg,
  data_o_298_sv2v_reg,data_o_297_sv2v_reg,data_o_296_sv2v_reg,data_o_295_sv2v_reg,
  data_o_294_sv2v_reg,data_o_293_sv2v_reg,data_o_292_sv2v_reg,data_o_291_sv2v_reg,
  data_o_290_sv2v_reg,data_o_289_sv2v_reg,data_o_288_sv2v_reg,data_o_287_sv2v_reg,
  data_o_286_sv2v_reg,data_o_285_sv2v_reg,data_o_284_sv2v_reg,data_o_283_sv2v_reg,
  data_o_282_sv2v_reg,data_o_281_sv2v_reg,data_o_280_sv2v_reg,data_o_279_sv2v_reg,
  data_o_278_sv2v_reg,data_o_277_sv2v_reg,data_o_276_sv2v_reg,data_o_275_sv2v_reg,
  data_o_274_sv2v_reg,data_o_273_sv2v_reg,data_o_272_sv2v_reg,data_o_271_sv2v_reg,
  data_o_270_sv2v_reg,data_o_269_sv2v_reg,data_o_268_sv2v_reg,data_o_267_sv2v_reg,
  data_o_266_sv2v_reg,data_o_265_sv2v_reg,data_o_264_sv2v_reg,data_o_263_sv2v_reg,
  data_o_262_sv2v_reg,data_o_261_sv2v_reg,data_o_260_sv2v_reg,data_o_259_sv2v_reg,
  data_o_258_sv2v_reg,data_o_257_sv2v_reg,data_o_256_sv2v_reg,data_o_255_sv2v_reg,
  data_o_254_sv2v_reg,data_o_253_sv2v_reg,data_o_252_sv2v_reg,data_o_251_sv2v_reg,
  data_o_250_sv2v_reg,data_o_249_sv2v_reg,data_o_248_sv2v_reg,data_o_247_sv2v_reg,
  data_o_246_sv2v_reg,data_o_245_sv2v_reg,data_o_244_sv2v_reg,data_o_243_sv2v_reg,
  data_o_242_sv2v_reg,data_o_241_sv2v_reg,data_o_240_sv2v_reg,data_o_239_sv2v_reg,
  data_o_238_sv2v_reg,data_o_237_sv2v_reg,data_o_236_sv2v_reg,data_o_235_sv2v_reg,
  data_o_234_sv2v_reg,data_o_233_sv2v_reg,data_o_232_sv2v_reg,data_o_231_sv2v_reg,
  data_o_230_sv2v_reg,data_o_229_sv2v_reg,data_o_228_sv2v_reg,data_o_227_sv2v_reg,
  data_o_226_sv2v_reg,data_o_225_sv2v_reg,data_o_224_sv2v_reg,data_o_223_sv2v_reg,
  data_o_222_sv2v_reg,data_o_221_sv2v_reg,data_o_220_sv2v_reg,data_o_219_sv2v_reg,
  data_o_218_sv2v_reg,data_o_217_sv2v_reg,data_o_216_sv2v_reg,data_o_215_sv2v_reg,
  data_o_214_sv2v_reg,data_o_213_sv2v_reg,data_o_212_sv2v_reg,data_o_211_sv2v_reg,
  data_o_210_sv2v_reg,data_o_209_sv2v_reg,data_o_208_sv2v_reg,data_o_207_sv2v_reg,
  data_o_206_sv2v_reg,data_o_205_sv2v_reg,data_o_204_sv2v_reg,data_o_203_sv2v_reg,
  data_o_202_sv2v_reg,data_o_201_sv2v_reg,data_o_200_sv2v_reg,data_o_199_sv2v_reg,
  data_o_198_sv2v_reg,data_o_197_sv2v_reg,data_o_196_sv2v_reg,data_o_195_sv2v_reg,
  data_o_194_sv2v_reg,data_o_193_sv2v_reg,data_o_192_sv2v_reg,data_o_191_sv2v_reg,
  data_o_190_sv2v_reg,data_o_189_sv2v_reg,data_o_188_sv2v_reg,data_o_187_sv2v_reg,
  data_o_186_sv2v_reg,data_o_185_sv2v_reg,data_o_184_sv2v_reg,data_o_183_sv2v_reg,
  data_o_182_sv2v_reg,data_o_181_sv2v_reg,data_o_180_sv2v_reg,data_o_179_sv2v_reg,
  data_o_178_sv2v_reg,data_o_177_sv2v_reg,data_o_176_sv2v_reg,data_o_175_sv2v_reg,
  data_o_174_sv2v_reg,data_o_173_sv2v_reg,data_o_172_sv2v_reg,data_o_171_sv2v_reg,
  data_o_170_sv2v_reg,data_o_169_sv2v_reg,data_o_168_sv2v_reg,data_o_167_sv2v_reg,
  data_o_166_sv2v_reg,data_o_165_sv2v_reg,data_o_164_sv2v_reg,data_o_163_sv2v_reg,
  data_o_162_sv2v_reg,data_o_161_sv2v_reg,data_o_160_sv2v_reg,data_o_159_sv2v_reg,
  data_o_158_sv2v_reg,data_o_157_sv2v_reg,data_o_156_sv2v_reg,data_o_155_sv2v_reg,
  data_o_154_sv2v_reg,data_o_153_sv2v_reg,data_o_152_sv2v_reg,data_o_151_sv2v_reg,
  data_o_150_sv2v_reg,data_o_149_sv2v_reg,data_o_148_sv2v_reg,data_o_147_sv2v_reg,
  data_o_146_sv2v_reg,data_o_145_sv2v_reg,data_o_144_sv2v_reg,data_o_143_sv2v_reg,
  data_o_142_sv2v_reg,data_o_141_sv2v_reg,data_o_140_sv2v_reg,data_o_139_sv2v_reg,
  data_o_138_sv2v_reg,data_o_137_sv2v_reg,data_o_136_sv2v_reg,data_o_135_sv2v_reg,
  data_o_134_sv2v_reg,data_o_133_sv2v_reg,data_o_132_sv2v_reg,data_o_131_sv2v_reg,
  data_o_130_sv2v_reg,data_o_129_sv2v_reg,data_o_128_sv2v_reg,data_o_127_sv2v_reg,
  data_o_126_sv2v_reg,data_o_125_sv2v_reg,data_o_124_sv2v_reg,data_o_123_sv2v_reg,
  data_o_122_sv2v_reg,data_o_121_sv2v_reg,data_o_120_sv2v_reg,data_o_119_sv2v_reg,
  data_o_118_sv2v_reg,data_o_117_sv2v_reg,data_o_116_sv2v_reg,data_o_115_sv2v_reg,
  data_o_114_sv2v_reg,data_o_113_sv2v_reg,data_o_112_sv2v_reg,data_o_111_sv2v_reg,
  data_o_110_sv2v_reg,data_o_109_sv2v_reg,data_o_108_sv2v_reg,data_o_107_sv2v_reg,
  data_o_106_sv2v_reg,data_o_105_sv2v_reg,data_o_104_sv2v_reg,data_o_103_sv2v_reg,
  data_o_102_sv2v_reg,data_o_101_sv2v_reg,data_o_100_sv2v_reg,data_o_99_sv2v_reg,
  data_o_98_sv2v_reg,data_o_97_sv2v_reg,data_o_96_sv2v_reg,data_o_95_sv2v_reg,
  data_o_94_sv2v_reg,data_o_93_sv2v_reg,data_o_92_sv2v_reg,data_o_91_sv2v_reg,
  data_o_90_sv2v_reg,data_o_89_sv2v_reg,data_o_88_sv2v_reg,data_o_87_sv2v_reg,
  data_o_86_sv2v_reg,data_o_85_sv2v_reg,data_o_84_sv2v_reg,data_o_83_sv2v_reg,
  data_o_82_sv2v_reg,data_o_81_sv2v_reg,data_o_80_sv2v_reg,data_o_79_sv2v_reg,data_o_78_sv2v_reg,
  data_o_77_sv2v_reg,data_o_76_sv2v_reg,data_o_75_sv2v_reg,data_o_74_sv2v_reg,
  data_o_73_sv2v_reg,data_o_72_sv2v_reg,data_o_71_sv2v_reg,data_o_70_sv2v_reg,
  data_o_69_sv2v_reg,data_o_68_sv2v_reg,data_o_67_sv2v_reg,data_o_66_sv2v_reg,
  data_o_65_sv2v_reg,data_o_64_sv2v_reg,data_o_63_sv2v_reg,data_o_62_sv2v_reg,
  data_o_61_sv2v_reg,data_o_60_sv2v_reg,data_o_59_sv2v_reg,data_o_58_sv2v_reg,data_o_57_sv2v_reg,
  data_o_56_sv2v_reg,data_o_55_sv2v_reg,data_o_54_sv2v_reg,data_o_53_sv2v_reg,
  data_o_52_sv2v_reg,data_o_51_sv2v_reg,data_o_50_sv2v_reg,data_o_49_sv2v_reg,
  data_o_48_sv2v_reg,data_o_47_sv2v_reg,data_o_46_sv2v_reg,data_o_45_sv2v_reg,
  data_o_44_sv2v_reg,data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,
  data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,
  data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,
  data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,
  data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,
  data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[394] = data_o_394_sv2v_reg;
  assign data_o[393] = data_o_393_sv2v_reg;
  assign data_o[392] = data_o_392_sv2v_reg;
  assign data_o[391] = data_o_391_sv2v_reg;
  assign data_o[390] = data_o_390_sv2v_reg;
  assign data_o[389] = data_o_389_sv2v_reg;
  assign data_o[388] = data_o_388_sv2v_reg;
  assign data_o[387] = data_o_387_sv2v_reg;
  assign data_o[386] = data_o_386_sv2v_reg;
  assign data_o[385] = data_o_385_sv2v_reg;
  assign data_o[384] = data_o_384_sv2v_reg;
  assign data_o[383] = data_o_383_sv2v_reg;
  assign data_o[382] = data_o_382_sv2v_reg;
  assign data_o[381] = data_o_381_sv2v_reg;
  assign data_o[380] = data_o_380_sv2v_reg;
  assign data_o[379] = data_o_379_sv2v_reg;
  assign data_o[378] = data_o_378_sv2v_reg;
  assign data_o[377] = data_o_377_sv2v_reg;
  assign data_o[376] = data_o_376_sv2v_reg;
  assign data_o[375] = data_o_375_sv2v_reg;
  assign data_o[374] = data_o_374_sv2v_reg;
  assign data_o[373] = data_o_373_sv2v_reg;
  assign data_o[372] = data_o_372_sv2v_reg;
  assign data_o[371] = data_o_371_sv2v_reg;
  assign data_o[370] = data_o_370_sv2v_reg;
  assign data_o[369] = data_o_369_sv2v_reg;
  assign data_o[368] = data_o_368_sv2v_reg;
  assign data_o[367] = data_o_367_sv2v_reg;
  assign data_o[366] = data_o_366_sv2v_reg;
  assign data_o[365] = data_o_365_sv2v_reg;
  assign data_o[364] = data_o_364_sv2v_reg;
  assign data_o[363] = data_o_363_sv2v_reg;
  assign data_o[362] = data_o_362_sv2v_reg;
  assign data_o[361] = data_o_361_sv2v_reg;
  assign data_o[360] = data_o_360_sv2v_reg;
  assign data_o[359] = data_o_359_sv2v_reg;
  assign data_o[358] = data_o_358_sv2v_reg;
  assign data_o[357] = data_o_357_sv2v_reg;
  assign data_o[356] = data_o_356_sv2v_reg;
  assign data_o[355] = data_o_355_sv2v_reg;
  assign data_o[354] = data_o_354_sv2v_reg;
  assign data_o[353] = data_o_353_sv2v_reg;
  assign data_o[352] = data_o_352_sv2v_reg;
  assign data_o[351] = data_o_351_sv2v_reg;
  assign data_o[350] = data_o_350_sv2v_reg;
  assign data_o[349] = data_o_349_sv2v_reg;
  assign data_o[348] = data_o_348_sv2v_reg;
  assign data_o[347] = data_o_347_sv2v_reg;
  assign data_o[346] = data_o_346_sv2v_reg;
  assign data_o[345] = data_o_345_sv2v_reg;
  assign data_o[344] = data_o_344_sv2v_reg;
  assign data_o[343] = data_o_343_sv2v_reg;
  assign data_o[342] = data_o_342_sv2v_reg;
  assign data_o[341] = data_o_341_sv2v_reg;
  assign data_o[340] = data_o_340_sv2v_reg;
  assign data_o[339] = data_o_339_sv2v_reg;
  assign data_o[338] = data_o_338_sv2v_reg;
  assign data_o[337] = data_o_337_sv2v_reg;
  assign data_o[336] = data_o_336_sv2v_reg;
  assign data_o[335] = data_o_335_sv2v_reg;
  assign data_o[334] = data_o_334_sv2v_reg;
  assign data_o[333] = data_o_333_sv2v_reg;
  assign data_o[332] = data_o_332_sv2v_reg;
  assign data_o[331] = data_o_331_sv2v_reg;
  assign data_o[330] = data_o_330_sv2v_reg;
  assign data_o[329] = data_o_329_sv2v_reg;
  assign data_o[328] = data_o_328_sv2v_reg;
  assign data_o[327] = data_o_327_sv2v_reg;
  assign data_o[326] = data_o_326_sv2v_reg;
  assign data_o[325] = data_o_325_sv2v_reg;
  assign data_o[324] = data_o_324_sv2v_reg;
  assign data_o[323] = data_o_323_sv2v_reg;
  assign data_o[322] = data_o_322_sv2v_reg;
  assign data_o[321] = data_o_321_sv2v_reg;
  assign data_o[320] = data_o_320_sv2v_reg;
  assign data_o[319] = data_o_319_sv2v_reg;
  assign data_o[318] = data_o_318_sv2v_reg;
  assign data_o[317] = data_o_317_sv2v_reg;
  assign data_o[316] = data_o_316_sv2v_reg;
  assign data_o[315] = data_o_315_sv2v_reg;
  assign data_o[314] = data_o_314_sv2v_reg;
  assign data_o[313] = data_o_313_sv2v_reg;
  assign data_o[312] = data_o_312_sv2v_reg;
  assign data_o[311] = data_o_311_sv2v_reg;
  assign data_o[310] = data_o_310_sv2v_reg;
  assign data_o[309] = data_o_309_sv2v_reg;
  assign data_o[308] = data_o_308_sv2v_reg;
  assign data_o[307] = data_o_307_sv2v_reg;
  assign data_o[306] = data_o_306_sv2v_reg;
  assign data_o[305] = data_o_305_sv2v_reg;
  assign data_o[304] = data_o_304_sv2v_reg;
  assign data_o[303] = data_o_303_sv2v_reg;
  assign data_o[302] = data_o_302_sv2v_reg;
  assign data_o[301] = data_o_301_sv2v_reg;
  assign data_o[300] = data_o_300_sv2v_reg;
  assign data_o[299] = data_o_299_sv2v_reg;
  assign data_o[298] = data_o_298_sv2v_reg;
  assign data_o[297] = data_o_297_sv2v_reg;
  assign data_o[296] = data_o_296_sv2v_reg;
  assign data_o[295] = data_o_295_sv2v_reg;
  assign data_o[294] = data_o_294_sv2v_reg;
  assign data_o[293] = data_o_293_sv2v_reg;
  assign data_o[292] = data_o_292_sv2v_reg;
  assign data_o[291] = data_o_291_sv2v_reg;
  assign data_o[290] = data_o_290_sv2v_reg;
  assign data_o[289] = data_o_289_sv2v_reg;
  assign data_o[288] = data_o_288_sv2v_reg;
  assign data_o[287] = data_o_287_sv2v_reg;
  assign data_o[286] = data_o_286_sv2v_reg;
  assign data_o[285] = data_o_285_sv2v_reg;
  assign data_o[284] = data_o_284_sv2v_reg;
  assign data_o[283] = data_o_283_sv2v_reg;
  assign data_o[282] = data_o_282_sv2v_reg;
  assign data_o[281] = data_o_281_sv2v_reg;
  assign data_o[280] = data_o_280_sv2v_reg;
  assign data_o[279] = data_o_279_sv2v_reg;
  assign data_o[278] = data_o_278_sv2v_reg;
  assign data_o[277] = data_o_277_sv2v_reg;
  assign data_o[276] = data_o_276_sv2v_reg;
  assign data_o[275] = data_o_275_sv2v_reg;
  assign data_o[274] = data_o_274_sv2v_reg;
  assign data_o[273] = data_o_273_sv2v_reg;
  assign data_o[272] = data_o_272_sv2v_reg;
  assign data_o[271] = data_o_271_sv2v_reg;
  assign data_o[270] = data_o_270_sv2v_reg;
  assign data_o[269] = data_o_269_sv2v_reg;
  assign data_o[268] = data_o_268_sv2v_reg;
  assign data_o[267] = data_o_267_sv2v_reg;
  assign data_o[266] = data_o_266_sv2v_reg;
  assign data_o[265] = data_o_265_sv2v_reg;
  assign data_o[264] = data_o_264_sv2v_reg;
  assign data_o[263] = data_o_263_sv2v_reg;
  assign data_o[262] = data_o_262_sv2v_reg;
  assign data_o[261] = data_o_261_sv2v_reg;
  assign data_o[260] = data_o_260_sv2v_reg;
  assign data_o[259] = data_o_259_sv2v_reg;
  assign data_o[258] = data_o_258_sv2v_reg;
  assign data_o[257] = data_o_257_sv2v_reg;
  assign data_o[256] = data_o_256_sv2v_reg;
  assign data_o[255] = data_o_255_sv2v_reg;
  assign data_o[254] = data_o_254_sv2v_reg;
  assign data_o[253] = data_o_253_sv2v_reg;
  assign data_o[252] = data_o_252_sv2v_reg;
  assign data_o[251] = data_o_251_sv2v_reg;
  assign data_o[250] = data_o_250_sv2v_reg;
  assign data_o[249] = data_o_249_sv2v_reg;
  assign data_o[248] = data_o_248_sv2v_reg;
  assign data_o[247] = data_o_247_sv2v_reg;
  assign data_o[246] = data_o_246_sv2v_reg;
  assign data_o[245] = data_o_245_sv2v_reg;
  assign data_o[244] = data_o_244_sv2v_reg;
  assign data_o[243] = data_o_243_sv2v_reg;
  assign data_o[242] = data_o_242_sv2v_reg;
  assign data_o[241] = data_o_241_sv2v_reg;
  assign data_o[240] = data_o_240_sv2v_reg;
  assign data_o[239] = data_o_239_sv2v_reg;
  assign data_o[238] = data_o_238_sv2v_reg;
  assign data_o[237] = data_o_237_sv2v_reg;
  assign data_o[236] = data_o_236_sv2v_reg;
  assign data_o[235] = data_o_235_sv2v_reg;
  assign data_o[234] = data_o_234_sv2v_reg;
  assign data_o[233] = data_o_233_sv2v_reg;
  assign data_o[232] = data_o_232_sv2v_reg;
  assign data_o[231] = data_o_231_sv2v_reg;
  assign data_o[230] = data_o_230_sv2v_reg;
  assign data_o[229] = data_o_229_sv2v_reg;
  assign data_o[228] = data_o_228_sv2v_reg;
  assign data_o[227] = data_o_227_sv2v_reg;
  assign data_o[226] = data_o_226_sv2v_reg;
  assign data_o[225] = data_o_225_sv2v_reg;
  assign data_o[224] = data_o_224_sv2v_reg;
  assign data_o[223] = data_o_223_sv2v_reg;
  assign data_o[222] = data_o_222_sv2v_reg;
  assign data_o[221] = data_o_221_sv2v_reg;
  assign data_o[220] = data_o_220_sv2v_reg;
  assign data_o[219] = data_o_219_sv2v_reg;
  assign data_o[218] = data_o_218_sv2v_reg;
  assign data_o[217] = data_o_217_sv2v_reg;
  assign data_o[216] = data_o_216_sv2v_reg;
  assign data_o[215] = data_o_215_sv2v_reg;
  assign data_o[214] = data_o_214_sv2v_reg;
  assign data_o[213] = data_o_213_sv2v_reg;
  assign data_o[212] = data_o_212_sv2v_reg;
  assign data_o[211] = data_o_211_sv2v_reg;
  assign data_o[210] = data_o_210_sv2v_reg;
  assign data_o[209] = data_o_209_sv2v_reg;
  assign data_o[208] = data_o_208_sv2v_reg;
  assign data_o[207] = data_o_207_sv2v_reg;
  assign data_o[206] = data_o_206_sv2v_reg;
  assign data_o[205] = data_o_205_sv2v_reg;
  assign data_o[204] = data_o_204_sv2v_reg;
  assign data_o[203] = data_o_203_sv2v_reg;
  assign data_o[202] = data_o_202_sv2v_reg;
  assign data_o[201] = data_o_201_sv2v_reg;
  assign data_o[200] = data_o_200_sv2v_reg;
  assign data_o[199] = data_o_199_sv2v_reg;
  assign data_o[198] = data_o_198_sv2v_reg;
  assign data_o[197] = data_o_197_sv2v_reg;
  assign data_o[196] = data_o_196_sv2v_reg;
  assign data_o[195] = data_o_195_sv2v_reg;
  assign data_o[194] = data_o_194_sv2v_reg;
  assign data_o[193] = data_o_193_sv2v_reg;
  assign data_o[192] = data_o_192_sv2v_reg;
  assign data_o[191] = data_o_191_sv2v_reg;
  assign data_o[190] = data_o_190_sv2v_reg;
  assign data_o[189] = data_o_189_sv2v_reg;
  assign data_o[188] = data_o_188_sv2v_reg;
  assign data_o[187] = data_o_187_sv2v_reg;
  assign data_o[186] = data_o_186_sv2v_reg;
  assign data_o[185] = data_o_185_sv2v_reg;
  assign data_o[184] = data_o_184_sv2v_reg;
  assign data_o[183] = data_o_183_sv2v_reg;
  assign data_o[182] = data_o_182_sv2v_reg;
  assign data_o[181] = data_o_181_sv2v_reg;
  assign data_o[180] = data_o_180_sv2v_reg;
  assign data_o[179] = data_o_179_sv2v_reg;
  assign data_o[178] = data_o_178_sv2v_reg;
  assign data_o[177] = data_o_177_sv2v_reg;
  assign data_o[176] = data_o_176_sv2v_reg;
  assign data_o[175] = data_o_175_sv2v_reg;
  assign data_o[174] = data_o_174_sv2v_reg;
  assign data_o[173] = data_o_173_sv2v_reg;
  assign data_o[172] = data_o_172_sv2v_reg;
  assign data_o[171] = data_o_171_sv2v_reg;
  assign data_o[170] = data_o_170_sv2v_reg;
  assign data_o[169] = data_o_169_sv2v_reg;
  assign data_o[168] = data_o_168_sv2v_reg;
  assign data_o[167] = data_o_167_sv2v_reg;
  assign data_o[166] = data_o_166_sv2v_reg;
  assign data_o[165] = data_o_165_sv2v_reg;
  assign data_o[164] = data_o_164_sv2v_reg;
  assign data_o[163] = data_o_163_sv2v_reg;
  assign data_o[162] = data_o_162_sv2v_reg;
  assign data_o[161] = data_o_161_sv2v_reg;
  assign data_o[160] = data_o_160_sv2v_reg;
  assign data_o[159] = data_o_159_sv2v_reg;
  assign data_o[158] = data_o_158_sv2v_reg;
  assign data_o[157] = data_o_157_sv2v_reg;
  assign data_o[156] = data_o_156_sv2v_reg;
  assign data_o[155] = data_o_155_sv2v_reg;
  assign data_o[154] = data_o_154_sv2v_reg;
  assign data_o[153] = data_o_153_sv2v_reg;
  assign data_o[152] = data_o_152_sv2v_reg;
  assign data_o[151] = data_o_151_sv2v_reg;
  assign data_o[150] = data_o_150_sv2v_reg;
  assign data_o[149] = data_o_149_sv2v_reg;
  assign data_o[148] = data_o_148_sv2v_reg;
  assign data_o[147] = data_o_147_sv2v_reg;
  assign data_o[146] = data_o_146_sv2v_reg;
  assign data_o[145] = data_o_145_sv2v_reg;
  assign data_o[144] = data_o_144_sv2v_reg;
  assign data_o[143] = data_o_143_sv2v_reg;
  assign data_o[142] = data_o_142_sv2v_reg;
  assign data_o[141] = data_o_141_sv2v_reg;
  assign data_o[140] = data_o_140_sv2v_reg;
  assign data_o[139] = data_o_139_sv2v_reg;
  assign data_o[138] = data_o_138_sv2v_reg;
  assign data_o[137] = data_o_137_sv2v_reg;
  assign data_o[136] = data_o_136_sv2v_reg;
  assign data_o[135] = data_o_135_sv2v_reg;
  assign data_o[134] = data_o_134_sv2v_reg;
  assign data_o[133] = data_o_133_sv2v_reg;
  assign data_o[132] = data_o_132_sv2v_reg;
  assign data_o[131] = data_o_131_sv2v_reg;
  assign data_o[130] = data_o_130_sv2v_reg;
  assign data_o[129] = data_o_129_sv2v_reg;
  assign data_o[128] = data_o_128_sv2v_reg;
  assign data_o[127] = data_o_127_sv2v_reg;
  assign data_o[126] = data_o_126_sv2v_reg;
  assign data_o[125] = data_o_125_sv2v_reg;
  assign data_o[124] = data_o_124_sv2v_reg;
  assign data_o[123] = data_o_123_sv2v_reg;
  assign data_o[122] = data_o_122_sv2v_reg;
  assign data_o[121] = data_o_121_sv2v_reg;
  assign data_o[120] = data_o_120_sv2v_reg;
  assign data_o[119] = data_o_119_sv2v_reg;
  assign data_o[118] = data_o_118_sv2v_reg;
  assign data_o[117] = data_o_117_sv2v_reg;
  assign data_o[116] = data_o_116_sv2v_reg;
  assign data_o[115] = data_o_115_sv2v_reg;
  assign data_o[114] = data_o_114_sv2v_reg;
  assign data_o[113] = data_o_113_sv2v_reg;
  assign data_o[112] = data_o_112_sv2v_reg;
  assign data_o[111] = data_o_111_sv2v_reg;
  assign data_o[110] = data_o_110_sv2v_reg;
  assign data_o[109] = data_o_109_sv2v_reg;
  assign data_o[108] = data_o_108_sv2v_reg;
  assign data_o[107] = data_o_107_sv2v_reg;
  assign data_o[106] = data_o_106_sv2v_reg;
  assign data_o[105] = data_o_105_sv2v_reg;
  assign data_o[104] = data_o_104_sv2v_reg;
  assign data_o[103] = data_o_103_sv2v_reg;
  assign data_o[102] = data_o_102_sv2v_reg;
  assign data_o[101] = data_o_101_sv2v_reg;
  assign data_o[100] = data_o_100_sv2v_reg;
  assign data_o[99] = data_o_99_sv2v_reg;
  assign data_o[98] = data_o_98_sv2v_reg;
  assign data_o[97] = data_o_97_sv2v_reg;
  assign data_o[96] = data_o_96_sv2v_reg;
  assign data_o[95] = data_o_95_sv2v_reg;
  assign data_o[94] = data_o_94_sv2v_reg;
  assign data_o[93] = data_o_93_sv2v_reg;
  assign data_o[92] = data_o_92_sv2v_reg;
  assign data_o[91] = data_o_91_sv2v_reg;
  assign data_o[90] = data_o_90_sv2v_reg;
  assign data_o[89] = data_o_89_sv2v_reg;
  assign data_o[88] = data_o_88_sv2v_reg;
  assign data_o[87] = data_o_87_sv2v_reg;
  assign data_o[86] = data_o_86_sv2v_reg;
  assign data_o[85] = data_o_85_sv2v_reg;
  assign data_o[84] = data_o_84_sv2v_reg;
  assign data_o[83] = data_o_83_sv2v_reg;
  assign data_o[82] = data_o_82_sv2v_reg;
  assign data_o[81] = data_o_81_sv2v_reg;
  assign data_o[80] = data_o_80_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_394_sv2v_reg <= data_i[394];
      data_o_393_sv2v_reg <= data_i[393];
      data_o_392_sv2v_reg <= data_i[392];
      data_o_391_sv2v_reg <= data_i[391];
      data_o_390_sv2v_reg <= data_i[390];
      data_o_389_sv2v_reg <= data_i[389];
      data_o_388_sv2v_reg <= data_i[388];
      data_o_387_sv2v_reg <= data_i[387];
      data_o_386_sv2v_reg <= data_i[386];
      data_o_385_sv2v_reg <= data_i[385];
      data_o_384_sv2v_reg <= data_i[384];
      data_o_383_sv2v_reg <= data_i[383];
      data_o_382_sv2v_reg <= data_i[382];
      data_o_381_sv2v_reg <= data_i[381];
      data_o_380_sv2v_reg <= data_i[380];
      data_o_379_sv2v_reg <= data_i[379];
      data_o_378_sv2v_reg <= data_i[378];
      data_o_377_sv2v_reg <= data_i[377];
      data_o_376_sv2v_reg <= data_i[376];
      data_o_375_sv2v_reg <= data_i[375];
      data_o_374_sv2v_reg <= data_i[374];
      data_o_373_sv2v_reg <= data_i[373];
      data_o_372_sv2v_reg <= data_i[372];
      data_o_371_sv2v_reg <= data_i[371];
      data_o_370_sv2v_reg <= data_i[370];
      data_o_369_sv2v_reg <= data_i[369];
      data_o_368_sv2v_reg <= data_i[368];
      data_o_367_sv2v_reg <= data_i[367];
      data_o_366_sv2v_reg <= data_i[366];
      data_o_365_sv2v_reg <= data_i[365];
      data_o_364_sv2v_reg <= data_i[364];
      data_o_363_sv2v_reg <= data_i[363];
      data_o_362_sv2v_reg <= data_i[362];
      data_o_361_sv2v_reg <= data_i[361];
      data_o_360_sv2v_reg <= data_i[360];
      data_o_359_sv2v_reg <= data_i[359];
      data_o_358_sv2v_reg <= data_i[358];
      data_o_357_sv2v_reg <= data_i[357];
      data_o_356_sv2v_reg <= data_i[356];
      data_o_355_sv2v_reg <= data_i[355];
      data_o_354_sv2v_reg <= data_i[354];
      data_o_353_sv2v_reg <= data_i[353];
      data_o_352_sv2v_reg <= data_i[352];
      data_o_351_sv2v_reg <= data_i[351];
      data_o_350_sv2v_reg <= data_i[350];
      data_o_349_sv2v_reg <= data_i[349];
      data_o_348_sv2v_reg <= data_i[348];
      data_o_347_sv2v_reg <= data_i[347];
      data_o_346_sv2v_reg <= data_i[346];
      data_o_345_sv2v_reg <= data_i[345];
      data_o_344_sv2v_reg <= data_i[344];
      data_o_343_sv2v_reg <= data_i[343];
      data_o_342_sv2v_reg <= data_i[342];
      data_o_341_sv2v_reg <= data_i[341];
      data_o_340_sv2v_reg <= data_i[340];
      data_o_339_sv2v_reg <= data_i[339];
      data_o_338_sv2v_reg <= data_i[338];
      data_o_337_sv2v_reg <= data_i[337];
      data_o_336_sv2v_reg <= data_i[336];
      data_o_335_sv2v_reg <= data_i[335];
      data_o_334_sv2v_reg <= data_i[334];
      data_o_333_sv2v_reg <= data_i[333];
      data_o_332_sv2v_reg <= data_i[332];
      data_o_331_sv2v_reg <= data_i[331];
      data_o_330_sv2v_reg <= data_i[330];
      data_o_329_sv2v_reg <= data_i[329];
      data_o_328_sv2v_reg <= data_i[328];
      data_o_327_sv2v_reg <= data_i[327];
      data_o_326_sv2v_reg <= data_i[326];
      data_o_325_sv2v_reg <= data_i[325];
      data_o_324_sv2v_reg <= data_i[324];
      data_o_323_sv2v_reg <= data_i[323];
      data_o_322_sv2v_reg <= data_i[322];
      data_o_321_sv2v_reg <= data_i[321];
      data_o_320_sv2v_reg <= data_i[320];
      data_o_319_sv2v_reg <= data_i[319];
      data_o_318_sv2v_reg <= data_i[318];
      data_o_317_sv2v_reg <= data_i[317];
      data_o_316_sv2v_reg <= data_i[316];
      data_o_315_sv2v_reg <= data_i[315];
      data_o_314_sv2v_reg <= data_i[314];
      data_o_313_sv2v_reg <= data_i[313];
      data_o_312_sv2v_reg <= data_i[312];
      data_o_311_sv2v_reg <= data_i[311];
      data_o_310_sv2v_reg <= data_i[310];
      data_o_309_sv2v_reg <= data_i[309];
      data_o_308_sv2v_reg <= data_i[308];
      data_o_307_sv2v_reg <= data_i[307];
      data_o_306_sv2v_reg <= data_i[306];
      data_o_305_sv2v_reg <= data_i[305];
      data_o_304_sv2v_reg <= data_i[304];
      data_o_303_sv2v_reg <= data_i[303];
      data_o_302_sv2v_reg <= data_i[302];
      data_o_301_sv2v_reg <= data_i[301];
      data_o_300_sv2v_reg <= data_i[300];
      data_o_299_sv2v_reg <= data_i[299];
      data_o_298_sv2v_reg <= data_i[298];
      data_o_297_sv2v_reg <= data_i[297];
      data_o_296_sv2v_reg <= data_i[296];
      data_o_295_sv2v_reg <= data_i[295];
      data_o_294_sv2v_reg <= data_i[294];
      data_o_293_sv2v_reg <= data_i[293];
      data_o_292_sv2v_reg <= data_i[292];
      data_o_291_sv2v_reg <= data_i[291];
      data_o_290_sv2v_reg <= data_i[290];
      data_o_289_sv2v_reg <= data_i[289];
      data_o_288_sv2v_reg <= data_i[288];
      data_o_287_sv2v_reg <= data_i[287];
      data_o_286_sv2v_reg <= data_i[286];
      data_o_285_sv2v_reg <= data_i[285];
      data_o_284_sv2v_reg <= data_i[284];
      data_o_283_sv2v_reg <= data_i[283];
      data_o_282_sv2v_reg <= data_i[282];
      data_o_281_sv2v_reg <= data_i[281];
      data_o_280_sv2v_reg <= data_i[280];
      data_o_279_sv2v_reg <= data_i[279];
      data_o_278_sv2v_reg <= data_i[278];
      data_o_277_sv2v_reg <= data_i[277];
      data_o_276_sv2v_reg <= data_i[276];
      data_o_275_sv2v_reg <= data_i[275];
      data_o_274_sv2v_reg <= data_i[274];
      data_o_273_sv2v_reg <= data_i[273];
      data_o_272_sv2v_reg <= data_i[272];
      data_o_271_sv2v_reg <= data_i[271];
      data_o_270_sv2v_reg <= data_i[270];
      data_o_269_sv2v_reg <= data_i[269];
      data_o_268_sv2v_reg <= data_i[268];
      data_o_267_sv2v_reg <= data_i[267];
      data_o_266_sv2v_reg <= data_i[266];
      data_o_265_sv2v_reg <= data_i[265];
      data_o_264_sv2v_reg <= data_i[264];
      data_o_263_sv2v_reg <= data_i[263];
      data_o_262_sv2v_reg <= data_i[262];
      data_o_261_sv2v_reg <= data_i[261];
      data_o_260_sv2v_reg <= data_i[260];
      data_o_259_sv2v_reg <= data_i[259];
      data_o_258_sv2v_reg <= data_i[258];
      data_o_257_sv2v_reg <= data_i[257];
      data_o_256_sv2v_reg <= data_i[256];
      data_o_255_sv2v_reg <= data_i[255];
      data_o_254_sv2v_reg <= data_i[254];
      data_o_253_sv2v_reg <= data_i[253];
      data_o_252_sv2v_reg <= data_i[252];
      data_o_251_sv2v_reg <= data_i[251];
      data_o_250_sv2v_reg <= data_i[250];
      data_o_249_sv2v_reg <= data_i[249];
      data_o_248_sv2v_reg <= data_i[248];
      data_o_247_sv2v_reg <= data_i[247];
      data_o_246_sv2v_reg <= data_i[246];
      data_o_245_sv2v_reg <= data_i[245];
      data_o_244_sv2v_reg <= data_i[244];
      data_o_243_sv2v_reg <= data_i[243];
      data_o_242_sv2v_reg <= data_i[242];
      data_o_241_sv2v_reg <= data_i[241];
      data_o_240_sv2v_reg <= data_i[240];
      data_o_239_sv2v_reg <= data_i[239];
      data_o_238_sv2v_reg <= data_i[238];
      data_o_237_sv2v_reg <= data_i[237];
      data_o_236_sv2v_reg <= data_i[236];
      data_o_235_sv2v_reg <= data_i[235];
      data_o_234_sv2v_reg <= data_i[234];
      data_o_233_sv2v_reg <= data_i[233];
      data_o_232_sv2v_reg <= data_i[232];
      data_o_231_sv2v_reg <= data_i[231];
      data_o_230_sv2v_reg <= data_i[230];
      data_o_229_sv2v_reg <= data_i[229];
      data_o_228_sv2v_reg <= data_i[228];
      data_o_227_sv2v_reg <= data_i[227];
      data_o_226_sv2v_reg <= data_i[226];
      data_o_225_sv2v_reg <= data_i[225];
      data_o_224_sv2v_reg <= data_i[224];
      data_o_223_sv2v_reg <= data_i[223];
      data_o_222_sv2v_reg <= data_i[222];
      data_o_221_sv2v_reg <= data_i[221];
      data_o_220_sv2v_reg <= data_i[220];
      data_o_219_sv2v_reg <= data_i[219];
      data_o_218_sv2v_reg <= data_i[218];
      data_o_217_sv2v_reg <= data_i[217];
      data_o_216_sv2v_reg <= data_i[216];
      data_o_215_sv2v_reg <= data_i[215];
      data_o_214_sv2v_reg <= data_i[214];
      data_o_213_sv2v_reg <= data_i[213];
      data_o_212_sv2v_reg <= data_i[212];
      data_o_211_sv2v_reg <= data_i[211];
      data_o_210_sv2v_reg <= data_i[210];
      data_o_209_sv2v_reg <= data_i[209];
      data_o_208_sv2v_reg <= data_i[208];
      data_o_207_sv2v_reg <= data_i[207];
      data_o_206_sv2v_reg <= data_i[206];
      data_o_205_sv2v_reg <= data_i[205];
      data_o_204_sv2v_reg <= data_i[204];
      data_o_203_sv2v_reg <= data_i[203];
      data_o_202_sv2v_reg <= data_i[202];
      data_o_201_sv2v_reg <= data_i[201];
      data_o_200_sv2v_reg <= data_i[200];
      data_o_199_sv2v_reg <= data_i[199];
      data_o_198_sv2v_reg <= data_i[198];
      data_o_197_sv2v_reg <= data_i[197];
      data_o_196_sv2v_reg <= data_i[196];
      data_o_195_sv2v_reg <= data_i[195];
      data_o_194_sv2v_reg <= data_i[194];
      data_o_193_sv2v_reg <= data_i[193];
      data_o_192_sv2v_reg <= data_i[192];
      data_o_191_sv2v_reg <= data_i[191];
      data_o_190_sv2v_reg <= data_i[190];
      data_o_189_sv2v_reg <= data_i[189];
      data_o_188_sv2v_reg <= data_i[188];
      data_o_187_sv2v_reg <= data_i[187];
      data_o_186_sv2v_reg <= data_i[186];
      data_o_185_sv2v_reg <= data_i[185];
      data_o_184_sv2v_reg <= data_i[184];
      data_o_183_sv2v_reg <= data_i[183];
      data_o_182_sv2v_reg <= data_i[182];
      data_o_181_sv2v_reg <= data_i[181];
      data_o_180_sv2v_reg <= data_i[180];
      data_o_179_sv2v_reg <= data_i[179];
      data_o_178_sv2v_reg <= data_i[178];
      data_o_177_sv2v_reg <= data_i[177];
      data_o_176_sv2v_reg <= data_i[176];
      data_o_175_sv2v_reg <= data_i[175];
      data_o_174_sv2v_reg <= data_i[174];
      data_o_173_sv2v_reg <= data_i[173];
      data_o_172_sv2v_reg <= data_i[172];
      data_o_171_sv2v_reg <= data_i[171];
      data_o_170_sv2v_reg <= data_i[170];
      data_o_169_sv2v_reg <= data_i[169];
      data_o_168_sv2v_reg <= data_i[168];
      data_o_167_sv2v_reg <= data_i[167];
      data_o_166_sv2v_reg <= data_i[166];
      data_o_165_sv2v_reg <= data_i[165];
      data_o_164_sv2v_reg <= data_i[164];
      data_o_163_sv2v_reg <= data_i[163];
      data_o_162_sv2v_reg <= data_i[162];
      data_o_161_sv2v_reg <= data_i[161];
      data_o_160_sv2v_reg <= data_i[160];
      data_o_159_sv2v_reg <= data_i[159];
      data_o_158_sv2v_reg <= data_i[158];
      data_o_157_sv2v_reg <= data_i[157];
      data_o_156_sv2v_reg <= data_i[156];
      data_o_155_sv2v_reg <= data_i[155];
      data_o_154_sv2v_reg <= data_i[154];
      data_o_153_sv2v_reg <= data_i[153];
      data_o_152_sv2v_reg <= data_i[152];
      data_o_151_sv2v_reg <= data_i[151];
      data_o_150_sv2v_reg <= data_i[150];
      data_o_149_sv2v_reg <= data_i[149];
      data_o_148_sv2v_reg <= data_i[148];
      data_o_147_sv2v_reg <= data_i[147];
      data_o_146_sv2v_reg <= data_i[146];
      data_o_145_sv2v_reg <= data_i[145];
      data_o_144_sv2v_reg <= data_i[144];
      data_o_143_sv2v_reg <= data_i[143];
      data_o_142_sv2v_reg <= data_i[142];
      data_o_141_sv2v_reg <= data_i[141];
      data_o_140_sv2v_reg <= data_i[140];
      data_o_139_sv2v_reg <= data_i[139];
      data_o_138_sv2v_reg <= data_i[138];
      data_o_137_sv2v_reg <= data_i[137];
      data_o_136_sv2v_reg <= data_i[136];
      data_o_135_sv2v_reg <= data_i[135];
      data_o_134_sv2v_reg <= data_i[134];
      data_o_133_sv2v_reg <= data_i[133];
      data_o_132_sv2v_reg <= data_i[132];
      data_o_131_sv2v_reg <= data_i[131];
      data_o_130_sv2v_reg <= data_i[130];
      data_o_129_sv2v_reg <= data_i[129];
      data_o_128_sv2v_reg <= data_i[128];
      data_o_127_sv2v_reg <= data_i[127];
      data_o_126_sv2v_reg <= data_i[126];
      data_o_125_sv2v_reg <= data_i[125];
      data_o_124_sv2v_reg <= data_i[124];
      data_o_123_sv2v_reg <= data_i[123];
      data_o_122_sv2v_reg <= data_i[122];
      data_o_121_sv2v_reg <= data_i[121];
      data_o_120_sv2v_reg <= data_i[120];
      data_o_119_sv2v_reg <= data_i[119];
      data_o_118_sv2v_reg <= data_i[118];
      data_o_117_sv2v_reg <= data_i[117];
      data_o_116_sv2v_reg <= data_i[116];
      data_o_115_sv2v_reg <= data_i[115];
      data_o_114_sv2v_reg <= data_i[114];
      data_o_113_sv2v_reg <= data_i[113];
      data_o_112_sv2v_reg <= data_i[112];
      data_o_111_sv2v_reg <= data_i[111];
      data_o_110_sv2v_reg <= data_i[110];
      data_o_109_sv2v_reg <= data_i[109];
      data_o_108_sv2v_reg <= data_i[108];
      data_o_107_sv2v_reg <= data_i[107];
      data_o_106_sv2v_reg <= data_i[106];
      data_o_105_sv2v_reg <= data_i[105];
      data_o_104_sv2v_reg <= data_i[104];
      data_o_103_sv2v_reg <= data_i[103];
      data_o_102_sv2v_reg <= data_i[102];
      data_o_101_sv2v_reg <= data_i[101];
      data_o_100_sv2v_reg <= data_i[100];
      data_o_99_sv2v_reg <= data_i[99];
      data_o_98_sv2v_reg <= data_i[98];
      data_o_97_sv2v_reg <= data_i[97];
      data_o_96_sv2v_reg <= data_i[96];
      data_o_95_sv2v_reg <= data_i[95];
      data_o_94_sv2v_reg <= data_i[94];
      data_o_93_sv2v_reg <= data_i[93];
      data_o_92_sv2v_reg <= data_i[92];
      data_o_91_sv2v_reg <= data_i[91];
      data_o_90_sv2v_reg <= data_i[90];
      data_o_89_sv2v_reg <= data_i[89];
      data_o_88_sv2v_reg <= data_i[88];
      data_o_87_sv2v_reg <= data_i[87];
      data_o_86_sv2v_reg <= data_i[86];
      data_o_85_sv2v_reg <= data_i[85];
      data_o_84_sv2v_reg <= data_i[84];
      data_o_83_sv2v_reg <= data_i[83];
      data_o_82_sv2v_reg <= data_i[82];
      data_o_81_sv2v_reg <= data_i[81];
      data_o_80_sv2v_reg <= data_i[80];
      data_o_79_sv2v_reg <= data_i[79];
      data_o_78_sv2v_reg <= data_i[78];
      data_o_77_sv2v_reg <= data_i[77];
      data_o_76_sv2v_reg <= data_i[76];
      data_o_75_sv2v_reg <= data_i[75];
      data_o_74_sv2v_reg <= data_i[74];
      data_o_73_sv2v_reg <= data_i[73];
      data_o_72_sv2v_reg <= data_i[72];
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_width_p190
(
  clk_i,
  data_i,
  data_o
);

  input [189:0] data_i;
  output [189:0] data_o;
  input clk_i;
  wire [189:0] data_o;
  reg data_o_189_sv2v_reg,data_o_188_sv2v_reg,data_o_187_sv2v_reg,data_o_186_sv2v_reg,
  data_o_185_sv2v_reg,data_o_184_sv2v_reg,data_o_183_sv2v_reg,data_o_182_sv2v_reg,
  data_o_181_sv2v_reg,data_o_180_sv2v_reg,data_o_179_sv2v_reg,data_o_178_sv2v_reg,
  data_o_177_sv2v_reg,data_o_176_sv2v_reg,data_o_175_sv2v_reg,data_o_174_sv2v_reg,
  data_o_173_sv2v_reg,data_o_172_sv2v_reg,data_o_171_sv2v_reg,data_o_170_sv2v_reg,
  data_o_169_sv2v_reg,data_o_168_sv2v_reg,data_o_167_sv2v_reg,data_o_166_sv2v_reg,
  data_o_165_sv2v_reg,data_o_164_sv2v_reg,data_o_163_sv2v_reg,data_o_162_sv2v_reg,
  data_o_161_sv2v_reg,data_o_160_sv2v_reg,data_o_159_sv2v_reg,data_o_158_sv2v_reg,
  data_o_157_sv2v_reg,data_o_156_sv2v_reg,data_o_155_sv2v_reg,data_o_154_sv2v_reg,
  data_o_153_sv2v_reg,data_o_152_sv2v_reg,data_o_151_sv2v_reg,data_o_150_sv2v_reg,
  data_o_149_sv2v_reg,data_o_148_sv2v_reg,data_o_147_sv2v_reg,data_o_146_sv2v_reg,
  data_o_145_sv2v_reg,data_o_144_sv2v_reg,data_o_143_sv2v_reg,data_o_142_sv2v_reg,
  data_o_141_sv2v_reg,data_o_140_sv2v_reg,data_o_139_sv2v_reg,data_o_138_sv2v_reg,
  data_o_137_sv2v_reg,data_o_136_sv2v_reg,data_o_135_sv2v_reg,data_o_134_sv2v_reg,
  data_o_133_sv2v_reg,data_o_132_sv2v_reg,data_o_131_sv2v_reg,data_o_130_sv2v_reg,
  data_o_129_sv2v_reg,data_o_128_sv2v_reg,data_o_127_sv2v_reg,data_o_126_sv2v_reg,
  data_o_125_sv2v_reg,data_o_124_sv2v_reg,data_o_123_sv2v_reg,data_o_122_sv2v_reg,
  data_o_121_sv2v_reg,data_o_120_sv2v_reg,data_o_119_sv2v_reg,data_o_118_sv2v_reg,
  data_o_117_sv2v_reg,data_o_116_sv2v_reg,data_o_115_sv2v_reg,data_o_114_sv2v_reg,
  data_o_113_sv2v_reg,data_o_112_sv2v_reg,data_o_111_sv2v_reg,data_o_110_sv2v_reg,
  data_o_109_sv2v_reg,data_o_108_sv2v_reg,data_o_107_sv2v_reg,data_o_106_sv2v_reg,
  data_o_105_sv2v_reg,data_o_104_sv2v_reg,data_o_103_sv2v_reg,data_o_102_sv2v_reg,
  data_o_101_sv2v_reg,data_o_100_sv2v_reg,data_o_99_sv2v_reg,data_o_98_sv2v_reg,
  data_o_97_sv2v_reg,data_o_96_sv2v_reg,data_o_95_sv2v_reg,data_o_94_sv2v_reg,
  data_o_93_sv2v_reg,data_o_92_sv2v_reg,data_o_91_sv2v_reg,data_o_90_sv2v_reg,
  data_o_89_sv2v_reg,data_o_88_sv2v_reg,data_o_87_sv2v_reg,data_o_86_sv2v_reg,
  data_o_85_sv2v_reg,data_o_84_sv2v_reg,data_o_83_sv2v_reg,data_o_82_sv2v_reg,
  data_o_81_sv2v_reg,data_o_80_sv2v_reg,data_o_79_sv2v_reg,data_o_78_sv2v_reg,data_o_77_sv2v_reg,
  data_o_76_sv2v_reg,data_o_75_sv2v_reg,data_o_74_sv2v_reg,data_o_73_sv2v_reg,
  data_o_72_sv2v_reg,data_o_71_sv2v_reg,data_o_70_sv2v_reg,data_o_69_sv2v_reg,
  data_o_68_sv2v_reg,data_o_67_sv2v_reg,data_o_66_sv2v_reg,data_o_65_sv2v_reg,
  data_o_64_sv2v_reg,data_o_63_sv2v_reg,data_o_62_sv2v_reg,data_o_61_sv2v_reg,data_o_60_sv2v_reg,
  data_o_59_sv2v_reg,data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,
  data_o_55_sv2v_reg,data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,
  data_o_51_sv2v_reg,data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,
  data_o_47_sv2v_reg,data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,
  data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,
  data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,
  data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,
  data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,
  data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,
  data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,
  data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[189] = data_o_189_sv2v_reg;
  assign data_o[188] = data_o_188_sv2v_reg;
  assign data_o[187] = data_o_187_sv2v_reg;
  assign data_o[186] = data_o_186_sv2v_reg;
  assign data_o[185] = data_o_185_sv2v_reg;
  assign data_o[184] = data_o_184_sv2v_reg;
  assign data_o[183] = data_o_183_sv2v_reg;
  assign data_o[182] = data_o_182_sv2v_reg;
  assign data_o[181] = data_o_181_sv2v_reg;
  assign data_o[180] = data_o_180_sv2v_reg;
  assign data_o[179] = data_o_179_sv2v_reg;
  assign data_o[178] = data_o_178_sv2v_reg;
  assign data_o[177] = data_o_177_sv2v_reg;
  assign data_o[176] = data_o_176_sv2v_reg;
  assign data_o[175] = data_o_175_sv2v_reg;
  assign data_o[174] = data_o_174_sv2v_reg;
  assign data_o[173] = data_o_173_sv2v_reg;
  assign data_o[172] = data_o_172_sv2v_reg;
  assign data_o[171] = data_o_171_sv2v_reg;
  assign data_o[170] = data_o_170_sv2v_reg;
  assign data_o[169] = data_o_169_sv2v_reg;
  assign data_o[168] = data_o_168_sv2v_reg;
  assign data_o[167] = data_o_167_sv2v_reg;
  assign data_o[166] = data_o_166_sv2v_reg;
  assign data_o[165] = data_o_165_sv2v_reg;
  assign data_o[164] = data_o_164_sv2v_reg;
  assign data_o[163] = data_o_163_sv2v_reg;
  assign data_o[162] = data_o_162_sv2v_reg;
  assign data_o[161] = data_o_161_sv2v_reg;
  assign data_o[160] = data_o_160_sv2v_reg;
  assign data_o[159] = data_o_159_sv2v_reg;
  assign data_o[158] = data_o_158_sv2v_reg;
  assign data_o[157] = data_o_157_sv2v_reg;
  assign data_o[156] = data_o_156_sv2v_reg;
  assign data_o[155] = data_o_155_sv2v_reg;
  assign data_o[154] = data_o_154_sv2v_reg;
  assign data_o[153] = data_o_153_sv2v_reg;
  assign data_o[152] = data_o_152_sv2v_reg;
  assign data_o[151] = data_o_151_sv2v_reg;
  assign data_o[150] = data_o_150_sv2v_reg;
  assign data_o[149] = data_o_149_sv2v_reg;
  assign data_o[148] = data_o_148_sv2v_reg;
  assign data_o[147] = data_o_147_sv2v_reg;
  assign data_o[146] = data_o_146_sv2v_reg;
  assign data_o[145] = data_o_145_sv2v_reg;
  assign data_o[144] = data_o_144_sv2v_reg;
  assign data_o[143] = data_o_143_sv2v_reg;
  assign data_o[142] = data_o_142_sv2v_reg;
  assign data_o[141] = data_o_141_sv2v_reg;
  assign data_o[140] = data_o_140_sv2v_reg;
  assign data_o[139] = data_o_139_sv2v_reg;
  assign data_o[138] = data_o_138_sv2v_reg;
  assign data_o[137] = data_o_137_sv2v_reg;
  assign data_o[136] = data_o_136_sv2v_reg;
  assign data_o[135] = data_o_135_sv2v_reg;
  assign data_o[134] = data_o_134_sv2v_reg;
  assign data_o[133] = data_o_133_sv2v_reg;
  assign data_o[132] = data_o_132_sv2v_reg;
  assign data_o[131] = data_o_131_sv2v_reg;
  assign data_o[130] = data_o_130_sv2v_reg;
  assign data_o[129] = data_o_129_sv2v_reg;
  assign data_o[128] = data_o_128_sv2v_reg;
  assign data_o[127] = data_o_127_sv2v_reg;
  assign data_o[126] = data_o_126_sv2v_reg;
  assign data_o[125] = data_o_125_sv2v_reg;
  assign data_o[124] = data_o_124_sv2v_reg;
  assign data_o[123] = data_o_123_sv2v_reg;
  assign data_o[122] = data_o_122_sv2v_reg;
  assign data_o[121] = data_o_121_sv2v_reg;
  assign data_o[120] = data_o_120_sv2v_reg;
  assign data_o[119] = data_o_119_sv2v_reg;
  assign data_o[118] = data_o_118_sv2v_reg;
  assign data_o[117] = data_o_117_sv2v_reg;
  assign data_o[116] = data_o_116_sv2v_reg;
  assign data_o[115] = data_o_115_sv2v_reg;
  assign data_o[114] = data_o_114_sv2v_reg;
  assign data_o[113] = data_o_113_sv2v_reg;
  assign data_o[112] = data_o_112_sv2v_reg;
  assign data_o[111] = data_o_111_sv2v_reg;
  assign data_o[110] = data_o_110_sv2v_reg;
  assign data_o[109] = data_o_109_sv2v_reg;
  assign data_o[108] = data_o_108_sv2v_reg;
  assign data_o[107] = data_o_107_sv2v_reg;
  assign data_o[106] = data_o_106_sv2v_reg;
  assign data_o[105] = data_o_105_sv2v_reg;
  assign data_o[104] = data_o_104_sv2v_reg;
  assign data_o[103] = data_o_103_sv2v_reg;
  assign data_o[102] = data_o_102_sv2v_reg;
  assign data_o[101] = data_o_101_sv2v_reg;
  assign data_o[100] = data_o_100_sv2v_reg;
  assign data_o[99] = data_o_99_sv2v_reg;
  assign data_o[98] = data_o_98_sv2v_reg;
  assign data_o[97] = data_o_97_sv2v_reg;
  assign data_o[96] = data_o_96_sv2v_reg;
  assign data_o[95] = data_o_95_sv2v_reg;
  assign data_o[94] = data_o_94_sv2v_reg;
  assign data_o[93] = data_o_93_sv2v_reg;
  assign data_o[92] = data_o_92_sv2v_reg;
  assign data_o[91] = data_o_91_sv2v_reg;
  assign data_o[90] = data_o_90_sv2v_reg;
  assign data_o[89] = data_o_89_sv2v_reg;
  assign data_o[88] = data_o_88_sv2v_reg;
  assign data_o[87] = data_o_87_sv2v_reg;
  assign data_o[86] = data_o_86_sv2v_reg;
  assign data_o[85] = data_o_85_sv2v_reg;
  assign data_o[84] = data_o_84_sv2v_reg;
  assign data_o[83] = data_o_83_sv2v_reg;
  assign data_o[82] = data_o_82_sv2v_reg;
  assign data_o[81] = data_o_81_sv2v_reg;
  assign data_o[80] = data_o_80_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_189_sv2v_reg <= data_i[189];
      data_o_188_sv2v_reg <= data_i[188];
      data_o_187_sv2v_reg <= data_i[187];
      data_o_186_sv2v_reg <= data_i[186];
      data_o_185_sv2v_reg <= data_i[185];
      data_o_184_sv2v_reg <= data_i[184];
      data_o_183_sv2v_reg <= data_i[183];
      data_o_182_sv2v_reg <= data_i[182];
      data_o_181_sv2v_reg <= data_i[181];
      data_o_180_sv2v_reg <= data_i[180];
      data_o_179_sv2v_reg <= data_i[179];
      data_o_178_sv2v_reg <= data_i[178];
      data_o_177_sv2v_reg <= data_i[177];
      data_o_176_sv2v_reg <= data_i[176];
      data_o_175_sv2v_reg <= data_i[175];
      data_o_174_sv2v_reg <= data_i[174];
      data_o_173_sv2v_reg <= data_i[173];
      data_o_172_sv2v_reg <= data_i[172];
      data_o_171_sv2v_reg <= data_i[171];
      data_o_170_sv2v_reg <= data_i[170];
      data_o_169_sv2v_reg <= data_i[169];
      data_o_168_sv2v_reg <= data_i[168];
      data_o_167_sv2v_reg <= data_i[167];
      data_o_166_sv2v_reg <= data_i[166];
      data_o_165_sv2v_reg <= data_i[165];
      data_o_164_sv2v_reg <= data_i[164];
      data_o_163_sv2v_reg <= data_i[163];
      data_o_162_sv2v_reg <= data_i[162];
      data_o_161_sv2v_reg <= data_i[161];
      data_o_160_sv2v_reg <= data_i[160];
      data_o_159_sv2v_reg <= data_i[159];
      data_o_158_sv2v_reg <= data_i[158];
      data_o_157_sv2v_reg <= data_i[157];
      data_o_156_sv2v_reg <= data_i[156];
      data_o_155_sv2v_reg <= data_i[155];
      data_o_154_sv2v_reg <= data_i[154];
      data_o_153_sv2v_reg <= data_i[153];
      data_o_152_sv2v_reg <= data_i[152];
      data_o_151_sv2v_reg <= data_i[151];
      data_o_150_sv2v_reg <= data_i[150];
      data_o_149_sv2v_reg <= data_i[149];
      data_o_148_sv2v_reg <= data_i[148];
      data_o_147_sv2v_reg <= data_i[147];
      data_o_146_sv2v_reg <= data_i[146];
      data_o_145_sv2v_reg <= data_i[145];
      data_o_144_sv2v_reg <= data_i[144];
      data_o_143_sv2v_reg <= data_i[143];
      data_o_142_sv2v_reg <= data_i[142];
      data_o_141_sv2v_reg <= data_i[141];
      data_o_140_sv2v_reg <= data_i[140];
      data_o_139_sv2v_reg <= data_i[139];
      data_o_138_sv2v_reg <= data_i[138];
      data_o_137_sv2v_reg <= data_i[137];
      data_o_136_sv2v_reg <= data_i[136];
      data_o_135_sv2v_reg <= data_i[135];
      data_o_134_sv2v_reg <= data_i[134];
      data_o_133_sv2v_reg <= data_i[133];
      data_o_132_sv2v_reg <= data_i[132];
      data_o_131_sv2v_reg <= data_i[131];
      data_o_130_sv2v_reg <= data_i[130];
      data_o_129_sv2v_reg <= data_i[129];
      data_o_128_sv2v_reg <= data_i[128];
      data_o_127_sv2v_reg <= data_i[127];
      data_o_126_sv2v_reg <= data_i[126];
      data_o_125_sv2v_reg <= data_i[125];
      data_o_124_sv2v_reg <= data_i[124];
      data_o_123_sv2v_reg <= data_i[123];
      data_o_122_sv2v_reg <= data_i[122];
      data_o_121_sv2v_reg <= data_i[121];
      data_o_120_sv2v_reg <= data_i[120];
      data_o_119_sv2v_reg <= data_i[119];
      data_o_118_sv2v_reg <= data_i[118];
      data_o_117_sv2v_reg <= data_i[117];
      data_o_116_sv2v_reg <= data_i[116];
      data_o_115_sv2v_reg <= data_i[115];
      data_o_114_sv2v_reg <= data_i[114];
      data_o_113_sv2v_reg <= data_i[113];
      data_o_112_sv2v_reg <= data_i[112];
      data_o_111_sv2v_reg <= data_i[111];
      data_o_110_sv2v_reg <= data_i[110];
      data_o_109_sv2v_reg <= data_i[109];
      data_o_108_sv2v_reg <= data_i[108];
      data_o_107_sv2v_reg <= data_i[107];
      data_o_106_sv2v_reg <= data_i[106];
      data_o_105_sv2v_reg <= data_i[105];
      data_o_104_sv2v_reg <= data_i[104];
      data_o_103_sv2v_reg <= data_i[103];
      data_o_102_sv2v_reg <= data_i[102];
      data_o_101_sv2v_reg <= data_i[101];
      data_o_100_sv2v_reg <= data_i[100];
      data_o_99_sv2v_reg <= data_i[99];
      data_o_98_sv2v_reg <= data_i[98];
      data_o_97_sv2v_reg <= data_i[97];
      data_o_96_sv2v_reg <= data_i[96];
      data_o_95_sv2v_reg <= data_i[95];
      data_o_94_sv2v_reg <= data_i[94];
      data_o_93_sv2v_reg <= data_i[93];
      data_o_92_sv2v_reg <= data_i[92];
      data_o_91_sv2v_reg <= data_i[91];
      data_o_90_sv2v_reg <= data_i[90];
      data_o_89_sv2v_reg <= data_i[89];
      data_o_88_sv2v_reg <= data_i[88];
      data_o_87_sv2v_reg <= data_i[87];
      data_o_86_sv2v_reg <= data_i[86];
      data_o_85_sv2v_reg <= data_i[85];
      data_o_84_sv2v_reg <= data_i[84];
      data_o_83_sv2v_reg <= data_i[83];
      data_o_82_sv2v_reg <= data_i[82];
      data_o_81_sv2v_reg <= data_i[81];
      data_o_80_sv2v_reg <= data_i[80];
      data_o_79_sv2v_reg <= data_i[79];
      data_o_78_sv2v_reg <= data_i[78];
      data_o_77_sv2v_reg <= data_i[77];
      data_o_76_sv2v_reg <= data_i[76];
      data_o_75_sv2v_reg <= data_i[75];
      data_o_74_sv2v_reg <= data_i[74];
      data_o_73_sv2v_reg <= data_i[73];
      data_o_72_sv2v_reg <= data_i[72];
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bp_be_calculator_top_00
(
  clk_i,
  reset_i,
  cfg_bus_i,
  dispatch_pkt_i,
  idiv_busy_o,
  fdiv_busy_o,
  mem_busy_o,
  mem_ordered_o,
  decode_info_o,
  trans_info_o,
  cmd_full_n_i,
  commit_pkt_o,
  br_pkt_o,
  iwb_pkt_o,
  fwb_pkt_o,
  late_wb_pkt_o,
  late_wb_v_o,
  late_wb_force_o,
  late_wb_yumi_i,
  debug_irq_i,
  timer_irq_i,
  software_irq_i,
  m_external_irq_i,
  s_external_irq_i,
  irq_waiting_o,
  irq_pending_o,
  cache_req_o,
  cache_req_v_o,
  cache_req_yumi_i,
  cache_req_lock_i,
  cache_req_metadata_o,
  cache_req_metadata_v_o,
  cache_req_id_i,
  cache_req_critical_i,
  cache_req_last_i,
  cache_req_credits_full_i,
  cache_req_credits_empty_i,
  data_mem_pkt_v_i,
  data_mem_pkt_i,
  data_mem_pkt_yumi_o,
  data_mem_o,
  tag_mem_pkt_v_i,
  tag_mem_pkt_i,
  tag_mem_pkt_yumi_o,
  tag_mem_o,
  stat_mem_pkt_v_i,
  stat_mem_pkt_i,
  stat_mem_pkt_yumi_o,
  stat_mem_o
);

  input [60:0] cfg_bus_i;
  input [365:0] dispatch_pkt_i;
  output [12:0] decode_info_o;
  output [32:0] trans_info_o;
  output [213:0] commit_pkt_o;
  output [42:0] br_pkt_o;
  output [78:0] iwb_pkt_o;
  output [78:0] fwb_pkt_o;
  output [78:0] late_wb_pkt_o;
  output [116:0] cache_req_o;
  output [3:0] cache_req_metadata_o;
  input [0:0] cache_req_id_i;
  input [142:0] data_mem_pkt_i;
  output [511:0] data_mem_o;
  input [34:0] tag_mem_pkt_i;
  output [22:0] tag_mem_o;
  input [10:0] stat_mem_pkt_i;
  output [14:0] stat_mem_o;
  input clk_i;
  input reset_i;
  input cmd_full_n_i;
  input late_wb_yumi_i;
  input debug_irq_i;
  input timer_irq_i;
  input software_irq_i;
  input m_external_irq_i;
  input s_external_irq_i;
  input cache_req_yumi_i;
  input cache_req_lock_i;
  input cache_req_critical_i;
  input cache_req_last_i;
  input cache_req_credits_full_i;
  input cache_req_credits_empty_i;
  input data_mem_pkt_v_i;
  input tag_mem_pkt_v_i;
  input stat_mem_pkt_v_i;
  output idiv_busy_o;
  output fdiv_busy_o;
  output mem_busy_o;
  output mem_ordered_o;
  output late_wb_v_o;
  output late_wb_force_o;
  output irq_waiting_o;
  output irq_pending_o;
  output cache_req_v_o;
  output cache_req_metadata_v_o;
  output data_mem_pkt_yumi_o;
  output tag_mem_pkt_yumi_o;
  output stat_mem_pkt_yumi_o;
  wire [12:0] decode_info_o;
  wire [32:0] trans_info_o;
  wire [213:0] commit_pkt_o;
  wire [42:0] br_pkt_o;
  wire [78:0] iwb_pkt_o,fwb_pkt_o,late_wb_pkt_o,pipe_mem_late_wb_pkt,pipe_long_iwb_pkt,
  pipe_long_fwb_pkt;
  wire [116:0] cache_req_o;
  wire [3:0] cache_req_metadata_o;
  wire [511:0] data_mem_o;
  wire [22:0] tag_mem_o;
  wire [14:0] stat_mem_o,match_rs;
  wire idiv_busy_o,fdiv_busy_o,mem_busy_o,mem_ordered_o,late_wb_v_o,late_wb_force_o,
  irq_waiting_o,irq_pending_o,cache_req_v_o,cache_req_metadata_v_o,
  data_mem_pkt_yumi_o,tag_mem_pkt_yumi_o,stat_mem_pkt_yumi_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,
  N12,N13,N14,N15,N16,N17,N18,N19,N20,comp_stage_r_2__ird_w_v_,
  comp_stage_r_2__frd_w_v_,comp_stage_r_2__rd_data__65_,comp_stage_r_2__rd_data__64_,
  comp_stage_r_2__rd_data__63_,comp_stage_r_2__rd_data__62_,comp_stage_r_2__rd_data__61_,
  comp_stage_r_2__rd_data__60_,comp_stage_r_2__rd_data__59_,comp_stage_r_2__rd_data__58_,
  comp_stage_r_2__rd_data__57_,comp_stage_r_2__rd_data__56_,
  comp_stage_r_2__rd_data__55_,comp_stage_r_2__rd_data__54_,comp_stage_r_2__rd_data__53_,
  comp_stage_r_2__rd_data__52_,comp_stage_r_2__rd_data__51_,comp_stage_r_2__rd_data__50_,
  comp_stage_r_2__rd_data__49_,comp_stage_r_2__rd_data__48_,comp_stage_r_2__rd_data__47_,
  comp_stage_r_2__rd_data__46_,comp_stage_r_2__rd_data__45_,
  comp_stage_r_2__rd_data__44_,comp_stage_r_2__rd_data__43_,comp_stage_r_2__rd_data__42_,
  comp_stage_r_2__rd_data__41_,comp_stage_r_2__rd_data__40_,comp_stage_r_2__rd_data__39_,
  comp_stage_r_2__rd_data__38_,comp_stage_r_2__rd_data__37_,comp_stage_r_2__rd_data__36_,
  comp_stage_r_2__rd_data__35_,comp_stage_r_2__rd_data__34_,
  comp_stage_r_2__rd_data__33_,comp_stage_r_2__rd_data__32_,comp_stage_r_2__rd_data__31_,
  comp_stage_r_2__rd_data__30_,comp_stage_r_2__rd_data__29_,comp_stage_r_2__rd_data__28_,
  comp_stage_r_2__rd_data__27_,comp_stage_r_2__rd_data__26_,comp_stage_r_2__rd_data__25_,
  comp_stage_r_2__rd_data__24_,comp_stage_r_2__rd_data__23_,
  comp_stage_r_2__rd_data__22_,comp_stage_r_2__rd_data__21_,comp_stage_r_2__rd_data__20_,
  comp_stage_r_2__rd_data__19_,comp_stage_r_2__rd_data__18_,comp_stage_r_2__rd_data__17_,
  comp_stage_r_2__rd_data__16_,comp_stage_r_2__rd_data__15_,comp_stage_r_2__rd_data__14_,
  comp_stage_r_2__rd_data__13_,comp_stage_r_2__rd_data__12_,comp_stage_r_2__rd_data__11_,
  comp_stage_r_2__rd_data__10_,comp_stage_r_2__rd_data__9_,
  comp_stage_r_2__rd_data__8_,comp_stage_r_2__rd_data__7_,comp_stage_r_2__rd_data__6_,
  comp_stage_r_2__rd_data__5_,comp_stage_r_2__rd_data__4_,comp_stage_r_2__rd_data__3_,
  comp_stage_r_2__rd_data__2_,comp_stage_r_2__rd_data__1_,comp_stage_r_2__rd_data__0_,
  comp_stage_r_2__fflags__nv_,comp_stage_r_2__fflags__dz_,comp_stage_r_2__fflags__of_,
  comp_stage_r_2__fflags__uf_,comp_stage_r_2__fflags__nx_,comp_stage_r_1__ird_w_v_,
  comp_stage_r_1__frd_w_v_,comp_stage_r_1__rd_data__65_,comp_stage_r_1__rd_data__64_,
  comp_stage_r_1__rd_data__63_,comp_stage_r_1__rd_data__62_,
  comp_stage_r_1__rd_data__61_,comp_stage_r_1__rd_data__60_,comp_stage_r_1__rd_data__59_,
  comp_stage_r_1__rd_data__58_,comp_stage_r_1__rd_data__57_,comp_stage_r_1__rd_data__56_,
  comp_stage_r_1__rd_data__55_,comp_stage_r_1__rd_data__54_,comp_stage_r_1__rd_data__53_,
  comp_stage_r_1__rd_data__52_,comp_stage_r_1__rd_data__51_,
  comp_stage_r_1__rd_data__50_,comp_stage_r_1__rd_data__49_,comp_stage_r_1__rd_data__48_,
  comp_stage_r_1__rd_data__47_,comp_stage_r_1__rd_data__46_,comp_stage_r_1__rd_data__45_,
  comp_stage_r_1__rd_data__44_,comp_stage_r_1__rd_data__43_,comp_stage_r_1__rd_data__42_,
  comp_stage_r_1__rd_data__41_,comp_stage_r_1__rd_data__40_,
  comp_stage_r_1__rd_data__39_,comp_stage_r_1__rd_data__38_,comp_stage_r_1__rd_data__37_,
  comp_stage_r_1__rd_data__36_,comp_stage_r_1__rd_data__35_,comp_stage_r_1__rd_data__34_,
  comp_stage_r_1__rd_data__33_,comp_stage_r_1__rd_data__32_,comp_stage_r_1__rd_data__31_,
  comp_stage_r_1__rd_data__30_,comp_stage_r_1__rd_data__29_,
  comp_stage_r_1__rd_data__28_,comp_stage_r_1__rd_data__27_,comp_stage_r_1__rd_data__26_,
  comp_stage_r_1__rd_data__25_,comp_stage_r_1__rd_data__24_,comp_stage_r_1__rd_data__23_,
  comp_stage_r_1__rd_data__22_,comp_stage_r_1__rd_data__21_,comp_stage_r_1__rd_data__20_,
  comp_stage_r_1__rd_data__19_,comp_stage_r_1__rd_data__18_,comp_stage_r_1__rd_data__17_,
  comp_stage_r_1__rd_data__16_,comp_stage_r_1__rd_data__15_,
  comp_stage_r_1__rd_data__14_,comp_stage_r_1__rd_data__13_,comp_stage_r_1__rd_data__12_,
  comp_stage_r_1__rd_data__11_,comp_stage_r_1__rd_data__10_,comp_stage_r_1__rd_data__9_,
  comp_stage_r_1__rd_data__8_,comp_stage_r_1__rd_data__7_,comp_stage_r_1__rd_data__6_,
  comp_stage_r_1__rd_data__5_,comp_stage_r_1__rd_data__4_,comp_stage_r_1__rd_data__3_,
  comp_stage_r_1__rd_data__2_,comp_stage_r_1__rd_data__1_,
  comp_stage_r_1__rd_data__0_,comp_stage_r_1__fflags__nv_,comp_stage_r_1__fflags__dz_,
  comp_stage_r_1__fflags__of_,comp_stage_r_1__fflags__uf_,comp_stage_r_1__fflags__nx_,
  comp_stage_r_0__ird_w_v_,comp_stage_r_0__frd_w_v_,comp_stage_r_0__rd_data__65_,
  comp_stage_r_0__rd_data__64_,comp_stage_r_0__rd_data__63_,comp_stage_r_0__rd_data__62_,
  comp_stage_r_0__rd_data__61_,comp_stage_r_0__rd_data__60_,comp_stage_r_0__rd_data__59_,
  comp_stage_r_0__rd_data__58_,comp_stage_r_0__rd_data__57_,
  comp_stage_r_0__rd_data__56_,comp_stage_r_0__rd_data__55_,comp_stage_r_0__rd_data__54_,
  comp_stage_r_0__rd_data__53_,comp_stage_r_0__rd_data__52_,comp_stage_r_0__rd_data__51_,
  comp_stage_r_0__rd_data__50_,comp_stage_r_0__rd_data__49_,comp_stage_r_0__rd_data__48_,
  comp_stage_r_0__rd_data__47_,comp_stage_r_0__rd_data__46_,
  comp_stage_r_0__rd_data__45_,comp_stage_r_0__rd_data__44_,comp_stage_r_0__rd_data__43_,
  comp_stage_r_0__rd_data__42_,comp_stage_r_0__rd_data__41_,comp_stage_r_0__rd_data__40_,
  comp_stage_r_0__rd_data__39_,comp_stage_r_0__rd_data__38_,comp_stage_r_0__rd_data__37_,
  comp_stage_r_0__rd_data__36_,comp_stage_r_0__rd_data__35_,
  comp_stage_r_0__rd_data__34_,comp_stage_r_0__rd_data__33_,comp_stage_r_0__rd_data__32_,
  comp_stage_r_0__rd_data__31_,comp_stage_r_0__rd_data__30_,comp_stage_r_0__rd_data__29_,
  comp_stage_r_0__rd_data__28_,comp_stage_r_0__rd_data__27_,comp_stage_r_0__rd_data__26_,
  comp_stage_r_0__rd_data__25_,comp_stage_r_0__rd_data__24_,comp_stage_r_0__rd_data__23_,
  comp_stage_r_0__rd_data__22_,comp_stage_r_0__rd_data__21_,
  comp_stage_r_0__rd_data__20_,comp_stage_r_0__rd_data__19_,comp_stage_r_0__rd_data__18_,
  comp_stage_r_0__rd_data__17_,comp_stage_r_0__rd_data__16_,comp_stage_r_0__rd_data__15_,
  comp_stage_r_0__rd_data__14_,comp_stage_r_0__rd_data__13_,comp_stage_r_0__rd_data__12_,
  comp_stage_r_0__rd_data__11_,comp_stage_r_0__rd_data__10_,
  comp_stage_r_0__rd_data__9_,comp_stage_r_0__rd_data__8_,comp_stage_r_0__rd_data__7_,
  comp_stage_r_0__rd_data__6_,comp_stage_r_0__rd_data__5_,comp_stage_r_0__rd_data__4_,
  comp_stage_r_0__rd_data__3_,comp_stage_r_0__rd_data__2_,comp_stage_r_0__rd_data__1_,
  comp_stage_r_0__rd_data__0_,comp_stage_r_0__fflags__nv_,comp_stage_r_0__fflags__dz_,
  comp_stage_r_0__fflags__of_,comp_stage_r_0__fflags__uf_,comp_stage_r_0__fflags__nx_,
  N21,N22,N23,N24,N25,comp_stage_n_4__ird_w_v_,comp_stage_n_4__frd_w_v_,
  comp_stage_n_4__fflags__nv_,comp_stage_n_4__fflags__dz_,comp_stage_n_4__fflags__of_,
  comp_stage_n_4__fflags__uf_,comp_stage_n_4__fflags__nx_,comp_stage_n_3__ird_w_v_,
  comp_stage_n_3__frd_w_v_,comp_stage_n_3__ptw_w_v_,comp_stage_n_3__rd_addr__4_,
  comp_stage_n_3__rd_addr__3_,comp_stage_n_3__rd_addr__2_,comp_stage_n_3__rd_addr__1_,
  comp_stage_n_3__rd_addr__0_,comp_stage_n_3__fflags__nv_,comp_stage_n_3__fflags__dz_,
  comp_stage_n_3__fflags__of_,comp_stage_n_3__fflags__uf_,
  comp_stage_n_3__fflags__nx_,comp_stage_n_2__ird_w_v_,comp_stage_n_2__frd_w_v_,comp_stage_n_2__ptw_w_v_,
  comp_stage_n_2__rd_addr__4_,comp_stage_n_2__rd_addr__3_,
  comp_stage_n_2__rd_addr__2_,comp_stage_n_2__rd_addr__1_,comp_stage_n_2__rd_addr__0_,
  comp_stage_n_2__fflags__nv_,comp_stage_n_2__fflags__dz_,comp_stage_n_2__fflags__of_,
  comp_stage_n_2__fflags__uf_,comp_stage_n_2__fflags__nx_,comp_stage_n_1__ird_w_v_,
  comp_stage_n_1__frd_w_v_,comp_stage_n_1__ptw_w_v_,comp_stage_n_1__rd_addr__4_,
  comp_stage_n_1__rd_addr__3_,comp_stage_n_1__rd_addr__2_,comp_stage_n_1__rd_addr__1_,
  comp_stage_n_1__rd_addr__0_,comp_stage_n_1__fflags__nv_,comp_stage_n_1__fflags__dz_,
  comp_stage_n_1__fflags__of_,comp_stage_n_1__fflags__uf_,comp_stage_n_1__fflags__nx_,
  comp_stage_n_0__ird_w_v_,comp_stage_n_0__frd_w_v_,comp_stage_n_0__rd_data__65_,
  comp_stage_n_0__rd_data__64_,comp_stage_n_0__rd_data__63_,comp_stage_n_0__rd_data__62_,
  comp_stage_n_0__rd_data__61_,comp_stage_n_0__rd_data__60_,
  comp_stage_n_0__rd_data__59_,comp_stage_n_0__rd_data__58_,comp_stage_n_0__rd_data__57_,
  comp_stage_n_0__rd_data__56_,comp_stage_n_0__rd_data__55_,comp_stage_n_0__rd_data__54_,
  comp_stage_n_0__rd_data__53_,comp_stage_n_0__rd_data__52_,comp_stage_n_0__rd_data__51_,
  comp_stage_n_0__rd_data__50_,comp_stage_n_0__rd_data__49_,
  comp_stage_n_0__rd_data__48_,comp_stage_n_0__rd_data__47_,comp_stage_n_0__rd_data__46_,
  comp_stage_n_0__rd_data__45_,comp_stage_n_0__rd_data__44_,comp_stage_n_0__rd_data__43_,
  comp_stage_n_0__rd_data__42_,comp_stage_n_0__rd_data__41_,comp_stage_n_0__rd_data__40_,
  comp_stage_n_0__rd_data__39_,comp_stage_n_0__rd_data__38_,
  comp_stage_n_0__rd_data__37_,comp_stage_n_0__rd_data__36_,comp_stage_n_0__rd_data__35_,
  comp_stage_n_0__rd_data__34_,comp_stage_n_0__rd_data__33_,comp_stage_n_0__rd_data__32_,
  comp_stage_n_0__rd_data__31_,comp_stage_n_0__rd_data__30_,comp_stage_n_0__rd_data__29_,
  comp_stage_n_0__rd_data__28_,comp_stage_n_0__rd_data__27_,
  comp_stage_n_0__rd_data__26_,comp_stage_n_0__rd_data__25_,comp_stage_n_0__rd_data__24_,
  comp_stage_n_0__rd_data__23_,comp_stage_n_0__rd_data__22_,comp_stage_n_0__rd_data__21_,
  comp_stage_n_0__rd_data__20_,comp_stage_n_0__rd_data__19_,comp_stage_n_0__rd_data__18_,
  comp_stage_n_0__rd_data__17_,comp_stage_n_0__rd_data__16_,
  comp_stage_n_0__rd_data__15_,comp_stage_n_0__rd_data__14_,comp_stage_n_0__rd_data__13_,
  comp_stage_n_0__rd_data__12_,comp_stage_n_0__rd_data__11_,comp_stage_n_0__rd_data__10_,
  comp_stage_n_0__rd_data__9_,comp_stage_n_0__rd_data__8_,comp_stage_n_0__rd_data__7_,
  comp_stage_n_0__rd_data__6_,comp_stage_n_0__rd_data__5_,comp_stage_n_0__rd_data__4_,
  comp_stage_n_0__rd_data__3_,comp_stage_n_0__rd_data__2_,comp_stage_n_0__rd_data__1_,
  comp_stage_n_0__rd_data__0_,comp_stage_n_0__fflags__nv_,
  comp_stage_n_0__fflags__dz_,comp_stage_n_0__fflags__of_,comp_stage_n_0__fflags__uf_,
  comp_stage_n_0__fflags__nx_,forward_data_3__65_,forward_data_3__64_,forward_data_3__63_,
  forward_data_3__62_,forward_data_3__61_,forward_data_3__60_,forward_data_3__59_,
  forward_data_3__58_,forward_data_3__57_,forward_data_3__56_,forward_data_3__55_,
  forward_data_3__54_,forward_data_3__53_,forward_data_3__52_,forward_data_3__51_,
  forward_data_3__50_,forward_data_3__49_,forward_data_3__48_,forward_data_3__47_,
  forward_data_3__46_,forward_data_3__45_,forward_data_3__44_,forward_data_3__43_,
  forward_data_3__42_,forward_data_3__41_,forward_data_3__40_,forward_data_3__39_,
  forward_data_3__38_,forward_data_3__37_,forward_data_3__36_,forward_data_3__35_,
  forward_data_3__34_,forward_data_3__33_,forward_data_3__32_,forward_data_3__31_,
  forward_data_3__30_,forward_data_3__29_,forward_data_3__28_,forward_data_3__27_,
  forward_data_3__26_,forward_data_3__25_,forward_data_3__24_,forward_data_3__23_,
  forward_data_3__22_,forward_data_3__21_,forward_data_3__20_,forward_data_3__19_,
  forward_data_3__18_,forward_data_3__17_,forward_data_3__16_,forward_data_3__15_,
  forward_data_3__14_,forward_data_3__13_,forward_data_3__12_,forward_data_3__11_,
  forward_data_3__10_,forward_data_3__9_,forward_data_3__8_,forward_data_3__7_,
  forward_data_3__6_,forward_data_3__5_,forward_data_3__4_,forward_data_3__3_,forward_data_3__2_,
  forward_data_3__1_,forward_data_3__0_,forward_data_2__65_,forward_data_2__64_,
  forward_data_2__63_,forward_data_2__62_,forward_data_2__61_,forward_data_2__60_,
  forward_data_2__59_,forward_data_2__58_,forward_data_2__57_,forward_data_2__56_,
  forward_data_2__55_,forward_data_2__54_,forward_data_2__53_,forward_data_2__52_,
  forward_data_2__51_,forward_data_2__50_,forward_data_2__49_,forward_data_2__48_,
  forward_data_2__47_,forward_data_2__46_,forward_data_2__45_,forward_data_2__44_,
  forward_data_2__43_,forward_data_2__42_,forward_data_2__41_,forward_data_2__40_,
  forward_data_2__39_,forward_data_2__38_,forward_data_2__37_,forward_data_2__36_,
  forward_data_2__35_,forward_data_2__34_,forward_data_2__33_,forward_data_2__32_,
  forward_data_2__31_,forward_data_2__30_,forward_data_2__29_,forward_data_2__28_,
  forward_data_2__27_,forward_data_2__26_,forward_data_2__25_,forward_data_2__24_,
  forward_data_2__23_,forward_data_2__22_,forward_data_2__21_,forward_data_2__20_,
  forward_data_2__19_,forward_data_2__18_,forward_data_2__17_,forward_data_2__16_,
  forward_data_2__15_,forward_data_2__14_,forward_data_2__13_,forward_data_2__12_,
  forward_data_2__11_,forward_data_2__10_,forward_data_2__9_,forward_data_2__8_,
  forward_data_2__7_,forward_data_2__6_,forward_data_2__5_,forward_data_2__4_,
  forward_data_2__3_,forward_data_2__2_,forward_data_2__1_,forward_data_2__0_,
  forward_data_1__65_,forward_data_1__64_,forward_data_1__63_,forward_data_1__62_,
  forward_data_1__61_,forward_data_1__60_,forward_data_1__59_,forward_data_1__58_,
  forward_data_1__57_,forward_data_1__56_,forward_data_1__55_,forward_data_1__54_,
  forward_data_1__53_,forward_data_1__52_,forward_data_1__51_,forward_data_1__50_,
  forward_data_1__49_,forward_data_1__48_,forward_data_1__47_,forward_data_1__46_,
  forward_data_1__45_,forward_data_1__44_,forward_data_1__43_,forward_data_1__42_,
  forward_data_1__41_,forward_data_1__40_,forward_data_1__39_,forward_data_1__38_,
  forward_data_1__37_,forward_data_1__36_,forward_data_1__35_,forward_data_1__34_,
  forward_data_1__33_,forward_data_1__32_,forward_data_1__31_,forward_data_1__30_,
  forward_data_1__29_,forward_data_1__28_,forward_data_1__27_,forward_data_1__26_,
  forward_data_1__25_,forward_data_1__24_,forward_data_1__23_,forward_data_1__22_,
  forward_data_1__21_,forward_data_1__20_,forward_data_1__19_,forward_data_1__18_,
  forward_data_1__17_,forward_data_1__16_,forward_data_1__15_,forward_data_1__14_,
  forward_data_1__13_,forward_data_1__12_,forward_data_1__11_,forward_data_1__10_,
  forward_data_1__9_,forward_data_1__8_,forward_data_1__7_,forward_data_1__6_,
  forward_data_1__5_,forward_data_1__4_,forward_data_1__3_,forward_data_1__2_,forward_data_1__1_,
  forward_data_1__0_,forward_data_0__65_,forward_data_0__64_,forward_data_0__63_,
  forward_data_0__62_,forward_data_0__61_,forward_data_0__60_,forward_data_0__59_,
  forward_data_0__58_,forward_data_0__57_,forward_data_0__56_,forward_data_0__55_,
  forward_data_0__54_,forward_data_0__53_,forward_data_0__52_,forward_data_0__51_,
  forward_data_0__50_,forward_data_0__49_,forward_data_0__48_,forward_data_0__47_,
  forward_data_0__46_,forward_data_0__45_,forward_data_0__44_,forward_data_0__43_,
  forward_data_0__42_,forward_data_0__41_,forward_data_0__40_,forward_data_0__39_,
  forward_data_0__38_,forward_data_0__37_,forward_data_0__36_,forward_data_0__35_,
  forward_data_0__34_,forward_data_0__33_,forward_data_0__32_,forward_data_0__31_,
  forward_data_0__30_,forward_data_0__29_,forward_data_0__28_,forward_data_0__27_,
  forward_data_0__26_,forward_data_0__25_,forward_data_0__24_,forward_data_0__23_,
  forward_data_0__22_,forward_data_0__21_,forward_data_0__20_,forward_data_0__19_,
  forward_data_0__18_,forward_data_0__17_,forward_data_0__16_,forward_data_0__15_,
  forward_data_0__14_,forward_data_0__13_,forward_data_0__12_,forward_data_0__11_,
  forward_data_0__10_,forward_data_0__9_,forward_data_0__8_,forward_data_0__7_,
  forward_data_0__6_,forward_data_0__5_,forward_data_0__4_,forward_data_0__3_,
  forward_data_0__2_,forward_data_0__1_,forward_data_0__0_,N26,N27,N28,N29,N30,N31,N32,N33,
  N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,pipe_sys_illegal_instr_lo,
  pipe_sys_data_v_lo,exc_stage_r_2__v_,exc_stage_r_1__v_,exc_stage_r_1__queue_v_,
  exc_stage_r_1__exc__instr_misaligned_,exc_stage_r_1__exc__dcache_replay_,
  exc_stage_r_1__exc__cmd_full_,exc_stage_r_1__exc__mispredict_,exc_stage_r_1__spec__dcache_miss_,
  exc_stage_r_0__v_,exc_stage_r_0__queue_v_,exc_stage_r_0__exc__store_page_fault_,
  exc_stage_r_0__exc__load_page_fault_,exc_stage_r_0__exc__store_access_fault_,
  exc_stage_r_0__exc__store_misaligned_,exc_stage_r_0__exc__load_access_fault_,
  exc_stage_r_0__exc__load_misaligned_,exc_stage_r_0__exc__illegal_instr_,
  exc_stage_r_0__exc__instr_misaligned_,exc_stage_r_0__exc__dtlb_load_miss_,
  exc_stage_r_0__exc__dtlb_store_miss_,_12_net_,pipe_int_early_data_v_lo,pipe_int_early_branch_lo,
  pipe_int_early_btaken_lo,pipe_int_early_instr_misaligned_lo,
  \catchup.catchup_reservation_n_isrc1__64_ ,\catchup.catchup_reservation_n_isrc1__63_ ,
  \catchup.catchup_reservation_n_isrc1__62_ ,\catchup.catchup_reservation_n_isrc1__61_ ,
  \catchup.catchup_reservation_n_isrc1__60_ ,\catchup.catchup_reservation_n_isrc1__59_ ,
  \catchup.catchup_reservation_n_isrc1__58_ ,\catchup.catchup_reservation_n_isrc1__57_ ,
  \catchup.catchup_reservation_n_isrc1__56_ ,\catchup.catchup_reservation_n_isrc1__55_ ,
  \catchup.catchup_reservation_n_isrc1__54_ ,
  \catchup.catchup_reservation_n_isrc1__53_ ,\catchup.catchup_reservation_n_isrc1__52_ ,
  \catchup.catchup_reservation_n_isrc1__51_ ,\catchup.catchup_reservation_n_isrc1__50_ ,
  \catchup.catchup_reservation_n_isrc1__49_ ,\catchup.catchup_reservation_n_isrc1__48_ ,
  \catchup.catchup_reservation_n_isrc1__47_ ,\catchup.catchup_reservation_n_isrc1__46_ ,
  \catchup.catchup_reservation_n_isrc1__45_ ,\catchup.catchup_reservation_n_isrc1__44_ ,
  \catchup.catchup_reservation_n_isrc1__43_ ,\catchup.catchup_reservation_n_isrc1__42_ ,
  \catchup.catchup_reservation_n_isrc1__41_ ,
  \catchup.catchup_reservation_n_isrc1__40_ ,\catchup.catchup_reservation_n_isrc1__39_ ,
  \catchup.catchup_reservation_n_isrc1__38_ ,\catchup.catchup_reservation_n_isrc1__37_ ,
  \catchup.catchup_reservation_n_isrc1__36_ ,\catchup.catchup_reservation_n_isrc1__35_ ,
  \catchup.catchup_reservation_n_isrc1__34_ ,\catchup.catchup_reservation_n_isrc1__33_ ,
  \catchup.catchup_reservation_n_isrc1__32_ ,\catchup.catchup_reservation_n_isrc1__31_ ,
  \catchup.catchup_reservation_n_isrc1__30_ ,\catchup.catchup_reservation_n_isrc1__29_ ,
  \catchup.catchup_reservation_n_isrc1__28_ ,
  \catchup.catchup_reservation_n_isrc1__27_ ,\catchup.catchup_reservation_n_isrc1__26_ ,
  \catchup.catchup_reservation_n_isrc1__25_ ,\catchup.catchup_reservation_n_isrc1__24_ ,
  \catchup.catchup_reservation_n_isrc1__23_ ,\catchup.catchup_reservation_n_isrc1__22_ ,
  \catchup.catchup_reservation_n_isrc1__21_ ,\catchup.catchup_reservation_n_isrc1__20_ ,
  \catchup.catchup_reservation_n_isrc1__19_ ,\catchup.catchup_reservation_n_isrc1__18_ ,
  \catchup.catchup_reservation_n_isrc1__17_ ,\catchup.catchup_reservation_n_isrc1__16_ ,
  \catchup.catchup_reservation_n_isrc1__15_ ,
  \catchup.catchup_reservation_n_isrc1__14_ ,\catchup.catchup_reservation_n_isrc1__13_ ,
  \catchup.catchup_reservation_n_isrc1__12_ ,\catchup.catchup_reservation_n_isrc1__11_ ,
  \catchup.catchup_reservation_n_isrc1__10_ ,\catchup.catchup_reservation_n_isrc1__9_ ,
  \catchup.catchup_reservation_n_isrc1__8_ ,\catchup.catchup_reservation_n_isrc1__7_ ,
  \catchup.catchup_reservation_n_isrc1__6_ ,\catchup.catchup_reservation_n_isrc1__5_ ,
  \catchup.catchup_reservation_n_isrc1__4_ ,\catchup.catchup_reservation_n_isrc1__3_ ,
  \catchup.catchup_reservation_n_isrc1__2_ ,\catchup.catchup_reservation_n_isrc1__1_ ,
  \catchup.catchup_reservation_n_isrc1__0_ ,\catchup.catchup_reservation_n_isrc2__64_ ,
  \catchup.catchup_reservation_n_isrc2__63_ ,
  \catchup.catchup_reservation_n_isrc2__62_ ,\catchup.catchup_reservation_n_isrc2__61_ ,
  \catchup.catchup_reservation_n_isrc2__60_ ,\catchup.catchup_reservation_n_isrc2__59_ ,
  \catchup.catchup_reservation_n_isrc2__58_ ,\catchup.catchup_reservation_n_isrc2__57_ ,
  \catchup.catchup_reservation_n_isrc2__56_ ,\catchup.catchup_reservation_n_isrc2__55_ ,
  \catchup.catchup_reservation_n_isrc2__54_ ,\catchup.catchup_reservation_n_isrc2__53_ ,
  \catchup.catchup_reservation_n_isrc2__52_ ,\catchup.catchup_reservation_n_isrc2__51_ ,
  \catchup.catchup_reservation_n_isrc2__50_ ,
  \catchup.catchup_reservation_n_isrc2__49_ ,\catchup.catchup_reservation_n_isrc2__48_ ,
  \catchup.catchup_reservation_n_isrc2__47_ ,\catchup.catchup_reservation_n_isrc2__46_ ,
  \catchup.catchup_reservation_n_isrc2__45_ ,\catchup.catchup_reservation_n_isrc2__44_ ,
  \catchup.catchup_reservation_n_isrc2__43_ ,\catchup.catchup_reservation_n_isrc2__42_ ,
  \catchup.catchup_reservation_n_isrc2__41_ ,\catchup.catchup_reservation_n_isrc2__40_ ,
  \catchup.catchup_reservation_n_isrc2__39_ ,\catchup.catchup_reservation_n_isrc2__38_ ,
  \catchup.catchup_reservation_n_isrc2__37_ ,\catchup.catchup_reservation_n_isrc2__36_ ,
  \catchup.catchup_reservation_n_isrc2__35_ ,
  \catchup.catchup_reservation_n_isrc2__34_ ,\catchup.catchup_reservation_n_isrc2__33_ ,
  \catchup.catchup_reservation_n_isrc2__32_ ,\catchup.catchup_reservation_n_isrc2__31_ ,
  \catchup.catchup_reservation_n_isrc2__30_ ,\catchup.catchup_reservation_n_isrc2__29_ ,
  \catchup.catchup_reservation_n_isrc2__28_ ,\catchup.catchup_reservation_n_isrc2__27_ ,
  \catchup.catchup_reservation_n_isrc2__26_ ,\catchup.catchup_reservation_n_isrc2__25_ ,
  \catchup.catchup_reservation_n_isrc2__24_ ,\catchup.catchup_reservation_n_isrc2__23_ ,
  \catchup.catchup_reservation_n_isrc2__22_ ,
  \catchup.catchup_reservation_n_isrc2__21_ ,\catchup.catchup_reservation_n_isrc2__20_ ,
  \catchup.catchup_reservation_n_isrc2__19_ ,\catchup.catchup_reservation_n_isrc2__18_ ,
  \catchup.catchup_reservation_n_isrc2__17_ ,\catchup.catchup_reservation_n_isrc2__16_ ,
  \catchup.catchup_reservation_n_isrc2__15_ ,\catchup.catchup_reservation_n_isrc2__14_ ,
  \catchup.catchup_reservation_n_isrc2__13_ ,\catchup.catchup_reservation_n_isrc2__12_ ,
  \catchup.catchup_reservation_n_isrc2__11_ ,\catchup.catchup_reservation_n_isrc2__10_ ,
  \catchup.catchup_reservation_n_isrc2__9_ ,
  \catchup.catchup_reservation_n_isrc2__8_ ,\catchup.catchup_reservation_n_isrc2__7_ ,
  \catchup.catchup_reservation_n_isrc2__6_ ,\catchup.catchup_reservation_n_isrc2__5_ ,
  \catchup.catchup_reservation_n_isrc2__4_ ,\catchup.catchup_reservation_n_isrc2__3_ ,
  \catchup.catchup_reservation_n_isrc2__2_ ,\catchup.catchup_reservation_n_isrc2__1_ ,
  \catchup.catchup_reservation_n_isrc2__0_ ,N44,N45,N46,N47,N48,N49,pipe_int_catchup_data_v_lo,
  pipe_int_catchup_branch_lo,pipe_int_catchup_btaken_lo,pipe_int_catchup_instr_misaligned_lo,
  N50,pipe_int_catchup_mispredict_lo,N51,N52,pipe_aux_fflags_lo_nv_,
  pipe_aux_fflags_lo_dz_,pipe_aux_fflags_lo_of_,pipe_aux_fflags_lo_uf_,pipe_aux_fflags_lo_nx_,
  pipe_aux_data_v_lo,pipe_mem_dtlb_store_miss_lo,pipe_mem_dtlb_load_miss_lo,
  pipe_mem_dcache_replay_lo,pipe_mem_dcache_miss_lo,pipe_mem_load_misaligned_lo,
  pipe_mem_load_access_fault_lo,pipe_mem_load_page_fault_lo,pipe_mem_store_misaligned_lo,
  pipe_mem_store_access_fault_lo,pipe_mem_store_page_fault_lo,
  pipe_mem_early_data_v_lo,pipe_mem_final_data_v_lo,pipe_mul_data_v_lo,pipe_fma_fflags_lo_nv_,
  pipe_fma_fflags_lo_dz_,pipe_fma_fflags_lo_of_,pipe_fma_fflags_lo_uf_,
  pipe_fma_fflags_lo_nx_,pipe_fma_data_v_lo,pipe_long_idata_yumi_lo,pipe_long_fdata_yumi_lo,injection,
  N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,
  N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,
  N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,
  N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,
  N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,
  N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,
  N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,
  N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,
  N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,
  N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,
  N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,
  N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,
  N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
  N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,
  N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,
  N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,
  N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,
  N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,
  N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,
  N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,
  N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,
  N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,
  N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,
  N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,
  N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,
  N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,
  N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,
  N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
  N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,
  N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,
  N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,
  N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
  N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,
  N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,
  N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,
  N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,
  N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,
  N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,
  N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,
  N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,
  N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,
  N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
  N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,
  N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,
  N766,N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,
  N782,N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,
  N798,N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,
  N814,N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,
  N830,N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,
  N846,N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,
  N862,N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,
  N878,exc_stage_n_5__v_,exc_stage_n_5__queue_v_,exc_stage_n_5__ispec_v_,
  exc_stage_n_5__nspec_v_,exc_stage_n_5__exc__store_page_fault_,
  exc_stage_n_5__exc__load_page_fault_,exc_stage_n_5__exc__instr_page_fault_,exc_stage_n_5__exc__ecall_m_,
  exc_stage_n_5__exc__ecall_s_,exc_stage_n_5__exc__ecall_u_,
  exc_stage_n_5__exc__store_access_fault_,exc_stage_n_5__exc__store_misaligned_,
  exc_stage_n_5__exc__load_access_fault_,exc_stage_n_5__exc__load_misaligned_,exc_stage_n_5__exc__ebreak_,
  exc_stage_n_5__exc__illegal_instr_,exc_stage_n_5__exc__instr_access_fault_,
  exc_stage_n_5__exc__instr_misaligned_,exc_stage_n_5__exc__resume_,
  exc_stage_n_5__exc__itlb_miss_,exc_stage_n_5__exc__icache_miss_,exc_stage_n_5__exc__dcache_replay_,
  exc_stage_n_5__exc__dtlb_load_miss_,exc_stage_n_5__exc__dtlb_store_miss_,
  exc_stage_n_5__exc__itlb_fill_,exc_stage_n_5__exc__dtlb_fill_,exc_stage_n_5__exc___interrupt_,
  exc_stage_n_5__exc__cmd_full_,exc_stage_n_5__exc__mispredict_,
  exc_stage_n_5__spec__dcache_miss_,exc_stage_n_5__spec__fencei_,exc_stage_n_5__spec__sfence_vma_,
  exc_stage_n_5__spec__dbreak_,exc_stage_n_5__spec__dret_,
  exc_stage_n_5__spec__mret_,exc_stage_n_5__spec__sret_,exc_stage_n_5__spec__wfi_,
  exc_stage_n_5__spec__csrw_,exc_stage_n_4__v_,exc_stage_n_4__queue_v_,exc_stage_n_4__ispec_v_,
  exc_stage_n_4__nspec_v_,exc_stage_n_4__exc__store_page_fault_,
  exc_stage_n_4__exc__load_page_fault_,exc_stage_n_4__exc__instr_page_fault_,exc_stage_n_4__exc__ecall_m_,
  exc_stage_n_4__exc__ecall_s_,exc_stage_n_4__exc__ecall_u_,
  exc_stage_n_4__exc__store_access_fault_,exc_stage_n_4__exc__store_misaligned_,
  exc_stage_n_4__exc__load_access_fault_,exc_stage_n_4__exc__load_misaligned_,exc_stage_n_4__exc__ebreak_,
  exc_stage_n_4__exc__illegal_instr_,exc_stage_n_4__exc__instr_access_fault_,
  exc_stage_n_4__exc__instr_misaligned_,exc_stage_n_4__exc__resume_,
  exc_stage_n_4__exc__itlb_miss_,exc_stage_n_4__exc__icache_miss_,exc_stage_n_4__exc__dcache_replay_,
  exc_stage_n_4__exc__dtlb_load_miss_,exc_stage_n_4__exc__dtlb_store_miss_,
  exc_stage_n_4__exc__itlb_fill_,exc_stage_n_4__exc__dtlb_fill_,exc_stage_n_4__exc___interrupt_,
  exc_stage_n_4__exc__cmd_full_,exc_stage_n_4__exc__mispredict_,
  exc_stage_n_4__spec__dcache_miss_,exc_stage_n_4__spec__fencei_,exc_stage_n_4__spec__sfence_vma_,
  exc_stage_n_4__spec__dbreak_,exc_stage_n_4__spec__dret_,
  exc_stage_n_4__spec__mret_,exc_stage_n_4__spec__sret_,exc_stage_n_4__spec__wfi_,
  exc_stage_n_4__spec__csrw_,exc_stage_n_3__v_,exc_stage_n_3__queue_v_,exc_stage_n_3__ispec_v_,
  exc_stage_n_3__nspec_v_,exc_stage_n_3__exc__store_page_fault_,
  exc_stage_n_3__exc__load_page_fault_,exc_stage_n_3__exc__instr_page_fault_,exc_stage_n_3__exc__ecall_m_,
  exc_stage_n_3__exc__ecall_s_,exc_stage_n_3__exc__ecall_u_,
  exc_stage_n_3__exc__store_access_fault_,exc_stage_n_3__exc__store_misaligned_,
  exc_stage_n_3__exc__load_access_fault_,exc_stage_n_3__exc__load_misaligned_,exc_stage_n_3__exc__ebreak_,
  exc_stage_n_3__exc__illegal_instr_,exc_stage_n_3__exc__instr_access_fault_,
  exc_stage_n_3__exc__instr_misaligned_,exc_stage_n_3__exc__resume_,
  exc_stage_n_3__exc__itlb_miss_,exc_stage_n_3__exc__icache_miss_,exc_stage_n_3__exc__dcache_replay_,
  exc_stage_n_3__exc__dtlb_load_miss_,exc_stage_n_3__exc__dtlb_store_miss_,
  exc_stage_n_3__exc__itlb_fill_,exc_stage_n_3__exc__dtlb_fill_,exc_stage_n_3__exc___interrupt_,
  exc_stage_n_3__exc__cmd_full_,exc_stage_n_3__exc__mispredict_,
  exc_stage_n_3__spec__dcache_miss_,exc_stage_n_3__spec__fencei_,exc_stage_n_3__spec__sfence_vma_,
  exc_stage_n_3__spec__dbreak_,exc_stage_n_3__spec__dret_,
  exc_stage_n_3__spec__mret_,exc_stage_n_3__spec__sret_,exc_stage_n_3__spec__wfi_,
  exc_stage_n_3__spec__csrw_,exc_stage_n_2__v_,exc_stage_n_2__queue_v_,exc_stage_n_2__ispec_v_,
  exc_stage_n_2__nspec_v_,exc_stage_n_2__exc__store_page_fault_,
  exc_stage_n_2__exc__load_page_fault_,exc_stage_n_2__exc__instr_page_fault_,exc_stage_n_2__exc__ecall_m_,
  exc_stage_n_2__exc__ecall_s_,exc_stage_n_2__exc__ecall_u_,
  exc_stage_n_2__exc__store_access_fault_,exc_stage_n_2__exc__store_misaligned_,
  exc_stage_n_2__exc__load_access_fault_,exc_stage_n_2__exc__load_misaligned_,exc_stage_n_2__exc__ebreak_,
  exc_stage_n_2__exc__illegal_instr_,exc_stage_n_2__exc__instr_access_fault_,
  exc_stage_n_2__exc__instr_misaligned_,exc_stage_n_2__exc__resume_,
  exc_stage_n_2__exc__itlb_miss_,exc_stage_n_2__exc__icache_miss_,exc_stage_n_2__exc__dcache_replay_,
  exc_stage_n_2__exc__dtlb_load_miss_,exc_stage_n_2__exc__dtlb_store_miss_,
  exc_stage_n_2__exc__itlb_fill_,exc_stage_n_2__exc__dtlb_fill_,exc_stage_n_2__exc___interrupt_,
  exc_stage_n_2__exc__cmd_full_,exc_stage_n_2__exc__mispredict_,
  exc_stage_n_2__spec__dcache_miss_,exc_stage_n_2__spec__fencei_,exc_stage_n_2__spec__sfence_vma_,
  exc_stage_n_2__spec__dbreak_,exc_stage_n_2__spec__dret_,
  exc_stage_n_2__spec__mret_,exc_stage_n_2__spec__sret_,exc_stage_n_2__spec__wfi_,
  exc_stage_n_2__spec__csrw_,exc_stage_n_1__v_,exc_stage_n_1__queue_v_,exc_stage_n_1__ispec_v_,
  exc_stage_n_1__nspec_v_,exc_stage_n_1__exc__store_page_fault_,
  exc_stage_n_1__exc__load_page_fault_,exc_stage_n_1__exc__instr_page_fault_,exc_stage_n_1__exc__ecall_m_,
  exc_stage_n_1__exc__ecall_s_,exc_stage_n_1__exc__ecall_u_,
  exc_stage_n_1__exc__store_access_fault_,exc_stage_n_1__exc__store_misaligned_,
  exc_stage_n_1__exc__load_access_fault_,exc_stage_n_1__exc__load_misaligned_,exc_stage_n_1__exc__ebreak_,
  exc_stage_n_1__exc__illegal_instr_,exc_stage_n_1__exc__instr_access_fault_,
  exc_stage_n_1__exc__instr_misaligned_,exc_stage_n_1__exc__resume_,
  exc_stage_n_1__exc__itlb_miss_,exc_stage_n_1__exc__icache_miss_,exc_stage_n_1__exc__dcache_replay_,
  exc_stage_n_1__exc__dtlb_load_miss_,exc_stage_n_1__exc__dtlb_store_miss_,
  exc_stage_n_1__exc__itlb_fill_,exc_stage_n_1__exc__dtlb_fill_,exc_stage_n_1__exc___interrupt_,
  exc_stage_n_1__exc__cmd_full_,exc_stage_n_1__exc__mispredict_,
  exc_stage_n_1__spec__dcache_miss_,exc_stage_n_1__spec__fencei_,exc_stage_n_1__spec__sfence_vma_,
  exc_stage_n_1__spec__dbreak_,exc_stage_n_1__spec__dret_,
  exc_stage_n_1__spec__mret_,exc_stage_n_1__spec__sret_,exc_stage_n_1__spec__wfi_,
  exc_stage_n_1__spec__csrw_,exc_stage_n_0__v_,exc_stage_n_0__queue_v_,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969;
  wire [5:0] \pencode_0_.match_rs_onehot ,\pencode_1_.match_rs_onehot ,
  \pencode_2_.match_rs_onehot ;
  wire [197:0] bypass_rs;
  wire [520:0] reservation_r,\catchup.catchup_reservation_r ;
  wire [65:0] pipe_sys_data_lo,pipe_int_early_data_lo,pipe_int_catchup_data_lo,
  pipe_aux_data_lo,pipe_mem_early_data_lo,pipe_mem_final_data_lo,pipe_mul_data_lo,
  pipe_fma_data_lo;
  wire [2:0] frm_dyn_lo,late_wb_grants_lo;
  wire [64:0] \catchup.catchup_bypass_src1 ,\catchup.catchup_bypass_src2 ;
  wire [38:0] pipe_int_catchup_npc_lo;
  wire [63:0] rs2_val_r;
  wire [2:1] late_wb_reqs_li;
  assign N21 = dispatch_pkt_i[310:306] == { comp_stage_n_1__rd_addr__4_, comp_stage_n_1__rd_addr__3_, comp_stage_n_1__rd_addr__2_, comp_stage_n_1__rd_addr__1_, comp_stage_n_1__rd_addr__0_ };
  assign N22 = dispatch_pkt_i[310:306] == { comp_stage_n_1__rd_addr__4_, comp_stage_n_1__rd_addr__3_, comp_stage_n_1__rd_addr__2_, comp_stage_n_1__rd_addr__1_, comp_stage_n_1__rd_addr__0_ };
  assign N23 = dispatch_pkt_i[315:311] == { comp_stage_n_1__rd_addr__4_, comp_stage_n_1__rd_addr__3_, comp_stage_n_1__rd_addr__2_, comp_stage_n_1__rd_addr__1_, comp_stage_n_1__rd_addr__0_ };
  assign N24 = dispatch_pkt_i[315:311] == { comp_stage_n_1__rd_addr__4_, comp_stage_n_1__rd_addr__3_, comp_stage_n_1__rd_addr__2_, comp_stage_n_1__rd_addr__1_, comp_stage_n_1__rd_addr__0_ };
  assign N25 = dispatch_pkt_i[322:318] == { comp_stage_n_1__rd_addr__4_, comp_stage_n_1__rd_addr__3_, comp_stage_n_1__rd_addr__2_, comp_stage_n_1__rd_addr__1_, comp_stage_n_1__rd_addr__0_ };
  assign N26 = dispatch_pkt_i[310:306] == { comp_stage_n_2__rd_addr__4_, comp_stage_n_2__rd_addr__3_, comp_stage_n_2__rd_addr__2_, comp_stage_n_2__rd_addr__1_, comp_stage_n_2__rd_addr__0_ };
  assign N27 = dispatch_pkt_i[310:306] == { comp_stage_n_2__rd_addr__4_, comp_stage_n_2__rd_addr__3_, comp_stage_n_2__rd_addr__2_, comp_stage_n_2__rd_addr__1_, comp_stage_n_2__rd_addr__0_ };
  assign N28 = dispatch_pkt_i[315:311] == { comp_stage_n_2__rd_addr__4_, comp_stage_n_2__rd_addr__3_, comp_stage_n_2__rd_addr__2_, comp_stage_n_2__rd_addr__1_, comp_stage_n_2__rd_addr__0_ };
  assign N29 = dispatch_pkt_i[315:311] == { comp_stage_n_2__rd_addr__4_, comp_stage_n_2__rd_addr__3_, comp_stage_n_2__rd_addr__2_, comp_stage_n_2__rd_addr__1_, comp_stage_n_2__rd_addr__0_ };
  assign N30 = dispatch_pkt_i[322:318] == { comp_stage_n_2__rd_addr__4_, comp_stage_n_2__rd_addr__3_, comp_stage_n_2__rd_addr__2_, comp_stage_n_2__rd_addr__1_, comp_stage_n_2__rd_addr__0_ };
  assign N31 = dispatch_pkt_i[310:306] == { comp_stage_n_3__rd_addr__4_, comp_stage_n_3__rd_addr__3_, comp_stage_n_3__rd_addr__2_, comp_stage_n_3__rd_addr__1_, comp_stage_n_3__rd_addr__0_ };
  assign N32 = dispatch_pkt_i[310:306] == { comp_stage_n_3__rd_addr__4_, comp_stage_n_3__rd_addr__3_, comp_stage_n_3__rd_addr__2_, comp_stage_n_3__rd_addr__1_, comp_stage_n_3__rd_addr__0_ };
  assign N33 = dispatch_pkt_i[315:311] == { comp_stage_n_3__rd_addr__4_, comp_stage_n_3__rd_addr__3_, comp_stage_n_3__rd_addr__2_, comp_stage_n_3__rd_addr__1_, comp_stage_n_3__rd_addr__0_ };
  assign N34 = dispatch_pkt_i[315:311] == { comp_stage_n_3__rd_addr__4_, comp_stage_n_3__rd_addr__3_, comp_stage_n_3__rd_addr__2_, comp_stage_n_3__rd_addr__1_, comp_stage_n_3__rd_addr__0_ };
  assign N35 = dispatch_pkt_i[322:318] == { comp_stage_n_3__rd_addr__4_, comp_stage_n_3__rd_addr__3_, comp_stage_n_3__rd_addr__2_, comp_stage_n_3__rd_addr__1_, comp_stage_n_3__rd_addr__0_ };
  assign N36 = dispatch_pkt_i[310:306] == iwb_pkt_o[75:71];
  assign N37 = dispatch_pkt_i[310:306] == iwb_pkt_o[75:71];
  assign N38 = dispatch_pkt_i[315:311] == iwb_pkt_o[75:71];
  assign N39 = dispatch_pkt_i[315:311] == iwb_pkt_o[75:71];
  assign N40 = dispatch_pkt_i[322:318] == iwb_pkt_o[75:71];
  assign N41 = dispatch_pkt_i[310:306] == fwb_pkt_o[75:71];
  assign N42 = dispatch_pkt_i[315:311] == fwb_pkt_o[75:71];
  assign N43 = dispatch_pkt_i[322:318] == fwb_pkt_o[75:71];

  bsg_priority_encode_one_hot_out_width_p6_lo_to_hi_p1
  \pencode_0_.pencode_oh 
  (
    .i({ 1'b1, match_rs[4:0] }),
    .o(\pencode_0_.match_rs_onehot )
  );


  bsg_mux_one_hot_width_p66_els_p6
  \pencode_0_.fwd_mux_oh 
  (
    .data_i({ dispatch_pkt_i[231:166], fwb_pkt_o[70:5], forward_data_3__65_, forward_data_3__64_, forward_data_3__63_, forward_data_3__62_, forward_data_3__61_, forward_data_3__60_, forward_data_3__59_, forward_data_3__58_, forward_data_3__57_, forward_data_3__56_, forward_data_3__55_, forward_data_3__54_, forward_data_3__53_, forward_data_3__52_, forward_data_3__51_, forward_data_3__50_, forward_data_3__49_, forward_data_3__48_, forward_data_3__47_, forward_data_3__46_, forward_data_3__45_, forward_data_3__44_, forward_data_3__43_, forward_data_3__42_, forward_data_3__41_, forward_data_3__40_, forward_data_3__39_, forward_data_3__38_, forward_data_3__37_, forward_data_3__36_, forward_data_3__35_, forward_data_3__34_, forward_data_3__33_, forward_data_3__32_, forward_data_3__31_, forward_data_3__30_, forward_data_3__29_, forward_data_3__28_, forward_data_3__27_, forward_data_3__26_, forward_data_3__25_, forward_data_3__24_, forward_data_3__23_, forward_data_3__22_, forward_data_3__21_, forward_data_3__20_, forward_data_3__19_, forward_data_3__18_, forward_data_3__17_, forward_data_3__16_, forward_data_3__15_, forward_data_3__14_, forward_data_3__13_, forward_data_3__12_, forward_data_3__11_, forward_data_3__10_, forward_data_3__9_, forward_data_3__8_, forward_data_3__7_, forward_data_3__6_, forward_data_3__5_, forward_data_3__4_, forward_data_3__3_, forward_data_3__2_, forward_data_3__1_, forward_data_3__0_, forward_data_2__65_, forward_data_2__64_, forward_data_2__63_, forward_data_2__62_, forward_data_2__61_, forward_data_2__60_, forward_data_2__59_, forward_data_2__58_, forward_data_2__57_, forward_data_2__56_, forward_data_2__55_, forward_data_2__54_, forward_data_2__53_, forward_data_2__52_, forward_data_2__51_, forward_data_2__50_, forward_data_2__49_, forward_data_2__48_, forward_data_2__47_, forward_data_2__46_, forward_data_2__45_, forward_data_2__44_, forward_data_2__43_, forward_data_2__42_, forward_data_2__41_, forward_data_2__40_, forward_data_2__39_, forward_data_2__38_, forward_data_2__37_, forward_data_2__36_, forward_data_2__35_, forward_data_2__34_, forward_data_2__33_, forward_data_2__32_, forward_data_2__31_, forward_data_2__30_, forward_data_2__29_, forward_data_2__28_, forward_data_2__27_, forward_data_2__26_, forward_data_2__25_, forward_data_2__24_, forward_data_2__23_, forward_data_2__22_, forward_data_2__21_, forward_data_2__20_, forward_data_2__19_, forward_data_2__18_, forward_data_2__17_, forward_data_2__16_, forward_data_2__15_, forward_data_2__14_, forward_data_2__13_, forward_data_2__12_, forward_data_2__11_, forward_data_2__10_, forward_data_2__9_, forward_data_2__8_, forward_data_2__7_, forward_data_2__6_, forward_data_2__5_, forward_data_2__4_, forward_data_2__3_, forward_data_2__2_, forward_data_2__1_, forward_data_2__0_, forward_data_1__65_, forward_data_1__64_, forward_data_1__63_, forward_data_1__62_, forward_data_1__61_, forward_data_1__60_, forward_data_1__59_, forward_data_1__58_, forward_data_1__57_, forward_data_1__56_, forward_data_1__55_, forward_data_1__54_, forward_data_1__53_, forward_data_1__52_, forward_data_1__51_, forward_data_1__50_, forward_data_1__49_, forward_data_1__48_, forward_data_1__47_, forward_data_1__46_, forward_data_1__45_, forward_data_1__44_, forward_data_1__43_, forward_data_1__42_, forward_data_1__41_, forward_data_1__40_, forward_data_1__39_, forward_data_1__38_, forward_data_1__37_, forward_data_1__36_, forward_data_1__35_, forward_data_1__34_, forward_data_1__33_, forward_data_1__32_, forward_data_1__31_, forward_data_1__30_, forward_data_1__29_, forward_data_1__28_, forward_data_1__27_, forward_data_1__26_, forward_data_1__25_, forward_data_1__24_, forward_data_1__23_, forward_data_1__22_, forward_data_1__21_, forward_data_1__20_, forward_data_1__19_, forward_data_1__18_, forward_data_1__17_, forward_data_1__16_, forward_data_1__15_, forward_data_1__14_, forward_data_1__13_, forward_data_1__12_, forward_data_1__11_, forward_data_1__10_, forward_data_1__9_, forward_data_1__8_, forward_data_1__7_, forward_data_1__6_, forward_data_1__5_, forward_data_1__4_, forward_data_1__3_, forward_data_1__2_, forward_data_1__1_, forward_data_1__0_, forward_data_0__65_, forward_data_0__64_, forward_data_0__63_, forward_data_0__62_, forward_data_0__61_, forward_data_0__60_, forward_data_0__59_, forward_data_0__58_, forward_data_0__57_, forward_data_0__56_, forward_data_0__55_, forward_data_0__54_, forward_data_0__53_, forward_data_0__52_, forward_data_0__51_, forward_data_0__50_, forward_data_0__49_, forward_data_0__48_, forward_data_0__47_, forward_data_0__46_, forward_data_0__45_, forward_data_0__44_, forward_data_0__43_, forward_data_0__42_, forward_data_0__41_, forward_data_0__40_, forward_data_0__39_, forward_data_0__38_, forward_data_0__37_, forward_data_0__36_, forward_data_0__35_, forward_data_0__34_, forward_data_0__33_, forward_data_0__32_, forward_data_0__31_, forward_data_0__30_, forward_data_0__29_, forward_data_0__28_, forward_data_0__27_, forward_data_0__26_, forward_data_0__25_, forward_data_0__24_, forward_data_0__23_, forward_data_0__22_, forward_data_0__21_, forward_data_0__20_, forward_data_0__19_, forward_data_0__18_, forward_data_0__17_, forward_data_0__16_, forward_data_0__15_, forward_data_0__14_, forward_data_0__13_, forward_data_0__12_, forward_data_0__11_, forward_data_0__10_, forward_data_0__9_, forward_data_0__8_, forward_data_0__7_, forward_data_0__6_, forward_data_0__5_, forward_data_0__4_, forward_data_0__3_, forward_data_0__2_, forward_data_0__1_, forward_data_0__0_ }),
    .sel_one_hot_i(\pencode_0_.match_rs_onehot ),
    .data_o(bypass_rs[65:0])
  );


  bsg_priority_encode_one_hot_out_width_p6_lo_to_hi_p1
  \pencode_1_.pencode_oh 
  (
    .i({ 1'b1, match_rs[9:5] }),
    .o(\pencode_1_.match_rs_onehot )
  );


  bsg_mux_one_hot_width_p66_els_p6
  \pencode_1_.fwd_mux_oh 
  (
    .data_i({ dispatch_pkt_i[165:100], fwb_pkt_o[70:5], forward_data_3__65_, forward_data_3__64_, forward_data_3__63_, forward_data_3__62_, forward_data_3__61_, forward_data_3__60_, forward_data_3__59_, forward_data_3__58_, forward_data_3__57_, forward_data_3__56_, forward_data_3__55_, forward_data_3__54_, forward_data_3__53_, forward_data_3__52_, forward_data_3__51_, forward_data_3__50_, forward_data_3__49_, forward_data_3__48_, forward_data_3__47_, forward_data_3__46_, forward_data_3__45_, forward_data_3__44_, forward_data_3__43_, forward_data_3__42_, forward_data_3__41_, forward_data_3__40_, forward_data_3__39_, forward_data_3__38_, forward_data_3__37_, forward_data_3__36_, forward_data_3__35_, forward_data_3__34_, forward_data_3__33_, forward_data_3__32_, forward_data_3__31_, forward_data_3__30_, forward_data_3__29_, forward_data_3__28_, forward_data_3__27_, forward_data_3__26_, forward_data_3__25_, forward_data_3__24_, forward_data_3__23_, forward_data_3__22_, forward_data_3__21_, forward_data_3__20_, forward_data_3__19_, forward_data_3__18_, forward_data_3__17_, forward_data_3__16_, forward_data_3__15_, forward_data_3__14_, forward_data_3__13_, forward_data_3__12_, forward_data_3__11_, forward_data_3__10_, forward_data_3__9_, forward_data_3__8_, forward_data_3__7_, forward_data_3__6_, forward_data_3__5_, forward_data_3__4_, forward_data_3__3_, forward_data_3__2_, forward_data_3__1_, forward_data_3__0_, forward_data_2__65_, forward_data_2__64_, forward_data_2__63_, forward_data_2__62_, forward_data_2__61_, forward_data_2__60_, forward_data_2__59_, forward_data_2__58_, forward_data_2__57_, forward_data_2__56_, forward_data_2__55_, forward_data_2__54_, forward_data_2__53_, forward_data_2__52_, forward_data_2__51_, forward_data_2__50_, forward_data_2__49_, forward_data_2__48_, forward_data_2__47_, forward_data_2__46_, forward_data_2__45_, forward_data_2__44_, forward_data_2__43_, forward_data_2__42_, forward_data_2__41_, forward_data_2__40_, forward_data_2__39_, forward_data_2__38_, forward_data_2__37_, forward_data_2__36_, forward_data_2__35_, forward_data_2__34_, forward_data_2__33_, forward_data_2__32_, forward_data_2__31_, forward_data_2__30_, forward_data_2__29_, forward_data_2__28_, forward_data_2__27_, forward_data_2__26_, forward_data_2__25_, forward_data_2__24_, forward_data_2__23_, forward_data_2__22_, forward_data_2__21_, forward_data_2__20_, forward_data_2__19_, forward_data_2__18_, forward_data_2__17_, forward_data_2__16_, forward_data_2__15_, forward_data_2__14_, forward_data_2__13_, forward_data_2__12_, forward_data_2__11_, forward_data_2__10_, forward_data_2__9_, forward_data_2__8_, forward_data_2__7_, forward_data_2__6_, forward_data_2__5_, forward_data_2__4_, forward_data_2__3_, forward_data_2__2_, forward_data_2__1_, forward_data_2__0_, forward_data_1__65_, forward_data_1__64_, forward_data_1__63_, forward_data_1__62_, forward_data_1__61_, forward_data_1__60_, forward_data_1__59_, forward_data_1__58_, forward_data_1__57_, forward_data_1__56_, forward_data_1__55_, forward_data_1__54_, forward_data_1__53_, forward_data_1__52_, forward_data_1__51_, forward_data_1__50_, forward_data_1__49_, forward_data_1__48_, forward_data_1__47_, forward_data_1__46_, forward_data_1__45_, forward_data_1__44_, forward_data_1__43_, forward_data_1__42_, forward_data_1__41_, forward_data_1__40_, forward_data_1__39_, forward_data_1__38_, forward_data_1__37_, forward_data_1__36_, forward_data_1__35_, forward_data_1__34_, forward_data_1__33_, forward_data_1__32_, forward_data_1__31_, forward_data_1__30_, forward_data_1__29_, forward_data_1__28_, forward_data_1__27_, forward_data_1__26_, forward_data_1__25_, forward_data_1__24_, forward_data_1__23_, forward_data_1__22_, forward_data_1__21_, forward_data_1__20_, forward_data_1__19_, forward_data_1__18_, forward_data_1__17_, forward_data_1__16_, forward_data_1__15_, forward_data_1__14_, forward_data_1__13_, forward_data_1__12_, forward_data_1__11_, forward_data_1__10_, forward_data_1__9_, forward_data_1__8_, forward_data_1__7_, forward_data_1__6_, forward_data_1__5_, forward_data_1__4_, forward_data_1__3_, forward_data_1__2_, forward_data_1__1_, forward_data_1__0_, forward_data_0__65_, forward_data_0__64_, forward_data_0__63_, forward_data_0__62_, forward_data_0__61_, forward_data_0__60_, forward_data_0__59_, forward_data_0__58_, forward_data_0__57_, forward_data_0__56_, forward_data_0__55_, forward_data_0__54_, forward_data_0__53_, forward_data_0__52_, forward_data_0__51_, forward_data_0__50_, forward_data_0__49_, forward_data_0__48_, forward_data_0__47_, forward_data_0__46_, forward_data_0__45_, forward_data_0__44_, forward_data_0__43_, forward_data_0__42_, forward_data_0__41_, forward_data_0__40_, forward_data_0__39_, forward_data_0__38_, forward_data_0__37_, forward_data_0__36_, forward_data_0__35_, forward_data_0__34_, forward_data_0__33_, forward_data_0__32_, forward_data_0__31_, forward_data_0__30_, forward_data_0__29_, forward_data_0__28_, forward_data_0__27_, forward_data_0__26_, forward_data_0__25_, forward_data_0__24_, forward_data_0__23_, forward_data_0__22_, forward_data_0__21_, forward_data_0__20_, forward_data_0__19_, forward_data_0__18_, forward_data_0__17_, forward_data_0__16_, forward_data_0__15_, forward_data_0__14_, forward_data_0__13_, forward_data_0__12_, forward_data_0__11_, forward_data_0__10_, forward_data_0__9_, forward_data_0__8_, forward_data_0__7_, forward_data_0__6_, forward_data_0__5_, forward_data_0__4_, forward_data_0__3_, forward_data_0__2_, forward_data_0__1_, forward_data_0__0_ }),
    .sel_one_hot_i(\pencode_1_.match_rs_onehot ),
    .data_o(bypass_rs[131:66])
  );


  bsg_priority_encode_one_hot_out_width_p6_lo_to_hi_p1
  \pencode_2_.pencode_oh 
  (
    .i({ 1'b1, match_rs[14:10] }),
    .o(\pencode_2_.match_rs_onehot )
  );


  bsg_mux_one_hot_width_p66_els_p6
  \pencode_2_.fwd_mux_oh 
  (
    .data_i({ dispatch_pkt_i[99:34], fwb_pkt_o[70:5], forward_data_3__65_, forward_data_3__64_, forward_data_3__63_, forward_data_3__62_, forward_data_3__61_, forward_data_3__60_, forward_data_3__59_, forward_data_3__58_, forward_data_3__57_, forward_data_3__56_, forward_data_3__55_, forward_data_3__54_, forward_data_3__53_, forward_data_3__52_, forward_data_3__51_, forward_data_3__50_, forward_data_3__49_, forward_data_3__48_, forward_data_3__47_, forward_data_3__46_, forward_data_3__45_, forward_data_3__44_, forward_data_3__43_, forward_data_3__42_, forward_data_3__41_, forward_data_3__40_, forward_data_3__39_, forward_data_3__38_, forward_data_3__37_, forward_data_3__36_, forward_data_3__35_, forward_data_3__34_, forward_data_3__33_, forward_data_3__32_, forward_data_3__31_, forward_data_3__30_, forward_data_3__29_, forward_data_3__28_, forward_data_3__27_, forward_data_3__26_, forward_data_3__25_, forward_data_3__24_, forward_data_3__23_, forward_data_3__22_, forward_data_3__21_, forward_data_3__20_, forward_data_3__19_, forward_data_3__18_, forward_data_3__17_, forward_data_3__16_, forward_data_3__15_, forward_data_3__14_, forward_data_3__13_, forward_data_3__12_, forward_data_3__11_, forward_data_3__10_, forward_data_3__9_, forward_data_3__8_, forward_data_3__7_, forward_data_3__6_, forward_data_3__5_, forward_data_3__4_, forward_data_3__3_, forward_data_3__2_, forward_data_3__1_, forward_data_3__0_, forward_data_2__65_, forward_data_2__64_, forward_data_2__63_, forward_data_2__62_, forward_data_2__61_, forward_data_2__60_, forward_data_2__59_, forward_data_2__58_, forward_data_2__57_, forward_data_2__56_, forward_data_2__55_, forward_data_2__54_, forward_data_2__53_, forward_data_2__52_, forward_data_2__51_, forward_data_2__50_, forward_data_2__49_, forward_data_2__48_, forward_data_2__47_, forward_data_2__46_, forward_data_2__45_, forward_data_2__44_, forward_data_2__43_, forward_data_2__42_, forward_data_2__41_, forward_data_2__40_, forward_data_2__39_, forward_data_2__38_, forward_data_2__37_, forward_data_2__36_, forward_data_2__35_, forward_data_2__34_, forward_data_2__33_, forward_data_2__32_, forward_data_2__31_, forward_data_2__30_, forward_data_2__29_, forward_data_2__28_, forward_data_2__27_, forward_data_2__26_, forward_data_2__25_, forward_data_2__24_, forward_data_2__23_, forward_data_2__22_, forward_data_2__21_, forward_data_2__20_, forward_data_2__19_, forward_data_2__18_, forward_data_2__17_, forward_data_2__16_, forward_data_2__15_, forward_data_2__14_, forward_data_2__13_, forward_data_2__12_, forward_data_2__11_, forward_data_2__10_, forward_data_2__9_, forward_data_2__8_, forward_data_2__7_, forward_data_2__6_, forward_data_2__5_, forward_data_2__4_, forward_data_2__3_, forward_data_2__2_, forward_data_2__1_, forward_data_2__0_, forward_data_1__65_, forward_data_1__64_, forward_data_1__63_, forward_data_1__62_, forward_data_1__61_, forward_data_1__60_, forward_data_1__59_, forward_data_1__58_, forward_data_1__57_, forward_data_1__56_, forward_data_1__55_, forward_data_1__54_, forward_data_1__53_, forward_data_1__52_, forward_data_1__51_, forward_data_1__50_, forward_data_1__49_, forward_data_1__48_, forward_data_1__47_, forward_data_1__46_, forward_data_1__45_, forward_data_1__44_, forward_data_1__43_, forward_data_1__42_, forward_data_1__41_, forward_data_1__40_, forward_data_1__39_, forward_data_1__38_, forward_data_1__37_, forward_data_1__36_, forward_data_1__35_, forward_data_1__34_, forward_data_1__33_, forward_data_1__32_, forward_data_1__31_, forward_data_1__30_, forward_data_1__29_, forward_data_1__28_, forward_data_1__27_, forward_data_1__26_, forward_data_1__25_, forward_data_1__24_, forward_data_1__23_, forward_data_1__22_, forward_data_1__21_, forward_data_1__20_, forward_data_1__19_, forward_data_1__18_, forward_data_1__17_, forward_data_1__16_, forward_data_1__15_, forward_data_1__14_, forward_data_1__13_, forward_data_1__12_, forward_data_1__11_, forward_data_1__10_, forward_data_1__9_, forward_data_1__8_, forward_data_1__7_, forward_data_1__6_, forward_data_1__5_, forward_data_1__4_, forward_data_1__3_, forward_data_1__2_, forward_data_1__1_, forward_data_1__0_, forward_data_0__65_, forward_data_0__64_, forward_data_0__63_, forward_data_0__62_, forward_data_0__61_, forward_data_0__60_, forward_data_0__59_, forward_data_0__58_, forward_data_0__57_, forward_data_0__56_, forward_data_0__55_, forward_data_0__54_, forward_data_0__53_, forward_data_0__52_, forward_data_0__51_, forward_data_0__50_, forward_data_0__49_, forward_data_0__48_, forward_data_0__47_, forward_data_0__46_, forward_data_0__45_, forward_data_0__44_, forward_data_0__43_, forward_data_0__42_, forward_data_0__41_, forward_data_0__40_, forward_data_0__39_, forward_data_0__38_, forward_data_0__37_, forward_data_0__36_, forward_data_0__35_, forward_data_0__34_, forward_data_0__33_, forward_data_0__32_, forward_data_0__31_, forward_data_0__30_, forward_data_0__29_, forward_data_0__28_, forward_data_0__27_, forward_data_0__26_, forward_data_0__25_, forward_data_0__24_, forward_data_0__23_, forward_data_0__22_, forward_data_0__21_, forward_data_0__20_, forward_data_0__19_, forward_data_0__18_, forward_data_0__17_, forward_data_0__16_, forward_data_0__15_, forward_data_0__14_, forward_data_0__13_, forward_data_0__12_, forward_data_0__11_, forward_data_0__10_, forward_data_0__9_, forward_data_0__8_, forward_data_0__7_, forward_data_0__6_, forward_data_0__5_, forward_data_0__4_, forward_data_0__3_, forward_data_0__2_, forward_data_0__1_, forward_data_0__0_ }),
    .sel_one_hot_i(\pencode_2_.match_rs_onehot ),
    .data_o(bypass_rs[197:132])
  );


  bp_be_reservation_00
  reservation_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .dispatch_pkt_i(dispatch_pkt_i),
    .bypass_rs_i(bypass_rs),
    .reservation_o(reservation_r)
  );


  bp_be_pipe_sys_00
  pipe_sys
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .cfg_bus_i(cfg_bus_i),
    .reservation_i(reservation_r),
    .flush_i(commit_pkt_o[213]),
    .retire_v_i(exc_stage_r_2__v_),
    .retire_queue_v_i(exc_stage_n_3__queue_v_),
    .retire_data_i({ comp_stage_r_2__rd_data__65_, comp_stage_r_2__rd_data__64_, comp_stage_r_2__rd_data__63_, comp_stage_r_2__rd_data__62_, comp_stage_r_2__rd_data__61_, comp_stage_r_2__rd_data__60_, comp_stage_r_2__rd_data__59_, comp_stage_r_2__rd_data__58_, comp_stage_r_2__rd_data__57_, comp_stage_r_2__rd_data__56_, comp_stage_r_2__rd_data__55_, comp_stage_r_2__rd_data__54_, comp_stage_r_2__rd_data__53_, comp_stage_r_2__rd_data__52_, comp_stage_r_2__rd_data__51_, comp_stage_r_2__rd_data__50_, comp_stage_r_2__rd_data__49_, comp_stage_r_2__rd_data__48_, comp_stage_r_2__rd_data__47_, comp_stage_r_2__rd_data__46_, comp_stage_r_2__rd_data__45_, comp_stage_r_2__rd_data__44_, comp_stage_r_2__rd_data__43_, comp_stage_r_2__rd_data__42_, comp_stage_r_2__rd_data__41_, comp_stage_r_2__rd_data__40_, comp_stage_r_2__rd_data__39_, comp_stage_r_2__rd_data__38_, comp_stage_r_2__rd_data__37_, comp_stage_r_2__rd_data__36_, comp_stage_r_2__rd_data__35_, comp_stage_r_2__rd_data__34_, comp_stage_r_2__rd_data__33_, comp_stage_r_2__rd_data__32_, comp_stage_r_2__rd_data__31_, comp_stage_r_2__rd_data__30_, comp_stage_r_2__rd_data__29_, comp_stage_r_2__rd_data__28_, comp_stage_r_2__rd_data__27_, comp_stage_r_2__rd_data__26_, comp_stage_r_2__rd_data__25_, comp_stage_r_2__rd_data__24_, comp_stage_r_2__rd_data__23_, comp_stage_r_2__rd_data__22_, comp_stage_r_2__rd_data__21_, comp_stage_r_2__rd_data__20_, comp_stage_r_2__rd_data__19_, comp_stage_r_2__rd_data__18_, comp_stage_r_2__rd_data__17_, comp_stage_r_2__rd_data__16_, comp_stage_r_2__rd_data__15_, comp_stage_r_2__rd_data__14_, comp_stage_r_2__rd_data__13_, comp_stage_r_2__rd_data__12_, comp_stage_r_2__rd_data__11_, comp_stage_r_2__rd_data__10_, comp_stage_r_2__rd_data__9_, comp_stage_r_2__rd_data__8_, comp_stage_r_2__rd_data__7_, comp_stage_r_2__rd_data__6_, comp_stage_r_2__rd_data__5_, comp_stage_r_2__rd_data__4_, comp_stage_r_2__rd_data__3_, comp_stage_r_2__rd_data__2_, comp_stage_r_2__rd_data__1_, comp_stage_r_2__rd_data__0_ }),
    .retire_exception_i({ exc_stage_n_3__exc__store_page_fault_, exc_stage_n_3__exc__load_page_fault_, exc_stage_n_3__exc__instr_page_fault_, exc_stage_n_3__exc__ecall_m_, exc_stage_n_3__exc__ecall_s_, exc_stage_n_3__exc__ecall_u_, exc_stage_n_3__exc__store_access_fault_, exc_stage_n_3__exc__store_misaligned_, exc_stage_n_3__exc__load_access_fault_, exc_stage_n_3__exc__load_misaligned_, exc_stage_n_3__exc__ebreak_, exc_stage_n_3__exc__illegal_instr_, exc_stage_n_3__exc__instr_access_fault_, exc_stage_n_3__exc__instr_misaligned_, exc_stage_n_3__exc__resume_, exc_stage_n_3__exc__itlb_miss_, exc_stage_n_3__exc__icache_miss_, exc_stage_n_3__exc__dcache_replay_, exc_stage_n_3__exc__dtlb_load_miss_, exc_stage_n_3__exc__dtlb_store_miss_, exc_stage_n_3__exc__itlb_fill_, exc_stage_n_3__exc__dtlb_fill_, exc_stage_n_3__exc___interrupt_, exc_stage_n_3__exc__cmd_full_, exc_stage_n_3__exc__mispredict_ }),
    .retire_special_i({ exc_stage_n_3__spec__dcache_miss_, exc_stage_n_3__spec__fencei_, exc_stage_n_3__spec__sfence_vma_, exc_stage_n_3__spec__dbreak_, exc_stage_n_3__spec__dret_, exc_stage_n_3__spec__mret_, exc_stage_n_3__spec__sret_, exc_stage_n_3__spec__wfi_, exc_stage_n_3__spec__csrw_ }),
    .data_o(pipe_sys_data_lo),
    .v_o(pipe_sys_data_v_lo),
    .illegal_instr_o(pipe_sys_illegal_instr_lo),
    .iwb_pkt_i(iwb_pkt_o),
    .fwb_pkt_i(fwb_pkt_o),
    .commit_pkt_o(commit_pkt_o),
    .debug_irq_i(debug_irq_i),
    .timer_irq_i(timer_irq_i),
    .software_irq_i(software_irq_i),
    .m_external_irq_i(m_external_irq_i),
    .s_external_irq_i(s_external_irq_i),
    .irq_pending_o(irq_pending_o),
    .irq_waiting_o(irq_waiting_o),
    .decode_info_o(decode_info_o),
    .trans_info_o(trans_info_o),
    .frm_dyn_o(frm_dyn_lo)
  );


  bp_be_pipe_int_00
  pipe_int_early
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(_12_net_),
    .reservation_i(reservation_r),
    .flush_i(commit_pkt_o[213]),
    .data_o(pipe_int_early_data_lo),
    .v_o(pipe_int_early_data_v_lo),
    .branch_o(pipe_int_early_branch_lo),
    .btaken_o(pipe_int_early_btaken_lo),
    .npc_o(br_pkt_o[38:0]),
    .instr_misaligned_v_o(pipe_int_early_instr_misaligned_lo)
  );


  bp_be_int_unbox_00
  \catchup.irs1_unbox 
  (
    .reg_i({ forward_data_1__65_, forward_data_1__64_, forward_data_1__63_, forward_data_1__62_, forward_data_1__61_, forward_data_1__60_, forward_data_1__59_, forward_data_1__58_, forward_data_1__57_, forward_data_1__56_, forward_data_1__55_, forward_data_1__54_, forward_data_1__53_, forward_data_1__52_, forward_data_1__51_, forward_data_1__50_, forward_data_1__49_, forward_data_1__48_, forward_data_1__47_, forward_data_1__46_, forward_data_1__45_, forward_data_1__44_, forward_data_1__43_, forward_data_1__42_, forward_data_1__41_, forward_data_1__40_, forward_data_1__39_, forward_data_1__38_, forward_data_1__37_, forward_data_1__36_, forward_data_1__35_, forward_data_1__34_, forward_data_1__33_, forward_data_1__32_, forward_data_1__31_, forward_data_1__30_, forward_data_1__29_, forward_data_1__28_, forward_data_1__27_, forward_data_1__26_, forward_data_1__25_, forward_data_1__24_, forward_data_1__23_, forward_data_1__22_, forward_data_1__21_, forward_data_1__20_, forward_data_1__19_, forward_data_1__18_, forward_data_1__17_, forward_data_1__16_, forward_data_1__15_, forward_data_1__14_, forward_data_1__13_, forward_data_1__12_, forward_data_1__11_, forward_data_1__10_, forward_data_1__9_, forward_data_1__8_, forward_data_1__7_, forward_data_1__6_, forward_data_1__5_, forward_data_1__4_, forward_data_1__3_, forward_data_1__2_, forward_data_1__1_, forward_data_1__0_ }),
    .tag_i(reservation_r[417:416]),
    .unsigned_i(reservation_r[418]),
    .val_o(\catchup.catchup_bypass_src1 )
  );


  bp_be_int_unbox_00
  \catchup.irs2_unbox 
  (
    .reg_i({ forward_data_1__65_, forward_data_1__64_, forward_data_1__63_, forward_data_1__62_, forward_data_1__61_, forward_data_1__60_, forward_data_1__59_, forward_data_1__58_, forward_data_1__57_, forward_data_1__56_, forward_data_1__55_, forward_data_1__54_, forward_data_1__53_, forward_data_1__52_, forward_data_1__51_, forward_data_1__50_, forward_data_1__49_, forward_data_1__48_, forward_data_1__47_, forward_data_1__46_, forward_data_1__45_, forward_data_1__44_, forward_data_1__43_, forward_data_1__42_, forward_data_1__41_, forward_data_1__40_, forward_data_1__39_, forward_data_1__38_, forward_data_1__37_, forward_data_1__36_, forward_data_1__35_, forward_data_1__34_, forward_data_1__33_, forward_data_1__32_, forward_data_1__31_, forward_data_1__30_, forward_data_1__29_, forward_data_1__28_, forward_data_1__27_, forward_data_1__26_, forward_data_1__25_, forward_data_1__24_, forward_data_1__23_, forward_data_1__22_, forward_data_1__21_, forward_data_1__20_, forward_data_1__19_, forward_data_1__18_, forward_data_1__17_, forward_data_1__16_, forward_data_1__15_, forward_data_1__14_, forward_data_1__13_, forward_data_1__12_, forward_data_1__11_, forward_data_1__10_, forward_data_1__9_, forward_data_1__8_, forward_data_1__7_, forward_data_1__6_, forward_data_1__5_, forward_data_1__4_, forward_data_1__3_, forward_data_1__2_, forward_data_1__1_, forward_data_1__0_ }),
    .tag_i(reservation_r[414:413]),
    .unsigned_i(reservation_r[415]),
    .val_o(\catchup.catchup_bypass_src2 )
  );

  assign N44 = { comp_stage_n_2__rd_addr__4_, comp_stage_n_2__rd_addr__3_, comp_stage_n_2__rd_addr__2_, comp_stage_n_2__rd_addr__1_, comp_stage_n_2__rd_addr__0_ } == reservation_r[468:464];
  assign N47 = { comp_stage_n_2__rd_addr__4_, comp_stage_n_2__rd_addr__3_, comp_stage_n_2__rd_addr__2_, comp_stage_n_2__rd_addr__1_, comp_stage_n_2__rd_addr__0_ } == reservation_r[473:469];

  bsg_dff_width_p521
  \catchup.catchup_reservation_reg 
  (
    .clk_i(clk_i),
    .data_i({ reservation_r[520:390], \catchup.catchup_reservation_n_isrc1__64_ , \catchup.catchup_reservation_n_isrc1__63_ , \catchup.catchup_reservation_n_isrc1__62_ , \catchup.catchup_reservation_n_isrc1__61_ , \catchup.catchup_reservation_n_isrc1__60_ , \catchup.catchup_reservation_n_isrc1__59_ , \catchup.catchup_reservation_n_isrc1__58_ , \catchup.catchup_reservation_n_isrc1__57_ , \catchup.catchup_reservation_n_isrc1__56_ , \catchup.catchup_reservation_n_isrc1__55_ , \catchup.catchup_reservation_n_isrc1__54_ , \catchup.catchup_reservation_n_isrc1__53_ , \catchup.catchup_reservation_n_isrc1__52_ , \catchup.catchup_reservation_n_isrc1__51_ , \catchup.catchup_reservation_n_isrc1__50_ , \catchup.catchup_reservation_n_isrc1__49_ , \catchup.catchup_reservation_n_isrc1__48_ , \catchup.catchup_reservation_n_isrc1__47_ , \catchup.catchup_reservation_n_isrc1__46_ , \catchup.catchup_reservation_n_isrc1__45_ , \catchup.catchup_reservation_n_isrc1__44_ , \catchup.catchup_reservation_n_isrc1__43_ , \catchup.catchup_reservation_n_isrc1__42_ , \catchup.catchup_reservation_n_isrc1__41_ , \catchup.catchup_reservation_n_isrc1__40_ , \catchup.catchup_reservation_n_isrc1__39_ , \catchup.catchup_reservation_n_isrc1__38_ , \catchup.catchup_reservation_n_isrc1__37_ , \catchup.catchup_reservation_n_isrc1__36_ , \catchup.catchup_reservation_n_isrc1__35_ , \catchup.catchup_reservation_n_isrc1__34_ , \catchup.catchup_reservation_n_isrc1__33_ , \catchup.catchup_reservation_n_isrc1__32_ , \catchup.catchup_reservation_n_isrc1__31_ , \catchup.catchup_reservation_n_isrc1__30_ , \catchup.catchup_reservation_n_isrc1__29_ , \catchup.catchup_reservation_n_isrc1__28_ , \catchup.catchup_reservation_n_isrc1__27_ , \catchup.catchup_reservation_n_isrc1__26_ , \catchup.catchup_reservation_n_isrc1__25_ , \catchup.catchup_reservation_n_isrc1__24_ , \catchup.catchup_reservation_n_isrc1__23_ , \catchup.catchup_reservation_n_isrc1__22_ , \catchup.catchup_reservation_n_isrc1__21_ , \catchup.catchup_reservation_n_isrc1__20_ , \catchup.catchup_reservation_n_isrc1__19_ , \catchup.catchup_reservation_n_isrc1__18_ , \catchup.catchup_reservation_n_isrc1__17_ , \catchup.catchup_reservation_n_isrc1__16_ , \catchup.catchup_reservation_n_isrc1__15_ , \catchup.catchup_reservation_n_isrc1__14_ , \catchup.catchup_reservation_n_isrc1__13_ , \catchup.catchup_reservation_n_isrc1__12_ , \catchup.catchup_reservation_n_isrc1__11_ , \catchup.catchup_reservation_n_isrc1__10_ , \catchup.catchup_reservation_n_isrc1__9_ , \catchup.catchup_reservation_n_isrc1__8_ , \catchup.catchup_reservation_n_isrc1__7_ , \catchup.catchup_reservation_n_isrc1__6_ , \catchup.catchup_reservation_n_isrc1__5_ , \catchup.catchup_reservation_n_isrc1__4_ , \catchup.catchup_reservation_n_isrc1__3_ , \catchup.catchup_reservation_n_isrc1__2_ , \catchup.catchup_reservation_n_isrc1__1_ , \catchup.catchup_reservation_n_isrc1__0_ , \catchup.catchup_reservation_n_isrc2__64_ , \catchup.catchup_reservation_n_isrc2__63_ , \catchup.catchup_reservation_n_isrc2__62_ , \catchup.catchup_reservation_n_isrc2__61_ , \catchup.catchup_reservation_n_isrc2__60_ , \catchup.catchup_reservation_n_isrc2__59_ , \catchup.catchup_reservation_n_isrc2__58_ , \catchup.catchup_reservation_n_isrc2__57_ , \catchup.catchup_reservation_n_isrc2__56_ , \catchup.catchup_reservation_n_isrc2__55_ , \catchup.catchup_reservation_n_isrc2__54_ , \catchup.catchup_reservation_n_isrc2__53_ , \catchup.catchup_reservation_n_isrc2__52_ , \catchup.catchup_reservation_n_isrc2__51_ , \catchup.catchup_reservation_n_isrc2__50_ , \catchup.catchup_reservation_n_isrc2__49_ , \catchup.catchup_reservation_n_isrc2__48_ , \catchup.catchup_reservation_n_isrc2__47_ , \catchup.catchup_reservation_n_isrc2__46_ , \catchup.catchup_reservation_n_isrc2__45_ , \catchup.catchup_reservation_n_isrc2__44_ , \catchup.catchup_reservation_n_isrc2__43_ , \catchup.catchup_reservation_n_isrc2__42_ , \catchup.catchup_reservation_n_isrc2__41_ , \catchup.catchup_reservation_n_isrc2__40_ , \catchup.catchup_reservation_n_isrc2__39_ , \catchup.catchup_reservation_n_isrc2__38_ , \catchup.catchup_reservation_n_isrc2__37_ , \catchup.catchup_reservation_n_isrc2__36_ , \catchup.catchup_reservation_n_isrc2__35_ , \catchup.catchup_reservation_n_isrc2__34_ , \catchup.catchup_reservation_n_isrc2__33_ , \catchup.catchup_reservation_n_isrc2__32_ , \catchup.catchup_reservation_n_isrc2__31_ , \catchup.catchup_reservation_n_isrc2__30_ , \catchup.catchup_reservation_n_isrc2__29_ , \catchup.catchup_reservation_n_isrc2__28_ , \catchup.catchup_reservation_n_isrc2__27_ , \catchup.catchup_reservation_n_isrc2__26_ , \catchup.catchup_reservation_n_isrc2__25_ , \catchup.catchup_reservation_n_isrc2__24_ , \catchup.catchup_reservation_n_isrc2__23_ , \catchup.catchup_reservation_n_isrc2__22_ , \catchup.catchup_reservation_n_isrc2__21_ , \catchup.catchup_reservation_n_isrc2__20_ , \catchup.catchup_reservation_n_isrc2__19_ , \catchup.catchup_reservation_n_isrc2__18_ , \catchup.catchup_reservation_n_isrc2__17_ , \catchup.catchup_reservation_n_isrc2__16_ , \catchup.catchup_reservation_n_isrc2__15_ , \catchup.catchup_reservation_n_isrc2__14_ , \catchup.catchup_reservation_n_isrc2__13_ , \catchup.catchup_reservation_n_isrc2__12_ , \catchup.catchup_reservation_n_isrc2__11_ , \catchup.catchup_reservation_n_isrc2__10_ , \catchup.catchup_reservation_n_isrc2__9_ , \catchup.catchup_reservation_n_isrc2__8_ , \catchup.catchup_reservation_n_isrc2__7_ , \catchup.catchup_reservation_n_isrc2__6_ , \catchup.catchup_reservation_n_isrc2__5_ , \catchup.catchup_reservation_n_isrc2__4_ , \catchup.catchup_reservation_n_isrc2__3_ , \catchup.catchup_reservation_n_isrc2__2_ , \catchup.catchup_reservation_n_isrc2__1_ , \catchup.catchup_reservation_n_isrc2__0_ , reservation_r[259:0] }),
    .data_o(\catchup.catchup_reservation_r )
  );


  bp_be_pipe_int_00
  \catchup.pipe_int_catchup 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(exc_stage_n_2__ispec_v_),
    .reservation_i(\catchup.catchup_reservation_r ),
    .flush_i(commit_pkt_o[213]),
    .data_o(pipe_int_catchup_data_lo),
    .v_o(pipe_int_catchup_data_v_lo),
    .branch_o(pipe_int_catchup_branch_lo),
    .btaken_o(pipe_int_catchup_btaken_lo),
    .npc_o(pipe_int_catchup_npc_lo),
    .instr_misaligned_v_o(pipe_int_catchup_instr_misaligned_lo)
  );

  assign N50 = pipe_int_catchup_npc_lo != reservation_r[519:481];

  bp_be_pipe_aux_00
  pipe_aux
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .reservation_i(reservation_r),
    .flush_i(commit_pkt_o[213]),
    .frm_dyn_i(frm_dyn_lo),
    .data_o(pipe_aux_data_lo),
    .v_o(pipe_aux_data_v_lo),
    .fflags_o_nv_(pipe_aux_fflags_lo_nv_),
    .fflags_o_dz_(pipe_aux_fflags_lo_dz_),
    .fflags_o_of_(pipe_aux_fflags_lo_of_),
    .fflags_o_uf_(pipe_aux_fflags_lo_uf_),
    .fflags_o_nx_(pipe_aux_fflags_lo_nx_)
  );


  bp_be_pipe_mem_00
  pipe_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .cfg_bus_i(cfg_bus_i),
    .flush_i(commit_pkt_o[213]),
    .sfence_i(commit_pkt_o[12]),
    .busy_o(mem_busy_o),
    .ordered_o(mem_ordered_o),
    .reservation_i(reservation_r),
    .rs2_val_i(rs2_val_r),
    .commit_pkt_i(commit_pkt_o),
    .tlb_load_miss_v_o(pipe_mem_dtlb_load_miss_lo),
    .tlb_store_miss_v_o(pipe_mem_dtlb_store_miss_lo),
    .cache_miss_v_o(pipe_mem_dcache_miss_lo),
    .cache_replay_v_o(pipe_mem_dcache_replay_lo),
    .load_misaligned_v_o(pipe_mem_load_misaligned_lo),
    .load_access_fault_v_o(pipe_mem_load_access_fault_lo),
    .load_page_fault_v_o(pipe_mem_load_page_fault_lo),
    .store_misaligned_v_o(pipe_mem_store_misaligned_lo),
    .store_access_fault_v_o(pipe_mem_store_access_fault_lo),
    .store_page_fault_v_o(pipe_mem_store_page_fault_lo),
    .early_data_o(pipe_mem_early_data_lo),
    .early_v_o(pipe_mem_early_data_v_lo),
    .final_data_o(pipe_mem_final_data_lo),
    .final_v_o(pipe_mem_final_data_v_lo),
    .late_wb_pkt_o(pipe_mem_late_wb_pkt),
    .late_wb_v_o(late_wb_force_o),
    .trans_info_i(trans_info_o),
    .cache_req_o(cache_req_o),
    .cache_req_v_o(cache_req_v_o),
    .cache_req_yumi_i(cache_req_yumi_i),
    .cache_req_lock_i(cache_req_lock_i),
    .cache_req_metadata_o(cache_req_metadata_o),
    .cache_req_metadata_v_o(cache_req_metadata_v_o),
    .cache_req_id_i(cache_req_id_i[0]),
    .cache_req_critical_i(cache_req_critical_i),
    .cache_req_last_i(cache_req_last_i),
    .cache_req_credits_full_i(cache_req_credits_full_i),
    .cache_req_credits_empty_i(cache_req_credits_empty_i),
    .data_mem_pkt_v_i(data_mem_pkt_v_i),
    .data_mem_pkt_i(data_mem_pkt_i),
    .data_mem_pkt_yumi_o(data_mem_pkt_yumi_o),
    .data_mem_o(data_mem_o),
    .tag_mem_pkt_v_i(tag_mem_pkt_v_i),
    .tag_mem_pkt_i(tag_mem_pkt_i),
    .tag_mem_pkt_yumi_o(tag_mem_pkt_yumi_o),
    .tag_mem_o(tag_mem_o),
    .stat_mem_pkt_v_i(stat_mem_pkt_v_i),
    .stat_mem_pkt_i(stat_mem_pkt_i),
    .stat_mem_pkt_yumi_o(stat_mem_pkt_yumi_o),
    .stat_mem_o(stat_mem_o)
  );


  bp_be_pipe_fma_00
  pipe_fma
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .reservation_i(reservation_r),
    .flush_i(commit_pkt_o[213]),
    .frm_dyn_i(frm_dyn_lo),
    .imul_data_o(pipe_mul_data_lo),
    .imul_v_o(pipe_mul_data_v_lo),
    .fma_data_o(pipe_fma_data_lo),
    .fma_v_o(pipe_fma_data_v_lo),
    .fma_fflags_o_nv_(pipe_fma_fflags_lo_nv_),
    .fma_fflags_o_dz_(pipe_fma_fflags_lo_dz_),
    .fma_fflags_o_of_(pipe_fma_fflags_lo_of_),
    .fma_fflags_o_uf_(pipe_fma_fflags_lo_uf_),
    .fma_fflags_o_nx_(pipe_fma_fflags_lo_nx_)
  );


  bp_be_pipe_long_00
  pipe_long
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .reservation_i(reservation_r),
    .ibusy_o(idiv_busy_o),
    .fbusy_o(fdiv_busy_o),
    .frm_dyn_i(frm_dyn_lo),
    .flush_i(commit_pkt_o[213]),
    .iwb_pkt_o(pipe_long_iwb_pkt),
    .iwb_v_o(late_wb_reqs_li[1]),
    .iwb_yumi_i(pipe_long_idata_yumi_lo),
    .fwb_pkt_o(pipe_long_fwb_pkt),
    .fwb_v_o(late_wb_reqs_li[2]),
    .fwb_yumi_i(pipe_long_fdata_yumi_lo)
  );


  bsg_arb_fixed_inputs_p3_lo_to_hi_p1
  late_wb_arb
  (
    .ready_then_i(1'b1),
    .reqs_i({ late_wb_reqs_li, late_wb_force_o }),
    .grants_o(late_wb_grants_lo)
  );


  bsg_mux_one_hot_width_p79_els_p3
  late_wb_mux_oh
  (
    .data_i({ pipe_long_fwb_pkt, pipe_long_iwb_pkt, pipe_mem_late_wb_pkt }),
    .sel_one_hot_i(late_wb_grants_lo),
    .data_o(late_wb_pkt_o)
  );


  bsg_dff_width_p395
  comp_stage_reg
  (
    .clk_i(clk_i),
    .data_i({ comp_stage_n_4__ird_w_v_, comp_stage_n_4__frd_w_v_, iwb_pkt_o[76:71], forward_data_3__65_, forward_data_3__64_, forward_data_3__63_, forward_data_3__62_, forward_data_3__61_, forward_data_3__60_, forward_data_3__59_, forward_data_3__58_, forward_data_3__57_, forward_data_3__56_, forward_data_3__55_, forward_data_3__54_, forward_data_3__53_, forward_data_3__52_, forward_data_3__51_, forward_data_3__50_, forward_data_3__49_, forward_data_3__48_, forward_data_3__47_, forward_data_3__46_, forward_data_3__45_, forward_data_3__44_, forward_data_3__43_, forward_data_3__42_, forward_data_3__41_, forward_data_3__40_, forward_data_3__39_, forward_data_3__38_, forward_data_3__37_, forward_data_3__36_, forward_data_3__35_, forward_data_3__34_, forward_data_3__33_, forward_data_3__32_, forward_data_3__31_, forward_data_3__30_, forward_data_3__29_, forward_data_3__28_, forward_data_3__27_, forward_data_3__26_, forward_data_3__25_, forward_data_3__24_, forward_data_3__23_, forward_data_3__22_, forward_data_3__21_, forward_data_3__20_, forward_data_3__19_, forward_data_3__18_, forward_data_3__17_, forward_data_3__16_, forward_data_3__15_, forward_data_3__14_, forward_data_3__13_, forward_data_3__12_, forward_data_3__11_, forward_data_3__10_, forward_data_3__9_, forward_data_3__8_, forward_data_3__7_, forward_data_3__6_, forward_data_3__5_, forward_data_3__4_, forward_data_3__3_, forward_data_3__2_, forward_data_3__1_, forward_data_3__0_, comp_stage_n_4__fflags__nv_, comp_stage_n_4__fflags__dz_, comp_stage_n_4__fflags__of_, comp_stage_n_4__fflags__uf_, comp_stage_n_4__fflags__nx_, comp_stage_n_3__ird_w_v_, comp_stage_n_3__frd_w_v_, comp_stage_n_3__ptw_w_v_, comp_stage_n_3__rd_addr__4_, comp_stage_n_3__rd_addr__3_, comp_stage_n_3__rd_addr__2_, comp_stage_n_3__rd_addr__1_, comp_stage_n_3__rd_addr__0_, forward_data_2__65_, forward_data_2__64_, forward_data_2__63_, forward_data_2__62_, forward_data_2__61_, forward_data_2__60_, forward_data_2__59_, forward_data_2__58_, forward_data_2__57_, forward_data_2__56_, forward_data_2__55_, forward_data_2__54_, forward_data_2__53_, forward_data_2__52_, forward_data_2__51_, forward_data_2__50_, forward_data_2__49_, forward_data_2__48_, forward_data_2__47_, forward_data_2__46_, forward_data_2__45_, forward_data_2__44_, forward_data_2__43_, forward_data_2__42_, forward_data_2__41_, forward_data_2__40_, forward_data_2__39_, forward_data_2__38_, forward_data_2__37_, forward_data_2__36_, forward_data_2__35_, forward_data_2__34_, forward_data_2__33_, forward_data_2__32_, forward_data_2__31_, forward_data_2__30_, forward_data_2__29_, forward_data_2__28_, forward_data_2__27_, forward_data_2__26_, forward_data_2__25_, forward_data_2__24_, forward_data_2__23_, forward_data_2__22_, forward_data_2__21_, forward_data_2__20_, forward_data_2__19_, forward_data_2__18_, forward_data_2__17_, forward_data_2__16_, forward_data_2__15_, forward_data_2__14_, forward_data_2__13_, forward_data_2__12_, forward_data_2__11_, forward_data_2__10_, forward_data_2__9_, forward_data_2__8_, forward_data_2__7_, forward_data_2__6_, forward_data_2__5_, forward_data_2__4_, forward_data_2__3_, forward_data_2__2_, forward_data_2__1_, forward_data_2__0_, comp_stage_n_3__fflags__nv_, comp_stage_n_3__fflags__dz_, comp_stage_n_3__fflags__of_, comp_stage_n_3__fflags__uf_, comp_stage_n_3__fflags__nx_, comp_stage_n_2__ird_w_v_, comp_stage_n_2__frd_w_v_, comp_stage_n_2__ptw_w_v_, comp_stage_n_2__rd_addr__4_, comp_stage_n_2__rd_addr__3_, comp_stage_n_2__rd_addr__2_, comp_stage_n_2__rd_addr__1_, comp_stage_n_2__rd_addr__0_, forward_data_1__65_, forward_data_1__64_, forward_data_1__63_, forward_data_1__62_, forward_data_1__61_, forward_data_1__60_, forward_data_1__59_, forward_data_1__58_, forward_data_1__57_, forward_data_1__56_, forward_data_1__55_, forward_data_1__54_, forward_data_1__53_, forward_data_1__52_, forward_data_1__51_, forward_data_1__50_, forward_data_1__49_, forward_data_1__48_, forward_data_1__47_, forward_data_1__46_, forward_data_1__45_, forward_data_1__44_, forward_data_1__43_, forward_data_1__42_, forward_data_1__41_, forward_data_1__40_, forward_data_1__39_, forward_data_1__38_, forward_data_1__37_, forward_data_1__36_, forward_data_1__35_, forward_data_1__34_, forward_data_1__33_, forward_data_1__32_, forward_data_1__31_, forward_data_1__30_, forward_data_1__29_, forward_data_1__28_, forward_data_1__27_, forward_data_1__26_, forward_data_1__25_, forward_data_1__24_, forward_data_1__23_, forward_data_1__22_, forward_data_1__21_, forward_data_1__20_, forward_data_1__19_, forward_data_1__18_, forward_data_1__17_, forward_data_1__16_, forward_data_1__15_, forward_data_1__14_, forward_data_1__13_, forward_data_1__12_, forward_data_1__11_, forward_data_1__10_, forward_data_1__9_, forward_data_1__8_, forward_data_1__7_, forward_data_1__6_, forward_data_1__5_, forward_data_1__4_, forward_data_1__3_, forward_data_1__2_, forward_data_1__1_, forward_data_1__0_, comp_stage_n_2__fflags__nv_, comp_stage_n_2__fflags__dz_, comp_stage_n_2__fflags__of_, comp_stage_n_2__fflags__uf_, comp_stage_n_2__fflags__nx_, comp_stage_n_1__ird_w_v_, comp_stage_n_1__frd_w_v_, comp_stage_n_1__ptw_w_v_, comp_stage_n_1__rd_addr__4_, comp_stage_n_1__rd_addr__3_, comp_stage_n_1__rd_addr__2_, comp_stage_n_1__rd_addr__1_, comp_stage_n_1__rd_addr__0_, forward_data_0__65_, forward_data_0__64_, forward_data_0__63_, forward_data_0__62_, forward_data_0__61_, forward_data_0__60_, forward_data_0__59_, forward_data_0__58_, forward_data_0__57_, forward_data_0__56_, forward_data_0__55_, forward_data_0__54_, forward_data_0__53_, forward_data_0__52_, forward_data_0__51_, forward_data_0__50_, forward_data_0__49_, forward_data_0__48_, forward_data_0__47_, forward_data_0__46_, forward_data_0__45_, forward_data_0__44_, forward_data_0__43_, forward_data_0__42_, forward_data_0__41_, forward_data_0__40_, forward_data_0__39_, forward_data_0__38_, forward_data_0__37_, forward_data_0__36_, forward_data_0__35_, forward_data_0__34_, forward_data_0__33_, forward_data_0__32_, forward_data_0__31_, forward_data_0__30_, forward_data_0__29_, forward_data_0__28_, forward_data_0__27_, forward_data_0__26_, forward_data_0__25_, forward_data_0__24_, forward_data_0__23_, forward_data_0__22_, forward_data_0__21_, forward_data_0__20_, forward_data_0__19_, forward_data_0__18_, forward_data_0__17_, forward_data_0__16_, forward_data_0__15_, forward_data_0__14_, forward_data_0__13_, forward_data_0__12_, forward_data_0__11_, forward_data_0__10_, forward_data_0__9_, forward_data_0__8_, forward_data_0__7_, forward_data_0__6_, forward_data_0__5_, forward_data_0__4_, forward_data_0__3_, forward_data_0__2_, forward_data_0__1_, forward_data_0__0_, comp_stage_n_1__fflags__nv_, comp_stage_n_1__fflags__dz_, comp_stage_n_1__fflags__of_, comp_stage_n_1__fflags__uf_, comp_stage_n_1__fflags__nx_, comp_stage_n_0__ird_w_v_, comp_stage_n_0__frd_w_v_, 1'b0, dispatch_pkt_i[302:298], comp_stage_n_0__rd_data__65_, comp_stage_n_0__rd_data__64_, comp_stage_n_0__rd_data__63_, comp_stage_n_0__rd_data__62_, comp_stage_n_0__rd_data__61_, comp_stage_n_0__rd_data__60_, comp_stage_n_0__rd_data__59_, comp_stage_n_0__rd_data__58_, comp_stage_n_0__rd_data__57_, comp_stage_n_0__rd_data__56_, comp_stage_n_0__rd_data__55_, comp_stage_n_0__rd_data__54_, comp_stage_n_0__rd_data__53_, comp_stage_n_0__rd_data__52_, comp_stage_n_0__rd_data__51_, comp_stage_n_0__rd_data__50_, comp_stage_n_0__rd_data__49_, comp_stage_n_0__rd_data__48_, comp_stage_n_0__rd_data__47_, comp_stage_n_0__rd_data__46_, comp_stage_n_0__rd_data__45_, comp_stage_n_0__rd_data__44_, comp_stage_n_0__rd_data__43_, comp_stage_n_0__rd_data__42_, comp_stage_n_0__rd_data__41_, comp_stage_n_0__rd_data__40_, comp_stage_n_0__rd_data__39_, comp_stage_n_0__rd_data__38_, comp_stage_n_0__rd_data__37_, comp_stage_n_0__rd_data__36_, comp_stage_n_0__rd_data__35_, comp_stage_n_0__rd_data__34_, comp_stage_n_0__rd_data__33_, comp_stage_n_0__rd_data__32_, comp_stage_n_0__rd_data__31_, comp_stage_n_0__rd_data__30_, comp_stage_n_0__rd_data__29_, comp_stage_n_0__rd_data__28_, comp_stage_n_0__rd_data__27_, comp_stage_n_0__rd_data__26_, comp_stage_n_0__rd_data__25_, comp_stage_n_0__rd_data__24_, comp_stage_n_0__rd_data__23_, comp_stage_n_0__rd_data__22_, comp_stage_n_0__rd_data__21_, comp_stage_n_0__rd_data__20_, comp_stage_n_0__rd_data__19_, comp_stage_n_0__rd_data__18_, comp_stage_n_0__rd_data__17_, comp_stage_n_0__rd_data__16_, comp_stage_n_0__rd_data__15_, comp_stage_n_0__rd_data__14_, comp_stage_n_0__rd_data__13_, comp_stage_n_0__rd_data__12_, comp_stage_n_0__rd_data__11_, comp_stage_n_0__rd_data__10_, comp_stage_n_0__rd_data__9_, comp_stage_n_0__rd_data__8_, comp_stage_n_0__rd_data__7_, comp_stage_n_0__rd_data__6_, comp_stage_n_0__rd_data__5_, comp_stage_n_0__rd_data__4_, comp_stage_n_0__rd_data__3_, comp_stage_n_0__rd_data__2_, comp_stage_n_0__rd_data__1_, comp_stage_n_0__rd_data__0_, comp_stage_n_0__fflags__nv_, comp_stage_n_0__fflags__dz_, comp_stage_n_0__fflags__of_, comp_stage_n_0__fflags__uf_, comp_stage_n_0__fflags__nx_ }),
    .data_o({ fwb_pkt_o, iwb_pkt_o, comp_stage_r_2__ird_w_v_, comp_stage_r_2__frd_w_v_, comp_stage_n_3__ptw_w_v_, comp_stage_n_3__rd_addr__4_, comp_stage_n_3__rd_addr__3_, comp_stage_n_3__rd_addr__2_, comp_stage_n_3__rd_addr__1_, comp_stage_n_3__rd_addr__0_, comp_stage_r_2__rd_data__65_, comp_stage_r_2__rd_data__64_, comp_stage_r_2__rd_data__63_, comp_stage_r_2__rd_data__62_, comp_stage_r_2__rd_data__61_, comp_stage_r_2__rd_data__60_, comp_stage_r_2__rd_data__59_, comp_stage_r_2__rd_data__58_, comp_stage_r_2__rd_data__57_, comp_stage_r_2__rd_data__56_, comp_stage_r_2__rd_data__55_, comp_stage_r_2__rd_data__54_, comp_stage_r_2__rd_data__53_, comp_stage_r_2__rd_data__52_, comp_stage_r_2__rd_data__51_, comp_stage_r_2__rd_data__50_, comp_stage_r_2__rd_data__49_, comp_stage_r_2__rd_data__48_, comp_stage_r_2__rd_data__47_, comp_stage_r_2__rd_data__46_, comp_stage_r_2__rd_data__45_, comp_stage_r_2__rd_data__44_, comp_stage_r_2__rd_data__43_, comp_stage_r_2__rd_data__42_, comp_stage_r_2__rd_data__41_, comp_stage_r_2__rd_data__40_, comp_stage_r_2__rd_data__39_, comp_stage_r_2__rd_data__38_, comp_stage_r_2__rd_data__37_, comp_stage_r_2__rd_data__36_, comp_stage_r_2__rd_data__35_, comp_stage_r_2__rd_data__34_, comp_stage_r_2__rd_data__33_, comp_stage_r_2__rd_data__32_, comp_stage_r_2__rd_data__31_, comp_stage_r_2__rd_data__30_, comp_stage_r_2__rd_data__29_, comp_stage_r_2__rd_data__28_, comp_stage_r_2__rd_data__27_, comp_stage_r_2__rd_data__26_, comp_stage_r_2__rd_data__25_, comp_stage_r_2__rd_data__24_, comp_stage_r_2__rd_data__23_, comp_stage_r_2__rd_data__22_, comp_stage_r_2__rd_data__21_, comp_stage_r_2__rd_data__20_, comp_stage_r_2__rd_data__19_, comp_stage_r_2__rd_data__18_, comp_stage_r_2__rd_data__17_, comp_stage_r_2__rd_data__16_, comp_stage_r_2__rd_data__15_, comp_stage_r_2__rd_data__14_, comp_stage_r_2__rd_data__13_, comp_stage_r_2__rd_data__12_, comp_stage_r_2__rd_data__11_, comp_stage_r_2__rd_data__10_, comp_stage_r_2__rd_data__9_, comp_stage_r_2__rd_data__8_, comp_stage_r_2__rd_data__7_, comp_stage_r_2__rd_data__6_, comp_stage_r_2__rd_data__5_, comp_stage_r_2__rd_data__4_, comp_stage_r_2__rd_data__3_, comp_stage_r_2__rd_data__2_, comp_stage_r_2__rd_data__1_, comp_stage_r_2__rd_data__0_, comp_stage_r_2__fflags__nv_, comp_stage_r_2__fflags__dz_, comp_stage_r_2__fflags__of_, comp_stage_r_2__fflags__uf_, comp_stage_r_2__fflags__nx_, comp_stage_r_1__ird_w_v_, comp_stage_r_1__frd_w_v_, comp_stage_n_2__ptw_w_v_, comp_stage_n_2__rd_addr__4_, comp_stage_n_2__rd_addr__3_, comp_stage_n_2__rd_addr__2_, comp_stage_n_2__rd_addr__1_, comp_stage_n_2__rd_addr__0_, comp_stage_r_1__rd_data__65_, comp_stage_r_1__rd_data__64_, comp_stage_r_1__rd_data__63_, comp_stage_r_1__rd_data__62_, comp_stage_r_1__rd_data__61_, comp_stage_r_1__rd_data__60_, comp_stage_r_1__rd_data__59_, comp_stage_r_1__rd_data__58_, comp_stage_r_1__rd_data__57_, comp_stage_r_1__rd_data__56_, comp_stage_r_1__rd_data__55_, comp_stage_r_1__rd_data__54_, comp_stage_r_1__rd_data__53_, comp_stage_r_1__rd_data__52_, comp_stage_r_1__rd_data__51_, comp_stage_r_1__rd_data__50_, comp_stage_r_1__rd_data__49_, comp_stage_r_1__rd_data__48_, comp_stage_r_1__rd_data__47_, comp_stage_r_1__rd_data__46_, comp_stage_r_1__rd_data__45_, comp_stage_r_1__rd_data__44_, comp_stage_r_1__rd_data__43_, comp_stage_r_1__rd_data__42_, comp_stage_r_1__rd_data__41_, comp_stage_r_1__rd_data__40_, comp_stage_r_1__rd_data__39_, comp_stage_r_1__rd_data__38_, comp_stage_r_1__rd_data__37_, comp_stage_r_1__rd_data__36_, comp_stage_r_1__rd_data__35_, comp_stage_r_1__rd_data__34_, comp_stage_r_1__rd_data__33_, comp_stage_r_1__rd_data__32_, comp_stage_r_1__rd_data__31_, comp_stage_r_1__rd_data__30_, comp_stage_r_1__rd_data__29_, comp_stage_r_1__rd_data__28_, comp_stage_r_1__rd_data__27_, comp_stage_r_1__rd_data__26_, comp_stage_r_1__rd_data__25_, comp_stage_r_1__rd_data__24_, comp_stage_r_1__rd_data__23_, comp_stage_r_1__rd_data__22_, comp_stage_r_1__rd_data__21_, comp_stage_r_1__rd_data__20_, comp_stage_r_1__rd_data__19_, comp_stage_r_1__rd_data__18_, comp_stage_r_1__rd_data__17_, comp_stage_r_1__rd_data__16_, comp_stage_r_1__rd_data__15_, comp_stage_r_1__rd_data__14_, comp_stage_r_1__rd_data__13_, comp_stage_r_1__rd_data__12_, comp_stage_r_1__rd_data__11_, comp_stage_r_1__rd_data__10_, comp_stage_r_1__rd_data__9_, comp_stage_r_1__rd_data__8_, comp_stage_r_1__rd_data__7_, comp_stage_r_1__rd_data__6_, comp_stage_r_1__rd_data__5_, comp_stage_r_1__rd_data__4_, comp_stage_r_1__rd_data__3_, comp_stage_r_1__rd_data__2_, comp_stage_r_1__rd_data__1_, comp_stage_r_1__rd_data__0_, comp_stage_r_1__fflags__nv_, comp_stage_r_1__fflags__dz_, comp_stage_r_1__fflags__of_, comp_stage_r_1__fflags__uf_, comp_stage_r_1__fflags__nx_, comp_stage_r_0__ird_w_v_, comp_stage_r_0__frd_w_v_, comp_stage_n_1__ptw_w_v_, comp_stage_n_1__rd_addr__4_, comp_stage_n_1__rd_addr__3_, comp_stage_n_1__rd_addr__2_, comp_stage_n_1__rd_addr__1_, comp_stage_n_1__rd_addr__0_, comp_stage_r_0__rd_data__65_, comp_stage_r_0__rd_data__64_, comp_stage_r_0__rd_data__63_, comp_stage_r_0__rd_data__62_, comp_stage_r_0__rd_data__61_, comp_stage_r_0__rd_data__60_, comp_stage_r_0__rd_data__59_, comp_stage_r_0__rd_data__58_, comp_stage_r_0__rd_data__57_, comp_stage_r_0__rd_data__56_, comp_stage_r_0__rd_data__55_, comp_stage_r_0__rd_data__54_, comp_stage_r_0__rd_data__53_, comp_stage_r_0__rd_data__52_, comp_stage_r_0__rd_data__51_, comp_stage_r_0__rd_data__50_, comp_stage_r_0__rd_data__49_, comp_stage_r_0__rd_data__48_, comp_stage_r_0__rd_data__47_, comp_stage_r_0__rd_data__46_, comp_stage_r_0__rd_data__45_, comp_stage_r_0__rd_data__44_, comp_stage_r_0__rd_data__43_, comp_stage_r_0__rd_data__42_, comp_stage_r_0__rd_data__41_, comp_stage_r_0__rd_data__40_, comp_stage_r_0__rd_data__39_, comp_stage_r_0__rd_data__38_, comp_stage_r_0__rd_data__37_, comp_stage_r_0__rd_data__36_, comp_stage_r_0__rd_data__35_, comp_stage_r_0__rd_data__34_, comp_stage_r_0__rd_data__33_, comp_stage_r_0__rd_data__32_, comp_stage_r_0__rd_data__31_, comp_stage_r_0__rd_data__30_, comp_stage_r_0__rd_data__29_, comp_stage_r_0__rd_data__28_, comp_stage_r_0__rd_data__27_, comp_stage_r_0__rd_data__26_, comp_stage_r_0__rd_data__25_, comp_stage_r_0__rd_data__24_, comp_stage_r_0__rd_data__23_, comp_stage_r_0__rd_data__22_, comp_stage_r_0__rd_data__21_, comp_stage_r_0__rd_data__20_, comp_stage_r_0__rd_data__19_, comp_stage_r_0__rd_data__18_, comp_stage_r_0__rd_data__17_, comp_stage_r_0__rd_data__16_, comp_stage_r_0__rd_data__15_, comp_stage_r_0__rd_data__14_, comp_stage_r_0__rd_data__13_, comp_stage_r_0__rd_data__12_, comp_stage_r_0__rd_data__11_, comp_stage_r_0__rd_data__10_, comp_stage_r_0__rd_data__9_, comp_stage_r_0__rd_data__8_, comp_stage_r_0__rd_data__7_, comp_stage_r_0__rd_data__6_, comp_stage_r_0__rd_data__5_, comp_stage_r_0__rd_data__4_, comp_stage_r_0__rd_data__3_, comp_stage_r_0__rd_data__2_, comp_stage_r_0__rd_data__1_, comp_stage_r_0__rd_data__0_, comp_stage_r_0__fflags__nv_, comp_stage_r_0__fflags__dz_, comp_stage_r_0__fflags__of_, comp_stage_r_0__fflags__uf_, comp_stage_r_0__fflags__nx_ })
  );


  bsg_dff_width_p190
  exc_stage_reg
  (
    .clk_i(clk_i),
    .data_i({ exc_stage_n_4__v_, exc_stage_n_4__queue_v_, exc_stage_n_4__ispec_v_, exc_stage_n_4__nspec_v_, exc_stage_n_4__exc__store_page_fault_, exc_stage_n_4__exc__load_page_fault_, exc_stage_n_4__exc__instr_page_fault_, exc_stage_n_4__exc__ecall_m_, exc_stage_n_4__exc__ecall_s_, exc_stage_n_4__exc__ecall_u_, exc_stage_n_4__exc__store_access_fault_, exc_stage_n_4__exc__store_misaligned_, exc_stage_n_4__exc__load_access_fault_, exc_stage_n_4__exc__load_misaligned_, exc_stage_n_4__exc__ebreak_, exc_stage_n_4__exc__illegal_instr_, exc_stage_n_4__exc__instr_access_fault_, exc_stage_n_4__exc__instr_misaligned_, exc_stage_n_4__exc__resume_, exc_stage_n_4__exc__itlb_miss_, exc_stage_n_4__exc__icache_miss_, exc_stage_n_4__exc__dcache_replay_, exc_stage_n_4__exc__dtlb_load_miss_, exc_stage_n_4__exc__dtlb_store_miss_, exc_stage_n_4__exc__itlb_fill_, exc_stage_n_4__exc__dtlb_fill_, exc_stage_n_4__exc___interrupt_, exc_stage_n_4__exc__cmd_full_, exc_stage_n_4__exc__mispredict_, exc_stage_n_4__spec__dcache_miss_, exc_stage_n_4__spec__fencei_, exc_stage_n_4__spec__sfence_vma_, exc_stage_n_4__spec__dbreak_, exc_stage_n_4__spec__dret_, exc_stage_n_4__spec__mret_, exc_stage_n_4__spec__sret_, exc_stage_n_4__spec__wfi_, exc_stage_n_4__spec__csrw_, exc_stage_n_3__v_, exc_stage_n_3__queue_v_, exc_stage_n_3__ispec_v_, exc_stage_n_3__nspec_v_, exc_stage_n_3__exc__store_page_fault_, exc_stage_n_3__exc__load_page_fault_, exc_stage_n_3__exc__instr_page_fault_, exc_stage_n_3__exc__ecall_m_, exc_stage_n_3__exc__ecall_s_, exc_stage_n_3__exc__ecall_u_, exc_stage_n_3__exc__store_access_fault_, exc_stage_n_3__exc__store_misaligned_, exc_stage_n_3__exc__load_access_fault_, exc_stage_n_3__exc__load_misaligned_, exc_stage_n_3__exc__ebreak_, exc_stage_n_3__exc__illegal_instr_, exc_stage_n_3__exc__instr_access_fault_, exc_stage_n_3__exc__instr_misaligned_, exc_stage_n_3__exc__resume_, exc_stage_n_3__exc__itlb_miss_, exc_stage_n_3__exc__icache_miss_, exc_stage_n_3__exc__dcache_replay_, exc_stage_n_3__exc__dtlb_load_miss_, exc_stage_n_3__exc__dtlb_store_miss_, exc_stage_n_3__exc__itlb_fill_, exc_stage_n_3__exc__dtlb_fill_, exc_stage_n_3__exc___interrupt_, exc_stage_n_3__exc__cmd_full_, exc_stage_n_3__exc__mispredict_, exc_stage_n_3__spec__dcache_miss_, exc_stage_n_3__spec__fencei_, exc_stage_n_3__spec__sfence_vma_, exc_stage_n_3__spec__dbreak_, exc_stage_n_3__spec__dret_, exc_stage_n_3__spec__mret_, exc_stage_n_3__spec__sret_, exc_stage_n_3__spec__wfi_, exc_stage_n_3__spec__csrw_, exc_stage_n_2__v_, exc_stage_n_2__queue_v_, exc_stage_n_2__ispec_v_, exc_stage_n_2__nspec_v_, exc_stage_n_2__exc__store_page_fault_, exc_stage_n_2__exc__load_page_fault_, exc_stage_n_2__exc__instr_page_fault_, exc_stage_n_2__exc__ecall_m_, exc_stage_n_2__exc__ecall_s_, exc_stage_n_2__exc__ecall_u_, exc_stage_n_2__exc__store_access_fault_, exc_stage_n_2__exc__store_misaligned_, exc_stage_n_2__exc__load_access_fault_, exc_stage_n_2__exc__load_misaligned_, exc_stage_n_2__exc__ebreak_, exc_stage_n_2__exc__illegal_instr_, exc_stage_n_2__exc__instr_access_fault_, exc_stage_n_2__exc__instr_misaligned_, exc_stage_n_2__exc__resume_, exc_stage_n_2__exc__itlb_miss_, exc_stage_n_2__exc__icache_miss_, exc_stage_n_2__exc__dcache_replay_, exc_stage_n_2__exc__dtlb_load_miss_, exc_stage_n_2__exc__dtlb_store_miss_, exc_stage_n_2__exc__itlb_fill_, exc_stage_n_2__exc__dtlb_fill_, exc_stage_n_2__exc___interrupt_, exc_stage_n_2__exc__cmd_full_, exc_stage_n_2__exc__mispredict_, exc_stage_n_2__spec__dcache_miss_, exc_stage_n_2__spec__fencei_, exc_stage_n_2__spec__sfence_vma_, exc_stage_n_2__spec__dbreak_, exc_stage_n_2__spec__dret_, exc_stage_n_2__spec__mret_, exc_stage_n_2__spec__sret_, exc_stage_n_2__spec__wfi_, exc_stage_n_2__spec__csrw_, exc_stage_n_1__v_, exc_stage_n_1__queue_v_, exc_stage_n_1__ispec_v_, exc_stage_n_1__nspec_v_, exc_stage_n_1__exc__store_page_fault_, exc_stage_n_1__exc__load_page_fault_, exc_stage_n_1__exc__instr_page_fault_, exc_stage_n_1__exc__ecall_m_, exc_stage_n_1__exc__ecall_s_, exc_stage_n_1__exc__ecall_u_, exc_stage_n_1__exc__store_access_fault_, exc_stage_n_1__exc__store_misaligned_, exc_stage_n_1__exc__load_access_fault_, exc_stage_n_1__exc__load_misaligned_, exc_stage_n_1__exc__ebreak_, exc_stage_n_1__exc__illegal_instr_, exc_stage_n_1__exc__instr_access_fault_, exc_stage_n_1__exc__instr_misaligned_, exc_stage_n_1__exc__resume_, exc_stage_n_1__exc__itlb_miss_, exc_stage_n_1__exc__icache_miss_, exc_stage_n_1__exc__dcache_replay_, exc_stage_n_1__exc__dtlb_load_miss_, exc_stage_n_1__exc__dtlb_store_miss_, exc_stage_n_1__exc__itlb_fill_, exc_stage_n_1__exc__dtlb_fill_, exc_stage_n_1__exc___interrupt_, exc_stage_n_1__exc__cmd_full_, exc_stage_n_1__exc__mispredict_, exc_stage_n_1__spec__dcache_miss_, exc_stage_n_1__spec__fencei_, exc_stage_n_1__spec__sfence_vma_, exc_stage_n_1__spec__dbreak_, exc_stage_n_1__spec__dret_, exc_stage_n_1__spec__mret_, exc_stage_n_1__spec__sret_, exc_stage_n_1__spec__wfi_, exc_stage_n_1__spec__csrw_, exc_stage_n_0__v_, exc_stage_n_0__queue_v_, dispatch_pkt_i[363:362], dispatch_pkt_i[33:0] }),
    .data_o({ exc_stage_n_5__v_, exc_stage_n_5__queue_v_, exc_stage_n_5__ispec_v_, exc_stage_n_5__nspec_v_, exc_stage_n_5__exc__store_page_fault_, exc_stage_n_5__exc__load_page_fault_, exc_stage_n_5__exc__instr_page_fault_, exc_stage_n_5__exc__ecall_m_, exc_stage_n_5__exc__ecall_s_, exc_stage_n_5__exc__ecall_u_, exc_stage_n_5__exc__store_access_fault_, exc_stage_n_5__exc__store_misaligned_, exc_stage_n_5__exc__load_access_fault_, exc_stage_n_5__exc__load_misaligned_, exc_stage_n_5__exc__ebreak_, exc_stage_n_5__exc__illegal_instr_, exc_stage_n_5__exc__instr_access_fault_, exc_stage_n_5__exc__instr_misaligned_, exc_stage_n_5__exc__resume_, exc_stage_n_5__exc__itlb_miss_, exc_stage_n_5__exc__icache_miss_, exc_stage_n_5__exc__dcache_replay_, exc_stage_n_5__exc__dtlb_load_miss_, exc_stage_n_5__exc__dtlb_store_miss_, exc_stage_n_5__exc__itlb_fill_, exc_stage_n_5__exc__dtlb_fill_, exc_stage_n_5__exc___interrupt_, exc_stage_n_5__exc__cmd_full_, exc_stage_n_5__exc__mispredict_, exc_stage_n_5__spec__dcache_miss_, exc_stage_n_5__spec__fencei_, exc_stage_n_5__spec__sfence_vma_, exc_stage_n_5__spec__dbreak_, exc_stage_n_5__spec__dret_, exc_stage_n_5__spec__mret_, exc_stage_n_5__spec__sret_, exc_stage_n_5__spec__wfi_, exc_stage_n_5__spec__csrw_, exc_stage_n_4__v_, exc_stage_n_4__queue_v_, exc_stage_n_4__ispec_v_, exc_stage_n_4__nspec_v_, exc_stage_n_4__exc__store_page_fault_, exc_stage_n_4__exc__load_page_fault_, exc_stage_n_4__exc__instr_page_fault_, exc_stage_n_4__exc__ecall_m_, exc_stage_n_4__exc__ecall_s_, exc_stage_n_4__exc__ecall_u_, exc_stage_n_4__exc__store_access_fault_, exc_stage_n_4__exc__store_misaligned_, exc_stage_n_4__exc__load_access_fault_, exc_stage_n_4__exc__load_misaligned_, exc_stage_n_4__exc__ebreak_, exc_stage_n_4__exc__illegal_instr_, exc_stage_n_4__exc__instr_access_fault_, exc_stage_n_4__exc__instr_misaligned_, exc_stage_n_4__exc__resume_, exc_stage_n_4__exc__itlb_miss_, exc_stage_n_4__exc__icache_miss_, exc_stage_n_4__exc__dcache_replay_, exc_stage_n_4__exc__dtlb_load_miss_, exc_stage_n_4__exc__dtlb_store_miss_, exc_stage_n_4__exc__itlb_fill_, exc_stage_n_4__exc__dtlb_fill_, exc_stage_n_4__exc___interrupt_, exc_stage_n_4__exc__cmd_full_, exc_stage_n_4__exc__mispredict_, exc_stage_n_4__spec__dcache_miss_, exc_stage_n_4__spec__fencei_, exc_stage_n_4__spec__sfence_vma_, exc_stage_n_4__spec__dbreak_, exc_stage_n_4__spec__dret_, exc_stage_n_4__spec__mret_, exc_stage_n_4__spec__sret_, exc_stage_n_4__spec__wfi_, exc_stage_n_4__spec__csrw_, exc_stage_r_2__v_, exc_stage_n_3__queue_v_, exc_stage_n_3__ispec_v_, exc_stage_n_3__nspec_v_, exc_stage_n_3__exc__store_page_fault_, exc_stage_n_3__exc__load_page_fault_, exc_stage_n_3__exc__instr_page_fault_, exc_stage_n_3__exc__ecall_m_, exc_stage_n_3__exc__ecall_s_, exc_stage_n_3__exc__ecall_u_, exc_stage_n_3__exc__store_access_fault_, exc_stage_n_3__exc__store_misaligned_, exc_stage_n_3__exc__load_access_fault_, exc_stage_n_3__exc__load_misaligned_, exc_stage_n_3__exc__ebreak_, exc_stage_n_3__exc__illegal_instr_, exc_stage_n_3__exc__instr_access_fault_, exc_stage_n_3__exc__instr_misaligned_, exc_stage_n_3__exc__resume_, exc_stage_n_3__exc__itlb_miss_, exc_stage_n_3__exc__icache_miss_, exc_stage_n_3__exc__dcache_replay_, exc_stage_n_3__exc__dtlb_load_miss_, exc_stage_n_3__exc__dtlb_store_miss_, exc_stage_n_3__exc__itlb_fill_, exc_stage_n_3__exc__dtlb_fill_, exc_stage_n_3__exc___interrupt_, exc_stage_n_3__exc__cmd_full_, exc_stage_n_3__exc__mispredict_, exc_stage_n_3__spec__dcache_miss_, exc_stage_n_3__spec__fencei_, exc_stage_n_3__spec__sfence_vma_, exc_stage_n_3__spec__dbreak_, exc_stage_n_3__spec__dret_, exc_stage_n_3__spec__mret_, exc_stage_n_3__spec__sret_, exc_stage_n_3__spec__wfi_, exc_stage_n_3__spec__csrw_, exc_stage_r_1__v_, exc_stage_r_1__queue_v_, exc_stage_n_2__ispec_v_, exc_stage_n_2__nspec_v_, exc_stage_n_2__exc__store_page_fault_, exc_stage_n_2__exc__load_page_fault_, exc_stage_n_2__exc__instr_page_fault_, exc_stage_n_2__exc__ecall_m_, exc_stage_n_2__exc__ecall_s_, exc_stage_n_2__exc__ecall_u_, exc_stage_n_2__exc__store_access_fault_, exc_stage_n_2__exc__store_misaligned_, exc_stage_n_2__exc__load_access_fault_, exc_stage_n_2__exc__load_misaligned_, exc_stage_n_2__exc__ebreak_, exc_stage_n_2__exc__illegal_instr_, exc_stage_n_2__exc__instr_access_fault_, exc_stage_r_1__exc__instr_misaligned_, exc_stage_n_2__exc__resume_, exc_stage_n_2__exc__itlb_miss_, exc_stage_n_2__exc__icache_miss_, exc_stage_r_1__exc__dcache_replay_, exc_stage_n_2__exc__dtlb_load_miss_, exc_stage_n_2__exc__dtlb_store_miss_, exc_stage_n_2__exc__itlb_fill_, exc_stage_n_2__exc__dtlb_fill_, exc_stage_n_2__exc___interrupt_, exc_stage_r_1__exc__cmd_full_, exc_stage_r_1__exc__mispredict_, exc_stage_r_1__spec__dcache_miss_, exc_stage_n_2__spec__fencei_, exc_stage_n_2__spec__sfence_vma_, exc_stage_n_2__spec__dbreak_, exc_stage_n_2__spec__dret_, exc_stage_n_2__spec__mret_, exc_stage_n_2__spec__sret_, exc_stage_n_2__spec__wfi_, exc_stage_n_2__spec__csrw_, exc_stage_r_0__v_, exc_stage_r_0__queue_v_, exc_stage_n_1__ispec_v_, exc_stage_n_1__nspec_v_, exc_stage_r_0__exc__store_page_fault_, exc_stage_r_0__exc__load_page_fault_, exc_stage_n_1__exc__instr_page_fault_, exc_stage_n_1__exc__ecall_m_, exc_stage_n_1__exc__ecall_s_, exc_stage_n_1__exc__ecall_u_, exc_stage_r_0__exc__store_access_fault_, exc_stage_r_0__exc__store_misaligned_, exc_stage_r_0__exc__load_access_fault_, exc_stage_r_0__exc__load_misaligned_, exc_stage_n_1__exc__ebreak_, exc_stage_r_0__exc__illegal_instr_, exc_stage_n_1__exc__instr_access_fault_, exc_stage_r_0__exc__instr_misaligned_, exc_stage_n_1__exc__resume_, exc_stage_n_1__exc__itlb_miss_, exc_stage_n_1__exc__icache_miss_, exc_stage_n_1__exc__dcache_replay_, exc_stage_r_0__exc__dtlb_load_miss_, exc_stage_r_0__exc__dtlb_store_miss_, exc_stage_n_1__exc__itlb_fill_, exc_stage_n_1__exc__dtlb_fill_, exc_stage_n_1__exc___interrupt_, exc_stage_n_1__exc__cmd_full_, exc_stage_n_1__exc__mispredict_, exc_stage_n_1__spec__dcache_miss_, exc_stage_n_1__spec__fencei_, exc_stage_n_1__spec__sfence_vma_, exc_stage_n_1__spec__dbreak_, exc_stage_n_1__spec__dret_, exc_stage_n_1__spec__mret_, exc_stage_n_1__spec__sret_, exc_stage_n_1__spec__wfi_, exc_stage_n_1__spec__csrw_ })
  );

  assign { \catchup.catchup_reservation_n_isrc1__64_ , \catchup.catchup_reservation_n_isrc1__63_ , \catchup.catchup_reservation_n_isrc1__62_ , \catchup.catchup_reservation_n_isrc1__61_ , \catchup.catchup_reservation_n_isrc1__60_ , \catchup.catchup_reservation_n_isrc1__59_ , \catchup.catchup_reservation_n_isrc1__58_ , \catchup.catchup_reservation_n_isrc1__57_ , \catchup.catchup_reservation_n_isrc1__56_ , \catchup.catchup_reservation_n_isrc1__55_ , \catchup.catchup_reservation_n_isrc1__54_ , \catchup.catchup_reservation_n_isrc1__53_ , \catchup.catchup_reservation_n_isrc1__52_ , \catchup.catchup_reservation_n_isrc1__51_ , \catchup.catchup_reservation_n_isrc1__50_ , \catchup.catchup_reservation_n_isrc1__49_ , \catchup.catchup_reservation_n_isrc1__48_ , \catchup.catchup_reservation_n_isrc1__47_ , \catchup.catchup_reservation_n_isrc1__46_ , \catchup.catchup_reservation_n_isrc1__45_ , \catchup.catchup_reservation_n_isrc1__44_ , \catchup.catchup_reservation_n_isrc1__43_ , \catchup.catchup_reservation_n_isrc1__42_ , \catchup.catchup_reservation_n_isrc1__41_ , \catchup.catchup_reservation_n_isrc1__40_ , \catchup.catchup_reservation_n_isrc1__39_ , \catchup.catchup_reservation_n_isrc1__38_ , \catchup.catchup_reservation_n_isrc1__37_ , \catchup.catchup_reservation_n_isrc1__36_ , \catchup.catchup_reservation_n_isrc1__35_ , \catchup.catchup_reservation_n_isrc1__34_ , \catchup.catchup_reservation_n_isrc1__33_ , \catchup.catchup_reservation_n_isrc1__32_ , \catchup.catchup_reservation_n_isrc1__31_ , \catchup.catchup_reservation_n_isrc1__30_ , \catchup.catchup_reservation_n_isrc1__29_ , \catchup.catchup_reservation_n_isrc1__28_ , \catchup.catchup_reservation_n_isrc1__27_ , \catchup.catchup_reservation_n_isrc1__26_ , \catchup.catchup_reservation_n_isrc1__25_ , \catchup.catchup_reservation_n_isrc1__24_ , \catchup.catchup_reservation_n_isrc1__23_ , \catchup.catchup_reservation_n_isrc1__22_ , \catchup.catchup_reservation_n_isrc1__21_ , \catchup.catchup_reservation_n_isrc1__20_ , \catchup.catchup_reservation_n_isrc1__19_ , \catchup.catchup_reservation_n_isrc1__18_ , \catchup.catchup_reservation_n_isrc1__17_ , \catchup.catchup_reservation_n_isrc1__16_ , \catchup.catchup_reservation_n_isrc1__15_ , \catchup.catchup_reservation_n_isrc1__14_ , \catchup.catchup_reservation_n_isrc1__13_ , \catchup.catchup_reservation_n_isrc1__12_ , \catchup.catchup_reservation_n_isrc1__11_ , \catchup.catchup_reservation_n_isrc1__10_ , \catchup.catchup_reservation_n_isrc1__9_ , \catchup.catchup_reservation_n_isrc1__8_ , \catchup.catchup_reservation_n_isrc1__7_ , \catchup.catchup_reservation_n_isrc1__6_ , \catchup.catchup_reservation_n_isrc1__5_ , \catchup.catchup_reservation_n_isrc1__4_ , \catchup.catchup_reservation_n_isrc1__3_ , \catchup.catchup_reservation_n_isrc1__2_ , \catchup.catchup_reservation_n_isrc1__1_ , \catchup.catchup_reservation_n_isrc1__0_  } = (N0)? \catchup.catchup_bypass_src1  : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                (N46)? reservation_r[389:325] : 1'b0;
  assign N0 = N45;
  assign { \catchup.catchup_reservation_n_isrc2__64_ , \catchup.catchup_reservation_n_isrc2__63_ , \catchup.catchup_reservation_n_isrc2__62_ , \catchup.catchup_reservation_n_isrc2__61_ , \catchup.catchup_reservation_n_isrc2__60_ , \catchup.catchup_reservation_n_isrc2__59_ , \catchup.catchup_reservation_n_isrc2__58_ , \catchup.catchup_reservation_n_isrc2__57_ , \catchup.catchup_reservation_n_isrc2__56_ , \catchup.catchup_reservation_n_isrc2__55_ , \catchup.catchup_reservation_n_isrc2__54_ , \catchup.catchup_reservation_n_isrc2__53_ , \catchup.catchup_reservation_n_isrc2__52_ , \catchup.catchup_reservation_n_isrc2__51_ , \catchup.catchup_reservation_n_isrc2__50_ , \catchup.catchup_reservation_n_isrc2__49_ , \catchup.catchup_reservation_n_isrc2__48_ , \catchup.catchup_reservation_n_isrc2__47_ , \catchup.catchup_reservation_n_isrc2__46_ , \catchup.catchup_reservation_n_isrc2__45_ , \catchup.catchup_reservation_n_isrc2__44_ , \catchup.catchup_reservation_n_isrc2__43_ , \catchup.catchup_reservation_n_isrc2__42_ , \catchup.catchup_reservation_n_isrc2__41_ , \catchup.catchup_reservation_n_isrc2__40_ , \catchup.catchup_reservation_n_isrc2__39_ , \catchup.catchup_reservation_n_isrc2__38_ , \catchup.catchup_reservation_n_isrc2__37_ , \catchup.catchup_reservation_n_isrc2__36_ , \catchup.catchup_reservation_n_isrc2__35_ , \catchup.catchup_reservation_n_isrc2__34_ , \catchup.catchup_reservation_n_isrc2__33_ , \catchup.catchup_reservation_n_isrc2__32_ , \catchup.catchup_reservation_n_isrc2__31_ , \catchup.catchup_reservation_n_isrc2__30_ , \catchup.catchup_reservation_n_isrc2__29_ , \catchup.catchup_reservation_n_isrc2__28_ , \catchup.catchup_reservation_n_isrc2__27_ , \catchup.catchup_reservation_n_isrc2__26_ , \catchup.catchup_reservation_n_isrc2__25_ , \catchup.catchup_reservation_n_isrc2__24_ , \catchup.catchup_reservation_n_isrc2__23_ , \catchup.catchup_reservation_n_isrc2__22_ , \catchup.catchup_reservation_n_isrc2__21_ , \catchup.catchup_reservation_n_isrc2__20_ , \catchup.catchup_reservation_n_isrc2__19_ , \catchup.catchup_reservation_n_isrc2__18_ , \catchup.catchup_reservation_n_isrc2__17_ , \catchup.catchup_reservation_n_isrc2__16_ , \catchup.catchup_reservation_n_isrc2__15_ , \catchup.catchup_reservation_n_isrc2__14_ , \catchup.catchup_reservation_n_isrc2__13_ , \catchup.catchup_reservation_n_isrc2__12_ , \catchup.catchup_reservation_n_isrc2__11_ , \catchup.catchup_reservation_n_isrc2__10_ , \catchup.catchup_reservation_n_isrc2__9_ , \catchup.catchup_reservation_n_isrc2__8_ , \catchup.catchup_reservation_n_isrc2__7_ , \catchup.catchup_reservation_n_isrc2__6_ , \catchup.catchup_reservation_n_isrc2__5_ , \catchup.catchup_reservation_n_isrc2__4_ , \catchup.catchup_reservation_n_isrc2__3_ , \catchup.catchup_reservation_n_isrc2__2_ , \catchup.catchup_reservation_n_isrc2__1_ , \catchup.catchup_reservation_n_isrc2__0_  } = (N1)? \catchup.catchup_bypass_src2  : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                (N49)? reservation_r[324:260] : 1'b0;
  assign N1 = N48;
  assign rs2_val_r = (N2)? \catchup.catchup_reservation_r [323:260] : 
                     (N52)? \catchup.catchup_reservation_r [128:65] : 1'b0;
  assign N2 = N51;
  assign { comp_stage_n_0__rd_data__65_, comp_stage_n_0__rd_data__64_, comp_stage_n_0__rd_data__63_, comp_stage_n_0__rd_data__62_, comp_stage_n_0__rd_data__61_, comp_stage_n_0__rd_data__60_, comp_stage_n_0__rd_data__59_, comp_stage_n_0__rd_data__58_, comp_stage_n_0__rd_data__57_, comp_stage_n_0__rd_data__56_, comp_stage_n_0__rd_data__55_, comp_stage_n_0__rd_data__54_, comp_stage_n_0__rd_data__53_, comp_stage_n_0__rd_data__52_, comp_stage_n_0__rd_data__51_, comp_stage_n_0__rd_data__50_, comp_stage_n_0__rd_data__49_, comp_stage_n_0__rd_data__48_, comp_stage_n_0__rd_data__47_, comp_stage_n_0__rd_data__46_, comp_stage_n_0__rd_data__45_, comp_stage_n_0__rd_data__44_, comp_stage_n_0__rd_data__43_, comp_stage_n_0__rd_data__42_, comp_stage_n_0__rd_data__41_, comp_stage_n_0__rd_data__40_, comp_stage_n_0__rd_data__39_, comp_stage_n_0__rd_data__38_, comp_stage_n_0__rd_data__37_, comp_stage_n_0__rd_data__36_, comp_stage_n_0__rd_data__35_, comp_stage_n_0__rd_data__34_, comp_stage_n_0__rd_data__33_, comp_stage_n_0__rd_data__32_, comp_stage_n_0__rd_data__31_, comp_stage_n_0__rd_data__30_, comp_stage_n_0__rd_data__29_, comp_stage_n_0__rd_data__28_, comp_stage_n_0__rd_data__27_, comp_stage_n_0__rd_data__26_, comp_stage_n_0__rd_data__25_, comp_stage_n_0__rd_data__24_, comp_stage_n_0__rd_data__23_, comp_stage_n_0__rd_data__22_, comp_stage_n_0__rd_data__21_, comp_stage_n_0__rd_data__20_, comp_stage_n_0__rd_data__19_, comp_stage_n_0__rd_data__18_, comp_stage_n_0__rd_data__17_, comp_stage_n_0__rd_data__16_, comp_stage_n_0__rd_data__15_, comp_stage_n_0__rd_data__14_, comp_stage_n_0__rd_data__13_, comp_stage_n_0__rd_data__12_, comp_stage_n_0__rd_data__11_, comp_stage_n_0__rd_data__10_, comp_stage_n_0__rd_data__9_, comp_stage_n_0__rd_data__8_, comp_stage_n_0__rd_data__7_, comp_stage_n_0__rd_data__6_, comp_stage_n_0__rd_data__5_, comp_stage_n_0__rd_data__4_, comp_stage_n_0__rd_data__3_, comp_stage_n_0__rd_data__2_, comp_stage_n_0__rd_data__1_, comp_stage_n_0__rd_data__0_ } = (N3)? dispatch_pkt_i[165:100] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N3 = injection;
  assign N4 = N53;
  assign { N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55 } = (N5)? pipe_int_early_data_lo : 
                                                                                                                                                                                                                                                                                                                                                                             (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N5 = pipe_int_early_data_v_lo;
  assign N6 = N54;
  assign { N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188 } = (N7)? pipe_sys_data_lo : 
                                                                                                                                                                                                                                                                                                                                                                                                                          (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N7 = pipe_sys_data_v_lo;
  assign N8 = N187;
  assign { N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255 } = (N9)? pipe_mem_early_data_lo : 
                                                                                                                                                                                                                                                                                                                                                                                                                          (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N9 = pipe_mem_early_data_v_lo;
  assign N10 = N254;
  assign { N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388 } = (N11)? pipe_aux_data_lo : 
                                                                                                                                                                                                                                                                                                                                                                                                                          (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = pipe_aux_data_v_lo;
  assign N12 = N387;
  assign { N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521 } = (N13)? pipe_int_catchup_data_lo : 
                                                                                                                                                                                                                                                                                                                                                                                                                          (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = pipe_int_catchup_data_v_lo;
  assign N14 = N520;
  assign { N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588 } = (N15)? pipe_mem_final_data_lo : 
                                                                                                                                                                                                                                                                                                                                                                                                                          (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = pipe_mem_final_data_v_lo;
  assign N16 = N587;
  assign { N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721 } = (N17)? pipe_mul_data_lo : 
                                                                                                                                                                                                                                                                                                                                                                                                                          (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N17 = pipe_mul_data_v_lo;
  assign N18 = N720;
  assign { N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788 } = (N19)? pipe_fma_data_lo : 
                                                                                                                                                                                                                                                                                                                                                                                                                          (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N19 = pipe_fma_data_v_lo;
  assign N20 = N787;
  assign { N858, N857, N856, N855, N854 } = (N3)? dispatch_pkt_i[38:34] : 
                                            (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N863, N862, N861, N860, N859 } = (N11)? { pipe_aux_fflags_lo_nv_, pipe_aux_fflags_lo_dz_, pipe_aux_fflags_lo_of_, pipe_aux_fflags_lo_uf_, pipe_aux_fflags_lo_nx_ } : 
                                            (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N873, N872, N871, N870, N869 } = (N19)? { pipe_fma_fflags_lo_nv_, pipe_fma_fflags_lo_dz_, pipe_fma_fflags_lo_of_, pipe_fma_fflags_lo_uf_, pipe_fma_fflags_lo_nx_ } : 
                                            (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign match_rs[0] = N882 | N884;
  assign N882 = N881 & N21;
  assign N881 = dispatch_pkt_i[277] & comp_stage_r_0__ird_w_v_;
  assign N884 = N883 & N22;
  assign N883 = dispatch_pkt_i[275] & comp_stage_r_0__frd_w_v_;
  assign match_rs[5] = N886 | N888;
  assign N886 = N885 & N23;
  assign N885 = dispatch_pkt_i[276] & comp_stage_r_0__ird_w_v_;
  assign N888 = N887 & N24;
  assign N887 = dispatch_pkt_i[274] & comp_stage_r_0__frd_w_v_;
  assign match_rs[10] = N889 & N25;
  assign N889 = dispatch_pkt_i[273] & comp_stage_r_0__frd_w_v_;
  assign match_rs[1] = N891 | N893;
  assign N891 = N890 & N26;
  assign N890 = dispatch_pkt_i[277] & comp_stage_r_1__ird_w_v_;
  assign N893 = N892 & N27;
  assign N892 = dispatch_pkt_i[275] & comp_stage_r_1__frd_w_v_;
  assign match_rs[6] = N895 | N897;
  assign N895 = N894 & N28;
  assign N894 = dispatch_pkt_i[276] & comp_stage_r_1__ird_w_v_;
  assign N897 = N896 & N29;
  assign N896 = dispatch_pkt_i[274] & comp_stage_r_1__frd_w_v_;
  assign match_rs[11] = N898 & N30;
  assign N898 = dispatch_pkt_i[273] & comp_stage_r_1__frd_w_v_;
  assign match_rs[2] = N900 | N902;
  assign N900 = N899 & N31;
  assign N899 = dispatch_pkt_i[277] & comp_stage_r_2__ird_w_v_;
  assign N902 = N901 & N32;
  assign N901 = dispatch_pkt_i[275] & comp_stage_r_2__frd_w_v_;
  assign match_rs[7] = N904 | N906;
  assign N904 = N903 & N33;
  assign N903 = dispatch_pkt_i[276] & comp_stage_r_2__ird_w_v_;
  assign N906 = N905 & N34;
  assign N905 = dispatch_pkt_i[274] & comp_stage_r_2__frd_w_v_;
  assign match_rs[12] = N907 & N35;
  assign N907 = dispatch_pkt_i[273] & comp_stage_r_2__frd_w_v_;
  assign match_rs[3] = N909 | N911;
  assign N909 = N908 & N36;
  assign N908 = dispatch_pkt_i[277] & iwb_pkt_o[78];
  assign N911 = N910 & N37;
  assign N910 = dispatch_pkt_i[275] & iwb_pkt_o[77];
  assign match_rs[8] = N913 | N915;
  assign N913 = N912 & N38;
  assign N912 = dispatch_pkt_i[276] & iwb_pkt_o[78];
  assign N915 = N914 & N39;
  assign N914 = dispatch_pkt_i[274] & iwb_pkt_o[77];
  assign match_rs[13] = N916 & N40;
  assign N916 = dispatch_pkt_i[273] & iwb_pkt_o[77];
  assign match_rs[4] = N917 & N41;
  assign N917 = dispatch_pkt_i[275] & fwb_pkt_o[77];
  assign match_rs[9] = N918 & N42;
  assign N918 = dispatch_pkt_i[274] & fwb_pkt_o[77];
  assign match_rs[14] = N919 & N43;
  assign N919 = dispatch_pkt_i[273] & fwb_pkt_o[77];
  assign _12_net_ = ~exc_stage_n_1__ispec_v_;
  assign br_pkt_o[42] = exc_stage_r_0__v_ & exc_stage_r_0__queue_v_;
  assign br_pkt_o[41] = br_pkt_o[42] & pipe_int_early_branch_lo;
  assign br_pkt_o[40] = br_pkt_o[42] & pipe_int_early_btaken_lo;
  assign br_pkt_o[39] = br_pkt_o[42] & exc_stage_n_1__ispec_v_;
  assign N45 = N920 & N44;
  assign N920 = reservation_r[440] & comp_stage_r_1__ird_w_v_;
  assign N46 = ~N45;
  assign N48 = N921 & N47;
  assign N921 = reservation_r[439] & comp_stage_r_1__ird_w_v_;
  assign N49 = ~N48;
  assign pipe_int_catchup_mispredict_lo = exc_stage_n_2__ispec_v_ & N50;
  assign N51 = \catchup.catchup_reservation_r [439];
  assign N52 = ~N51;
  assign pipe_long_fdata_yumi_lo = late_wb_grants_lo[2] & late_wb_yumi_i;
  assign pipe_long_idata_yumi_lo = late_wb_grants_lo[1] & late_wb_yumi_i;
  assign late_wb_v_o = N922 | late_wb_grants_lo[0];
  assign N922 = late_wb_grants_lo[2] | late_wb_grants_lo[1];
  assign injection = dispatch_pkt_i[365] & N923;
  assign N923 = ~dispatch_pkt_i[364];
  assign N53 = ~injection;
  assign N54 = ~pipe_int_early_data_v_lo;
  assign N121 = comp_stage_r_0__rd_data__65_ | N120;
  assign N122 = comp_stage_r_0__rd_data__64_ | N119;
  assign N123 = comp_stage_r_0__rd_data__63_ | N118;
  assign N124 = comp_stage_r_0__rd_data__62_ | N117;
  assign N125 = comp_stage_r_0__rd_data__61_ | N116;
  assign N126 = comp_stage_r_0__rd_data__60_ | N115;
  assign N127 = comp_stage_r_0__rd_data__59_ | N114;
  assign N128 = comp_stage_r_0__rd_data__58_ | N113;
  assign N129 = comp_stage_r_0__rd_data__57_ | N112;
  assign N130 = comp_stage_r_0__rd_data__56_ | N111;
  assign N131 = comp_stage_r_0__rd_data__55_ | N110;
  assign N132 = comp_stage_r_0__rd_data__54_ | N109;
  assign N133 = comp_stage_r_0__rd_data__53_ | N108;
  assign N134 = comp_stage_r_0__rd_data__52_ | N107;
  assign N135 = comp_stage_r_0__rd_data__51_ | N106;
  assign N136 = comp_stage_r_0__rd_data__50_ | N105;
  assign N137 = comp_stage_r_0__rd_data__49_ | N104;
  assign N138 = comp_stage_r_0__rd_data__48_ | N103;
  assign N139 = comp_stage_r_0__rd_data__47_ | N102;
  assign N140 = comp_stage_r_0__rd_data__46_ | N101;
  assign N141 = comp_stage_r_0__rd_data__45_ | N100;
  assign N142 = comp_stage_r_0__rd_data__44_ | N99;
  assign N143 = comp_stage_r_0__rd_data__43_ | N98;
  assign N144 = comp_stage_r_0__rd_data__42_ | N97;
  assign N145 = comp_stage_r_0__rd_data__41_ | N96;
  assign N146 = comp_stage_r_0__rd_data__40_ | N95;
  assign N147 = comp_stage_r_0__rd_data__39_ | N94;
  assign N148 = comp_stage_r_0__rd_data__38_ | N93;
  assign N149 = comp_stage_r_0__rd_data__37_ | N92;
  assign N150 = comp_stage_r_0__rd_data__36_ | N91;
  assign N151 = comp_stage_r_0__rd_data__35_ | N90;
  assign N152 = comp_stage_r_0__rd_data__34_ | N89;
  assign N153 = comp_stage_r_0__rd_data__33_ | N88;
  assign N154 = comp_stage_r_0__rd_data__32_ | N87;
  assign N155 = comp_stage_r_0__rd_data__31_ | N86;
  assign N156 = comp_stage_r_0__rd_data__30_ | N85;
  assign N157 = comp_stage_r_0__rd_data__29_ | N84;
  assign N158 = comp_stage_r_0__rd_data__28_ | N83;
  assign N159 = comp_stage_r_0__rd_data__27_ | N82;
  assign N160 = comp_stage_r_0__rd_data__26_ | N81;
  assign N161 = comp_stage_r_0__rd_data__25_ | N80;
  assign N162 = comp_stage_r_0__rd_data__24_ | N79;
  assign N163 = comp_stage_r_0__rd_data__23_ | N78;
  assign N164 = comp_stage_r_0__rd_data__22_ | N77;
  assign N165 = comp_stage_r_0__rd_data__21_ | N76;
  assign N166 = comp_stage_r_0__rd_data__20_ | N75;
  assign N167 = comp_stage_r_0__rd_data__19_ | N74;
  assign N168 = comp_stage_r_0__rd_data__18_ | N73;
  assign N169 = comp_stage_r_0__rd_data__17_ | N72;
  assign N170 = comp_stage_r_0__rd_data__16_ | N71;
  assign N171 = comp_stage_r_0__rd_data__15_ | N70;
  assign N172 = comp_stage_r_0__rd_data__14_ | N69;
  assign N173 = comp_stage_r_0__rd_data__13_ | N68;
  assign N174 = comp_stage_r_0__rd_data__12_ | N67;
  assign N175 = comp_stage_r_0__rd_data__11_ | N66;
  assign N176 = comp_stage_r_0__rd_data__10_ | N65;
  assign N177 = comp_stage_r_0__rd_data__9_ | N64;
  assign N178 = comp_stage_r_0__rd_data__8_ | N63;
  assign N179 = comp_stage_r_0__rd_data__7_ | N62;
  assign N180 = comp_stage_r_0__rd_data__6_ | N61;
  assign N181 = comp_stage_r_0__rd_data__5_ | N60;
  assign N182 = comp_stage_r_0__rd_data__4_ | N59;
  assign N183 = comp_stage_r_0__rd_data__3_ | N58;
  assign N184 = comp_stage_r_0__rd_data__2_ | N57;
  assign N185 = comp_stage_r_0__rd_data__1_ | N56;
  assign N186 = comp_stage_r_0__rd_data__0_ | N55;
  assign N187 = ~pipe_sys_data_v_lo;
  assign forward_data_0__65_ = N121 | N253;
  assign forward_data_0__64_ = N122 | N252;
  assign forward_data_0__63_ = N123 | N251;
  assign forward_data_0__62_ = N124 | N250;
  assign forward_data_0__61_ = N125 | N249;
  assign forward_data_0__60_ = N126 | N248;
  assign forward_data_0__59_ = N127 | N247;
  assign forward_data_0__58_ = N128 | N246;
  assign forward_data_0__57_ = N129 | N245;
  assign forward_data_0__56_ = N130 | N244;
  assign forward_data_0__55_ = N131 | N243;
  assign forward_data_0__54_ = N132 | N242;
  assign forward_data_0__53_ = N133 | N241;
  assign forward_data_0__52_ = N134 | N240;
  assign forward_data_0__51_ = N135 | N239;
  assign forward_data_0__50_ = N136 | N238;
  assign forward_data_0__49_ = N137 | N237;
  assign forward_data_0__48_ = N138 | N236;
  assign forward_data_0__47_ = N139 | N235;
  assign forward_data_0__46_ = N140 | N234;
  assign forward_data_0__45_ = N141 | N233;
  assign forward_data_0__44_ = N142 | N232;
  assign forward_data_0__43_ = N143 | N231;
  assign forward_data_0__42_ = N144 | N230;
  assign forward_data_0__41_ = N145 | N229;
  assign forward_data_0__40_ = N146 | N228;
  assign forward_data_0__39_ = N147 | N227;
  assign forward_data_0__38_ = N148 | N226;
  assign forward_data_0__37_ = N149 | N225;
  assign forward_data_0__36_ = N150 | N224;
  assign forward_data_0__35_ = N151 | N223;
  assign forward_data_0__34_ = N152 | N222;
  assign forward_data_0__33_ = N153 | N221;
  assign forward_data_0__32_ = N154 | N220;
  assign forward_data_0__31_ = N155 | N219;
  assign forward_data_0__30_ = N156 | N218;
  assign forward_data_0__29_ = N157 | N217;
  assign forward_data_0__28_ = N158 | N216;
  assign forward_data_0__27_ = N159 | N215;
  assign forward_data_0__26_ = N160 | N214;
  assign forward_data_0__25_ = N161 | N213;
  assign forward_data_0__24_ = N162 | N212;
  assign forward_data_0__23_ = N163 | N211;
  assign forward_data_0__22_ = N164 | N210;
  assign forward_data_0__21_ = N165 | N209;
  assign forward_data_0__20_ = N166 | N208;
  assign forward_data_0__19_ = N167 | N207;
  assign forward_data_0__18_ = N168 | N206;
  assign forward_data_0__17_ = N169 | N205;
  assign forward_data_0__16_ = N170 | N204;
  assign forward_data_0__15_ = N171 | N203;
  assign forward_data_0__14_ = N172 | N202;
  assign forward_data_0__13_ = N173 | N201;
  assign forward_data_0__12_ = N174 | N200;
  assign forward_data_0__11_ = N175 | N199;
  assign forward_data_0__10_ = N176 | N198;
  assign forward_data_0__9_ = N177 | N197;
  assign forward_data_0__8_ = N178 | N196;
  assign forward_data_0__7_ = N179 | N195;
  assign forward_data_0__6_ = N180 | N194;
  assign forward_data_0__5_ = N181 | N193;
  assign forward_data_0__4_ = N182 | N192;
  assign forward_data_0__3_ = N183 | N191;
  assign forward_data_0__2_ = N184 | N190;
  assign forward_data_0__1_ = N185 | N189;
  assign forward_data_0__0_ = N186 | N188;
  assign N254 = ~pipe_mem_early_data_v_lo;
  assign N321 = comp_stage_r_1__rd_data__65_ | N320;
  assign N322 = comp_stage_r_1__rd_data__64_ | N319;
  assign N323 = comp_stage_r_1__rd_data__63_ | N318;
  assign N324 = comp_stage_r_1__rd_data__62_ | N317;
  assign N325 = comp_stage_r_1__rd_data__61_ | N316;
  assign N326 = comp_stage_r_1__rd_data__60_ | N315;
  assign N327 = comp_stage_r_1__rd_data__59_ | N314;
  assign N328 = comp_stage_r_1__rd_data__58_ | N313;
  assign N329 = comp_stage_r_1__rd_data__57_ | N312;
  assign N330 = comp_stage_r_1__rd_data__56_ | N311;
  assign N331 = comp_stage_r_1__rd_data__55_ | N310;
  assign N332 = comp_stage_r_1__rd_data__54_ | N309;
  assign N333 = comp_stage_r_1__rd_data__53_ | N308;
  assign N334 = comp_stage_r_1__rd_data__52_ | N307;
  assign N335 = comp_stage_r_1__rd_data__51_ | N306;
  assign N336 = comp_stage_r_1__rd_data__50_ | N305;
  assign N337 = comp_stage_r_1__rd_data__49_ | N304;
  assign N338 = comp_stage_r_1__rd_data__48_ | N303;
  assign N339 = comp_stage_r_1__rd_data__47_ | N302;
  assign N340 = comp_stage_r_1__rd_data__46_ | N301;
  assign N341 = comp_stage_r_1__rd_data__45_ | N300;
  assign N342 = comp_stage_r_1__rd_data__44_ | N299;
  assign N343 = comp_stage_r_1__rd_data__43_ | N298;
  assign N344 = comp_stage_r_1__rd_data__42_ | N297;
  assign N345 = comp_stage_r_1__rd_data__41_ | N296;
  assign N346 = comp_stage_r_1__rd_data__40_ | N295;
  assign N347 = comp_stage_r_1__rd_data__39_ | N294;
  assign N348 = comp_stage_r_1__rd_data__38_ | N293;
  assign N349 = comp_stage_r_1__rd_data__37_ | N292;
  assign N350 = comp_stage_r_1__rd_data__36_ | N291;
  assign N351 = comp_stage_r_1__rd_data__35_ | N290;
  assign N352 = comp_stage_r_1__rd_data__34_ | N289;
  assign N353 = comp_stage_r_1__rd_data__33_ | N288;
  assign N354 = comp_stage_r_1__rd_data__32_ | N287;
  assign N355 = comp_stage_r_1__rd_data__31_ | N286;
  assign N356 = comp_stage_r_1__rd_data__30_ | N285;
  assign N357 = comp_stage_r_1__rd_data__29_ | N284;
  assign N358 = comp_stage_r_1__rd_data__28_ | N283;
  assign N359 = comp_stage_r_1__rd_data__27_ | N282;
  assign N360 = comp_stage_r_1__rd_data__26_ | N281;
  assign N361 = comp_stage_r_1__rd_data__25_ | N280;
  assign N362 = comp_stage_r_1__rd_data__24_ | N279;
  assign N363 = comp_stage_r_1__rd_data__23_ | N278;
  assign N364 = comp_stage_r_1__rd_data__22_ | N277;
  assign N365 = comp_stage_r_1__rd_data__21_ | N276;
  assign N366 = comp_stage_r_1__rd_data__20_ | N275;
  assign N367 = comp_stage_r_1__rd_data__19_ | N274;
  assign N368 = comp_stage_r_1__rd_data__18_ | N273;
  assign N369 = comp_stage_r_1__rd_data__17_ | N272;
  assign N370 = comp_stage_r_1__rd_data__16_ | N271;
  assign N371 = comp_stage_r_1__rd_data__15_ | N270;
  assign N372 = comp_stage_r_1__rd_data__14_ | N269;
  assign N373 = comp_stage_r_1__rd_data__13_ | N268;
  assign N374 = comp_stage_r_1__rd_data__12_ | N267;
  assign N375 = comp_stage_r_1__rd_data__11_ | N266;
  assign N376 = comp_stage_r_1__rd_data__10_ | N265;
  assign N377 = comp_stage_r_1__rd_data__9_ | N264;
  assign N378 = comp_stage_r_1__rd_data__8_ | N263;
  assign N379 = comp_stage_r_1__rd_data__7_ | N262;
  assign N380 = comp_stage_r_1__rd_data__6_ | N261;
  assign N381 = comp_stage_r_1__rd_data__5_ | N260;
  assign N382 = comp_stage_r_1__rd_data__4_ | N259;
  assign N383 = comp_stage_r_1__rd_data__3_ | N258;
  assign N384 = comp_stage_r_1__rd_data__2_ | N257;
  assign N385 = comp_stage_r_1__rd_data__1_ | N256;
  assign N386 = comp_stage_r_1__rd_data__0_ | N255;
  assign N387 = ~pipe_aux_data_v_lo;
  assign N454 = N321 | N453;
  assign N455 = N322 | N452;
  assign N456 = N323 | N451;
  assign N457 = N324 | N450;
  assign N458 = N325 | N449;
  assign N459 = N326 | N448;
  assign N460 = N327 | N447;
  assign N461 = N328 | N446;
  assign N462 = N329 | N445;
  assign N463 = N330 | N444;
  assign N464 = N331 | N443;
  assign N465 = N332 | N442;
  assign N466 = N333 | N441;
  assign N467 = N334 | N440;
  assign N468 = N335 | N439;
  assign N469 = N336 | N438;
  assign N470 = N337 | N437;
  assign N471 = N338 | N436;
  assign N472 = N339 | N435;
  assign N473 = N340 | N434;
  assign N474 = N341 | N433;
  assign N475 = N342 | N432;
  assign N476 = N343 | N431;
  assign N477 = N344 | N430;
  assign N478 = N345 | N429;
  assign N479 = N346 | N428;
  assign N480 = N347 | N427;
  assign N481 = N348 | N426;
  assign N482 = N349 | N425;
  assign N483 = N350 | N424;
  assign N484 = N351 | N423;
  assign N485 = N352 | N422;
  assign N486 = N353 | N421;
  assign N487 = N354 | N420;
  assign N488 = N355 | N419;
  assign N489 = N356 | N418;
  assign N490 = N357 | N417;
  assign N491 = N358 | N416;
  assign N492 = N359 | N415;
  assign N493 = N360 | N414;
  assign N494 = N361 | N413;
  assign N495 = N362 | N412;
  assign N496 = N363 | N411;
  assign N497 = N364 | N410;
  assign N498 = N365 | N409;
  assign N499 = N366 | N408;
  assign N500 = N367 | N407;
  assign N501 = N368 | N406;
  assign N502 = N369 | N405;
  assign N503 = N370 | N404;
  assign N504 = N371 | N403;
  assign N505 = N372 | N402;
  assign N506 = N373 | N401;
  assign N507 = N374 | N400;
  assign N508 = N375 | N399;
  assign N509 = N376 | N398;
  assign N510 = N377 | N397;
  assign N511 = N378 | N396;
  assign N512 = N379 | N395;
  assign N513 = N380 | N394;
  assign N514 = N381 | N393;
  assign N515 = N382 | N392;
  assign N516 = N383 | N391;
  assign N517 = N384 | N390;
  assign N518 = N385 | N389;
  assign N519 = N386 | N388;
  assign N520 = ~pipe_int_catchup_data_v_lo;
  assign forward_data_1__65_ = N454 | N586;
  assign forward_data_1__64_ = N455 | N585;
  assign forward_data_1__63_ = N456 | N584;
  assign forward_data_1__62_ = N457 | N583;
  assign forward_data_1__61_ = N458 | N582;
  assign forward_data_1__60_ = N459 | N581;
  assign forward_data_1__59_ = N460 | N580;
  assign forward_data_1__58_ = N461 | N579;
  assign forward_data_1__57_ = N462 | N578;
  assign forward_data_1__56_ = N463 | N577;
  assign forward_data_1__55_ = N464 | N576;
  assign forward_data_1__54_ = N465 | N575;
  assign forward_data_1__53_ = N466 | N574;
  assign forward_data_1__52_ = N467 | N573;
  assign forward_data_1__51_ = N468 | N572;
  assign forward_data_1__50_ = N469 | N571;
  assign forward_data_1__49_ = N470 | N570;
  assign forward_data_1__48_ = N471 | N569;
  assign forward_data_1__47_ = N472 | N568;
  assign forward_data_1__46_ = N473 | N567;
  assign forward_data_1__45_ = N474 | N566;
  assign forward_data_1__44_ = N475 | N565;
  assign forward_data_1__43_ = N476 | N564;
  assign forward_data_1__42_ = N477 | N563;
  assign forward_data_1__41_ = N478 | N562;
  assign forward_data_1__40_ = N479 | N561;
  assign forward_data_1__39_ = N480 | N560;
  assign forward_data_1__38_ = N481 | N559;
  assign forward_data_1__37_ = N482 | N558;
  assign forward_data_1__36_ = N483 | N557;
  assign forward_data_1__35_ = N484 | N556;
  assign forward_data_1__34_ = N485 | N555;
  assign forward_data_1__33_ = N486 | N554;
  assign forward_data_1__32_ = N487 | N553;
  assign forward_data_1__31_ = N488 | N552;
  assign forward_data_1__30_ = N489 | N551;
  assign forward_data_1__29_ = N490 | N550;
  assign forward_data_1__28_ = N491 | N549;
  assign forward_data_1__27_ = N492 | N548;
  assign forward_data_1__26_ = N493 | N547;
  assign forward_data_1__25_ = N494 | N546;
  assign forward_data_1__24_ = N495 | N545;
  assign forward_data_1__23_ = N496 | N544;
  assign forward_data_1__22_ = N497 | N543;
  assign forward_data_1__21_ = N498 | N542;
  assign forward_data_1__20_ = N499 | N541;
  assign forward_data_1__19_ = N500 | N540;
  assign forward_data_1__18_ = N501 | N539;
  assign forward_data_1__17_ = N502 | N538;
  assign forward_data_1__16_ = N503 | N537;
  assign forward_data_1__15_ = N504 | N536;
  assign forward_data_1__14_ = N505 | N535;
  assign forward_data_1__13_ = N506 | N534;
  assign forward_data_1__12_ = N507 | N533;
  assign forward_data_1__11_ = N508 | N532;
  assign forward_data_1__10_ = N509 | N531;
  assign forward_data_1__9_ = N510 | N530;
  assign forward_data_1__8_ = N511 | N529;
  assign forward_data_1__7_ = N512 | N528;
  assign forward_data_1__6_ = N513 | N527;
  assign forward_data_1__5_ = N514 | N526;
  assign forward_data_1__4_ = N515 | N525;
  assign forward_data_1__3_ = N516 | N524;
  assign forward_data_1__2_ = N517 | N523;
  assign forward_data_1__1_ = N518 | N522;
  assign forward_data_1__0_ = N519 | N521;
  assign N587 = ~pipe_mem_final_data_v_lo;
  assign N654 = comp_stage_r_2__rd_data__65_ | N653;
  assign N655 = comp_stage_r_2__rd_data__64_ | N652;
  assign N656 = comp_stage_r_2__rd_data__63_ | N651;
  assign N657 = comp_stage_r_2__rd_data__62_ | N650;
  assign N658 = comp_stage_r_2__rd_data__61_ | N649;
  assign N659 = comp_stage_r_2__rd_data__60_ | N648;
  assign N660 = comp_stage_r_2__rd_data__59_ | N647;
  assign N661 = comp_stage_r_2__rd_data__58_ | N646;
  assign N662 = comp_stage_r_2__rd_data__57_ | N645;
  assign N663 = comp_stage_r_2__rd_data__56_ | N644;
  assign N664 = comp_stage_r_2__rd_data__55_ | N643;
  assign N665 = comp_stage_r_2__rd_data__54_ | N642;
  assign N666 = comp_stage_r_2__rd_data__53_ | N641;
  assign N667 = comp_stage_r_2__rd_data__52_ | N640;
  assign N668 = comp_stage_r_2__rd_data__51_ | N639;
  assign N669 = comp_stage_r_2__rd_data__50_ | N638;
  assign N670 = comp_stage_r_2__rd_data__49_ | N637;
  assign N671 = comp_stage_r_2__rd_data__48_ | N636;
  assign N672 = comp_stage_r_2__rd_data__47_ | N635;
  assign N673 = comp_stage_r_2__rd_data__46_ | N634;
  assign N674 = comp_stage_r_2__rd_data__45_ | N633;
  assign N675 = comp_stage_r_2__rd_data__44_ | N632;
  assign N676 = comp_stage_r_2__rd_data__43_ | N631;
  assign N677 = comp_stage_r_2__rd_data__42_ | N630;
  assign N678 = comp_stage_r_2__rd_data__41_ | N629;
  assign N679 = comp_stage_r_2__rd_data__40_ | N628;
  assign N680 = comp_stage_r_2__rd_data__39_ | N627;
  assign N681 = comp_stage_r_2__rd_data__38_ | N626;
  assign N682 = comp_stage_r_2__rd_data__37_ | N625;
  assign N683 = comp_stage_r_2__rd_data__36_ | N624;
  assign N684 = comp_stage_r_2__rd_data__35_ | N623;
  assign N685 = comp_stage_r_2__rd_data__34_ | N622;
  assign N686 = comp_stage_r_2__rd_data__33_ | N621;
  assign N687 = comp_stage_r_2__rd_data__32_ | N620;
  assign N688 = comp_stage_r_2__rd_data__31_ | N619;
  assign N689 = comp_stage_r_2__rd_data__30_ | N618;
  assign N690 = comp_stage_r_2__rd_data__29_ | N617;
  assign N691 = comp_stage_r_2__rd_data__28_ | N616;
  assign N692 = comp_stage_r_2__rd_data__27_ | N615;
  assign N693 = comp_stage_r_2__rd_data__26_ | N614;
  assign N694 = comp_stage_r_2__rd_data__25_ | N613;
  assign N695 = comp_stage_r_2__rd_data__24_ | N612;
  assign N696 = comp_stage_r_2__rd_data__23_ | N611;
  assign N697 = comp_stage_r_2__rd_data__22_ | N610;
  assign N698 = comp_stage_r_2__rd_data__21_ | N609;
  assign N699 = comp_stage_r_2__rd_data__20_ | N608;
  assign N700 = comp_stage_r_2__rd_data__19_ | N607;
  assign N701 = comp_stage_r_2__rd_data__18_ | N606;
  assign N702 = comp_stage_r_2__rd_data__17_ | N605;
  assign N703 = comp_stage_r_2__rd_data__16_ | N604;
  assign N704 = comp_stage_r_2__rd_data__15_ | N603;
  assign N705 = comp_stage_r_2__rd_data__14_ | N602;
  assign N706 = comp_stage_r_2__rd_data__13_ | N601;
  assign N707 = comp_stage_r_2__rd_data__12_ | N600;
  assign N708 = comp_stage_r_2__rd_data__11_ | N599;
  assign N709 = comp_stage_r_2__rd_data__10_ | N598;
  assign N710 = comp_stage_r_2__rd_data__9_ | N597;
  assign N711 = comp_stage_r_2__rd_data__8_ | N596;
  assign N712 = comp_stage_r_2__rd_data__7_ | N595;
  assign N713 = comp_stage_r_2__rd_data__6_ | N594;
  assign N714 = comp_stage_r_2__rd_data__5_ | N593;
  assign N715 = comp_stage_r_2__rd_data__4_ | N592;
  assign N716 = comp_stage_r_2__rd_data__3_ | N591;
  assign N717 = comp_stage_r_2__rd_data__2_ | N590;
  assign N718 = comp_stage_r_2__rd_data__1_ | N589;
  assign N719 = comp_stage_r_2__rd_data__0_ | N588;
  assign N720 = ~pipe_mul_data_v_lo;
  assign forward_data_2__65_ = N654 | N786;
  assign forward_data_2__64_ = N655 | N785;
  assign forward_data_2__63_ = N656 | N784;
  assign forward_data_2__62_ = N657 | N783;
  assign forward_data_2__61_ = N658 | N782;
  assign forward_data_2__60_ = N659 | N781;
  assign forward_data_2__59_ = N660 | N780;
  assign forward_data_2__58_ = N661 | N779;
  assign forward_data_2__57_ = N662 | N778;
  assign forward_data_2__56_ = N663 | N777;
  assign forward_data_2__55_ = N664 | N776;
  assign forward_data_2__54_ = N665 | N775;
  assign forward_data_2__53_ = N666 | N774;
  assign forward_data_2__52_ = N667 | N773;
  assign forward_data_2__51_ = N668 | N772;
  assign forward_data_2__50_ = N669 | N771;
  assign forward_data_2__49_ = N670 | N770;
  assign forward_data_2__48_ = N671 | N769;
  assign forward_data_2__47_ = N672 | N768;
  assign forward_data_2__46_ = N673 | N767;
  assign forward_data_2__45_ = N674 | N766;
  assign forward_data_2__44_ = N675 | N765;
  assign forward_data_2__43_ = N676 | N764;
  assign forward_data_2__42_ = N677 | N763;
  assign forward_data_2__41_ = N678 | N762;
  assign forward_data_2__40_ = N679 | N761;
  assign forward_data_2__39_ = N680 | N760;
  assign forward_data_2__38_ = N681 | N759;
  assign forward_data_2__37_ = N682 | N758;
  assign forward_data_2__36_ = N683 | N757;
  assign forward_data_2__35_ = N684 | N756;
  assign forward_data_2__34_ = N685 | N755;
  assign forward_data_2__33_ = N686 | N754;
  assign forward_data_2__32_ = N687 | N753;
  assign forward_data_2__31_ = N688 | N752;
  assign forward_data_2__30_ = N689 | N751;
  assign forward_data_2__29_ = N690 | N750;
  assign forward_data_2__28_ = N691 | N749;
  assign forward_data_2__27_ = N692 | N748;
  assign forward_data_2__26_ = N693 | N747;
  assign forward_data_2__25_ = N694 | N746;
  assign forward_data_2__24_ = N695 | N745;
  assign forward_data_2__23_ = N696 | N744;
  assign forward_data_2__22_ = N697 | N743;
  assign forward_data_2__21_ = N698 | N742;
  assign forward_data_2__20_ = N699 | N741;
  assign forward_data_2__19_ = N700 | N740;
  assign forward_data_2__18_ = N701 | N739;
  assign forward_data_2__17_ = N702 | N738;
  assign forward_data_2__16_ = N703 | N737;
  assign forward_data_2__15_ = N704 | N736;
  assign forward_data_2__14_ = N705 | N735;
  assign forward_data_2__13_ = N706 | N734;
  assign forward_data_2__12_ = N707 | N733;
  assign forward_data_2__11_ = N708 | N732;
  assign forward_data_2__10_ = N709 | N731;
  assign forward_data_2__9_ = N710 | N730;
  assign forward_data_2__8_ = N711 | N729;
  assign forward_data_2__7_ = N712 | N728;
  assign forward_data_2__6_ = N713 | N727;
  assign forward_data_2__5_ = N714 | N726;
  assign forward_data_2__4_ = N715 | N725;
  assign forward_data_2__3_ = N716 | N724;
  assign forward_data_2__2_ = N717 | N723;
  assign forward_data_2__1_ = N718 | N722;
  assign forward_data_2__0_ = N719 | N721;
  assign N787 = ~pipe_fma_data_v_lo;
  assign forward_data_3__65_ = iwb_pkt_o[70] | N853;
  assign forward_data_3__64_ = iwb_pkt_o[69] | N852;
  assign forward_data_3__63_ = iwb_pkt_o[68] | N851;
  assign forward_data_3__62_ = iwb_pkt_o[67] | N850;
  assign forward_data_3__61_ = iwb_pkt_o[66] | N849;
  assign forward_data_3__60_ = iwb_pkt_o[65] | N848;
  assign forward_data_3__59_ = iwb_pkt_o[64] | N847;
  assign forward_data_3__58_ = iwb_pkt_o[63] | N846;
  assign forward_data_3__57_ = iwb_pkt_o[62] | N845;
  assign forward_data_3__56_ = iwb_pkt_o[61] | N844;
  assign forward_data_3__55_ = iwb_pkt_o[60] | N843;
  assign forward_data_3__54_ = iwb_pkt_o[59] | N842;
  assign forward_data_3__53_ = iwb_pkt_o[58] | N841;
  assign forward_data_3__52_ = iwb_pkt_o[57] | N840;
  assign forward_data_3__51_ = iwb_pkt_o[56] | N839;
  assign forward_data_3__50_ = iwb_pkt_o[55] | N838;
  assign forward_data_3__49_ = iwb_pkt_o[54] | N837;
  assign forward_data_3__48_ = iwb_pkt_o[53] | N836;
  assign forward_data_3__47_ = iwb_pkt_o[52] | N835;
  assign forward_data_3__46_ = iwb_pkt_o[51] | N834;
  assign forward_data_3__45_ = iwb_pkt_o[50] | N833;
  assign forward_data_3__44_ = iwb_pkt_o[49] | N832;
  assign forward_data_3__43_ = iwb_pkt_o[48] | N831;
  assign forward_data_3__42_ = iwb_pkt_o[47] | N830;
  assign forward_data_3__41_ = iwb_pkt_o[46] | N829;
  assign forward_data_3__40_ = iwb_pkt_o[45] | N828;
  assign forward_data_3__39_ = iwb_pkt_o[44] | N827;
  assign forward_data_3__38_ = iwb_pkt_o[43] | N826;
  assign forward_data_3__37_ = iwb_pkt_o[42] | N825;
  assign forward_data_3__36_ = iwb_pkt_o[41] | N824;
  assign forward_data_3__35_ = iwb_pkt_o[40] | N823;
  assign forward_data_3__34_ = iwb_pkt_o[39] | N822;
  assign forward_data_3__33_ = iwb_pkt_o[38] | N821;
  assign forward_data_3__32_ = iwb_pkt_o[37] | N820;
  assign forward_data_3__31_ = iwb_pkt_o[36] | N819;
  assign forward_data_3__30_ = iwb_pkt_o[35] | N818;
  assign forward_data_3__29_ = iwb_pkt_o[34] | N817;
  assign forward_data_3__28_ = iwb_pkt_o[33] | N816;
  assign forward_data_3__27_ = iwb_pkt_o[32] | N815;
  assign forward_data_3__26_ = iwb_pkt_o[31] | N814;
  assign forward_data_3__25_ = iwb_pkt_o[30] | N813;
  assign forward_data_3__24_ = iwb_pkt_o[29] | N812;
  assign forward_data_3__23_ = iwb_pkt_o[28] | N811;
  assign forward_data_3__22_ = iwb_pkt_o[27] | N810;
  assign forward_data_3__21_ = iwb_pkt_o[26] | N809;
  assign forward_data_3__20_ = iwb_pkt_o[25] | N808;
  assign forward_data_3__19_ = iwb_pkt_o[24] | N807;
  assign forward_data_3__18_ = iwb_pkt_o[23] | N806;
  assign forward_data_3__17_ = iwb_pkt_o[22] | N805;
  assign forward_data_3__16_ = iwb_pkt_o[21] | N804;
  assign forward_data_3__15_ = iwb_pkt_o[20] | N803;
  assign forward_data_3__14_ = iwb_pkt_o[19] | N802;
  assign forward_data_3__13_ = iwb_pkt_o[18] | N801;
  assign forward_data_3__12_ = iwb_pkt_o[17] | N800;
  assign forward_data_3__11_ = iwb_pkt_o[16] | N799;
  assign forward_data_3__10_ = iwb_pkt_o[15] | N798;
  assign forward_data_3__9_ = iwb_pkt_o[14] | N797;
  assign forward_data_3__8_ = iwb_pkt_o[13] | N796;
  assign forward_data_3__7_ = iwb_pkt_o[12] | N795;
  assign forward_data_3__6_ = iwb_pkt_o[11] | N794;
  assign forward_data_3__5_ = iwb_pkt_o[10] | N793;
  assign forward_data_3__4_ = iwb_pkt_o[9] | N792;
  assign forward_data_3__3_ = iwb_pkt_o[8] | N791;
  assign forward_data_3__2_ = iwb_pkt_o[7] | N790;
  assign forward_data_3__1_ = iwb_pkt_o[6] | N789;
  assign forward_data_3__0_ = iwb_pkt_o[5] | N788;
  assign N864 = comp_stage_r_1__fflags__nv_ | N863;
  assign N865 = comp_stage_r_1__fflags__dz_ | N862;
  assign N866 = comp_stage_r_1__fflags__of_ | N861;
  assign N867 = comp_stage_r_1__fflags__uf_ | N860;
  assign N868 = comp_stage_r_1__fflags__nx_ | N859;
  assign N874 = iwb_pkt_o[4] | N873;
  assign N875 = iwb_pkt_o[3] | N872;
  assign N876 = iwb_pkt_o[2] | N871;
  assign N877 = iwb_pkt_o[1] | N870;
  assign N878 = iwb_pkt_o[0] | N869;
  assign comp_stage_n_0__ird_w_v_ = dispatch_pkt_i[272] & exc_stage_n_0__v_;
  assign comp_stage_n_1__ird_w_v_ = comp_stage_r_0__ird_w_v_ & exc_stage_n_1__v_;
  assign comp_stage_n_2__ird_w_v_ = comp_stage_r_1__ird_w_v_ & exc_stage_n_2__v_;
  assign N879 = comp_stage_r_2__ird_w_v_ & exc_stage_n_3__v_;
  assign comp_stage_n_4__ird_w_v_ = iwb_pkt_o[78] & exc_stage_n_4__v_;
  assign comp_stage_n_0__frd_w_v_ = dispatch_pkt_i[271] & exc_stage_n_0__v_;
  assign comp_stage_n_1__frd_w_v_ = comp_stage_r_0__frd_w_v_ & exc_stage_n_1__v_;
  assign comp_stage_n_2__frd_w_v_ = comp_stage_r_1__frd_w_v_ & exc_stage_n_2__v_;
  assign N880 = comp_stage_r_2__frd_w_v_ & exc_stage_n_3__v_;
  assign comp_stage_n_4__frd_w_v_ = iwb_pkt_o[77] & exc_stage_n_4__v_;
  assign comp_stage_n_0__fflags__nv_ = N858 & exc_stage_n_0__v_;
  assign comp_stage_n_0__fflags__dz_ = N857 & exc_stage_n_0__v_;
  assign comp_stage_n_0__fflags__of_ = N856 & exc_stage_n_0__v_;
  assign comp_stage_n_0__fflags__uf_ = N855 & exc_stage_n_0__v_;
  assign comp_stage_n_0__fflags__nx_ = N854 & exc_stage_n_0__v_;
  assign comp_stage_n_1__fflags__nv_ = comp_stage_r_0__fflags__nv_ & exc_stage_n_1__v_;
  assign comp_stage_n_1__fflags__dz_ = comp_stage_r_0__fflags__dz_ & exc_stage_n_1__v_;
  assign comp_stage_n_1__fflags__of_ = comp_stage_r_0__fflags__of_ & exc_stage_n_1__v_;
  assign comp_stage_n_1__fflags__uf_ = comp_stage_r_0__fflags__uf_ & exc_stage_n_1__v_;
  assign comp_stage_n_1__fflags__nx_ = comp_stage_r_0__fflags__nx_ & exc_stage_n_1__v_;
  assign comp_stage_n_2__fflags__nv_ = N864 & exc_stage_n_2__v_;
  assign comp_stage_n_2__fflags__dz_ = N865 & exc_stage_n_2__v_;
  assign comp_stage_n_2__fflags__of_ = N866 & exc_stage_n_2__v_;
  assign comp_stage_n_2__fflags__uf_ = N867 & exc_stage_n_2__v_;
  assign comp_stage_n_2__fflags__nx_ = N868 & exc_stage_n_2__v_;
  assign comp_stage_n_3__fflags__nv_ = comp_stage_r_2__fflags__nv_ & exc_stage_n_3__v_;
  assign comp_stage_n_3__fflags__dz_ = comp_stage_r_2__fflags__dz_ & exc_stage_n_3__v_;
  assign comp_stage_n_3__fflags__of_ = comp_stage_r_2__fflags__of_ & exc_stage_n_3__v_;
  assign comp_stage_n_3__fflags__uf_ = comp_stage_r_2__fflags__uf_ & exc_stage_n_3__v_;
  assign comp_stage_n_3__fflags__nx_ = comp_stage_r_2__fflags__nx_ & exc_stage_n_3__v_;
  assign comp_stage_n_4__fflags__nv_ = N874 & exc_stage_n_4__v_;
  assign comp_stage_n_4__fflags__dz_ = N875 & exc_stage_n_4__v_;
  assign comp_stage_n_4__fflags__of_ = N876 & exc_stage_n_4__v_;
  assign comp_stage_n_4__fflags__uf_ = N877 & exc_stage_n_4__v_;
  assign comp_stage_n_4__fflags__nx_ = N878 & exc_stage_n_4__v_;
  assign comp_stage_n_3__ird_w_v_ = N879 & N924;
  assign N924 = ~commit_pkt_o[1];
  assign comp_stage_n_3__frd_w_v_ = N880 & N925;
  assign N925 = ~commit_pkt_o[0];
  assign exc_stage_n_0__v_ = dispatch_pkt_i[365] & N927;
  assign N927 = N926 | dispatch_pkt_i[362];
  assign N926 = ~commit_pkt_o[213];
  assign exc_stage_n_1__v_ = exc_stage_r_0__v_ & N929;
  assign N929 = N928 | exc_stage_n_1__nspec_v_;
  assign N928 = ~commit_pkt_o[213];
  assign exc_stage_n_2__v_ = exc_stage_r_1__v_ & N931;
  assign N931 = N930 | exc_stage_n_2__nspec_v_;
  assign N930 = ~commit_pkt_o[213];
  assign exc_stage_n_3__v_ = exc_stage_r_2__v_ & N932;
  assign N932 = commit_pkt_o[211] | exc_stage_n_3__nspec_v_;
  assign exc_stage_n_0__queue_v_ = dispatch_pkt_i[364] & N933;
  assign N933 = ~commit_pkt_o[213];
  assign exc_stage_n_1__queue_v_ = exc_stage_r_0__queue_v_ & N934;
  assign N934 = ~commit_pkt_o[213];
  assign exc_stage_n_2__queue_v_ = exc_stage_r_1__queue_v_ & N935;
  assign N935 = ~commit_pkt_o[213];
  assign exc_stage_n_1__exc__illegal_instr_ = exc_stage_r_0__exc__illegal_instr_ | pipe_sys_illegal_instr_lo;
  assign exc_stage_n_1__exc__instr_misaligned_ = exc_stage_r_0__exc__instr_misaligned_ | pipe_int_early_instr_misaligned_lo;
  assign exc_stage_n_1__exc__dtlb_store_miss_ = exc_stage_r_0__exc__dtlb_store_miss_ | pipe_mem_dtlb_store_miss_lo;
  assign exc_stage_n_1__exc__dtlb_load_miss_ = exc_stage_r_0__exc__dtlb_load_miss_ | pipe_mem_dtlb_load_miss_lo;
  assign exc_stage_n_1__exc__load_misaligned_ = exc_stage_r_0__exc__load_misaligned_ | pipe_mem_load_misaligned_lo;
  assign exc_stage_n_1__exc__load_access_fault_ = exc_stage_r_0__exc__load_access_fault_ | pipe_mem_load_access_fault_lo;
  assign exc_stage_n_1__exc__load_page_fault_ = exc_stage_r_0__exc__load_page_fault_ | pipe_mem_load_page_fault_lo;
  assign exc_stage_n_1__exc__store_misaligned_ = exc_stage_r_0__exc__store_misaligned_ | pipe_mem_store_misaligned_lo;
  assign exc_stage_n_1__exc__store_access_fault_ = exc_stage_r_0__exc__store_access_fault_ | pipe_mem_store_access_fault_lo;
  assign exc_stage_n_1__exc__store_page_fault_ = exc_stage_r_0__exc__store_page_fault_ | pipe_mem_store_page_fault_lo;
  assign exc_stage_n_2__exc__instr_misaligned_ = exc_stage_r_1__exc__instr_misaligned_ | pipe_int_catchup_instr_misaligned_lo;
  assign exc_stage_n_2__exc__mispredict_ = exc_stage_r_1__exc__mispredict_ | pipe_int_catchup_mispredict_lo;
  assign exc_stage_n_2__exc__dcache_replay_ = exc_stage_r_1__exc__dcache_replay_ | pipe_mem_dcache_replay_lo;
  assign exc_stage_n_2__spec__dcache_miss_ = exc_stage_r_1__spec__dcache_miss_ | pipe_mem_dcache_miss_lo;
  assign exc_stage_n_2__exc__cmd_full_ = exc_stage_r_1__exc__cmd_full_ | N969;
  assign N969 = N968 & cmd_full_n_i;
  assign N968 = N967 | exc_stage_n_3__spec__csrw_;
  assign N967 = N966 | exc_stage_n_3__spec__wfi_;
  assign N966 = N965 | exc_stage_n_3__spec__sret_;
  assign N965 = N964 | exc_stage_n_3__spec__mret_;
  assign N964 = N963 | exc_stage_n_3__spec__dret_;
  assign N963 = N962 | exc_stage_n_3__spec__dbreak_;
  assign N962 = N961 | exc_stage_n_3__spec__sfence_vma_;
  assign N961 = N960 | exc_stage_n_3__spec__fencei_;
  assign N960 = N959 | exc_stage_n_3__spec__dcache_miss_;
  assign N959 = N958 | exc_stage_n_3__exc__mispredict_;
  assign N958 = N957 | exc_stage_n_3__exc__cmd_full_;
  assign N957 = N956 | exc_stage_n_3__exc___interrupt_;
  assign N956 = N955 | exc_stage_n_3__exc__dtlb_fill_;
  assign N955 = N954 | exc_stage_n_3__exc__itlb_fill_;
  assign N954 = N953 | exc_stage_n_3__exc__dtlb_store_miss_;
  assign N953 = N952 | exc_stage_n_3__exc__dtlb_load_miss_;
  assign N952 = N951 | exc_stage_n_3__exc__dcache_replay_;
  assign N951 = N950 | exc_stage_n_3__exc__icache_miss_;
  assign N950 = N949 | exc_stage_n_3__exc__itlb_miss_;
  assign N949 = N948 | exc_stage_n_3__exc__resume_;
  assign N948 = N947 | exc_stage_n_3__exc__instr_misaligned_;
  assign N947 = N946 | exc_stage_n_3__exc__instr_access_fault_;
  assign N946 = N945 | exc_stage_n_3__exc__illegal_instr_;
  assign N945 = N944 | exc_stage_n_3__exc__ebreak_;
  assign N944 = N943 | exc_stage_n_3__exc__load_misaligned_;
  assign N943 = N942 | exc_stage_n_3__exc__load_access_fault_;
  assign N942 = N941 | exc_stage_n_3__exc__store_misaligned_;
  assign N941 = N940 | exc_stage_n_3__exc__store_access_fault_;
  assign N940 = N939 | exc_stage_n_3__exc__ecall_u_;
  assign N939 = N938 | exc_stage_n_3__exc__ecall_s_;
  assign N938 = N937 | exc_stage_n_3__exc__ecall_m_;
  assign N937 = N936 | exc_stage_n_3__exc__instr_page_fault_;
  assign N936 = exc_stage_n_3__exc__store_page_fault_ | exc_stage_n_3__exc__load_page_fault_;

endmodule



module bp_be_top
(
  clk_i,
  reset_i,
  cfg_bus_i,
  fe_queue_i,
  fe_queue_v_i,
  fe_queue_ready_and_o,
  fe_cmd_o,
  fe_cmd_v_o,
  fe_cmd_yumi_i,
  cache_req_o,
  cache_req_v_o,
  cache_req_yumi_i,
  cache_req_lock_i,
  cache_req_metadata_o,
  cache_req_metadata_v_o,
  cache_req_id_i,
  cache_req_critical_i,
  cache_req_last_i,
  cache_req_credits_full_i,
  cache_req_credits_empty_i,
  tag_mem_pkt_v_i,
  tag_mem_pkt_i,
  tag_mem_o,
  tag_mem_pkt_yumi_o,
  data_mem_pkt_v_i,
  data_mem_pkt_i,
  data_mem_o,
  data_mem_pkt_yumi_o,
  stat_mem_pkt_v_i,
  stat_mem_pkt_i,
  stat_mem_o,
  stat_mem_pkt_yumi_o,
  debug_irq_i,
  timer_irq_i,
  software_irq_i,
  m_external_irq_i,
  s_external_irq_i
);

  input [60:0] cfg_bus_i;
  input [173:0] fe_queue_i;
  output [113:0] fe_cmd_o;
  output [116:0] cache_req_o;
  output [3:0] cache_req_metadata_o;
  input [0:0] cache_req_id_i;
  input [34:0] tag_mem_pkt_i;
  output [22:0] tag_mem_o;
  input [142:0] data_mem_pkt_i;
  output [511:0] data_mem_o;
  input [10:0] stat_mem_pkt_i;
  output [14:0] stat_mem_o;
  input clk_i;
  input reset_i;
  input fe_queue_v_i;
  input fe_cmd_yumi_i;
  input cache_req_yumi_i;
  input cache_req_lock_i;
  input cache_req_critical_i;
  input cache_req_last_i;
  input cache_req_credits_full_i;
  input cache_req_credits_empty_i;
  input tag_mem_pkt_v_i;
  input data_mem_pkt_v_i;
  input stat_mem_pkt_v_i;
  input debug_irq_i;
  input timer_irq_i;
  input software_irq_i;
  input m_external_irq_i;
  input s_external_irq_i;
  output fe_queue_ready_and_o;
  output fe_cmd_v_o;
  output cache_req_v_o;
  output cache_req_metadata_v_o;
  output tag_mem_pkt_yumi_o;
  output data_mem_pkt_yumi_o;
  output stat_mem_pkt_yumi_o;
  wire [113:0] fe_cmd_o;
  wire [116:0] cache_req_o;
  wire [3:0] cache_req_metadata_o;
  wire [22:0] tag_mem_o;
  wire [511:0] data_mem_o;
  wire [14:0] stat_mem_o;
  wire fe_queue_ready_and_o,fe_cmd_v_o,cache_req_v_o,cache_req_metadata_v_o,
  tag_mem_pkt_yumi_o,data_mem_pkt_yumi_o,stat_mem_pkt_yumi_o,resume_lo,poison_isd_lo,
  clear_iss_lo,suppress_iss_lo,irq_waiting_lo,mem_busy_lo,cmd_full_n_lo,cmd_full_r_lo,
  mem_ordered_lo,fdiv_busy_lo,idiv_busy_lo,ispec_v,hazard_v,ordered_v,late_wb_yumi_li,
  decode_info_lo_u_mode_,decode_info_lo_s_mode_,decode_info_lo_m_mode_,
  decode_info_lo_debug_mode_,decode_info_lo_tsr_,decode_info_lo_tw_,decode_info_lo_tvm_,
  decode_info_lo_ebreakm_,decode_info_lo_ebreaks_,decode_info_lo_ebreaku_,
  decode_info_lo_fpu_en_,decode_info_lo_cycle_en_,decode_info_lo_instret_en_,irq_pending_lo,
  late_wb_v_lo,late_wb_force_lo;
  wire [263:0] issue_pkt;
  wire [38:0] expected_npc_lo;
  wire [42:0] br_pkt;
  wire [213:0] commit_pkt;
  wire [365:0] dispatch_pkt;
  wire [78:0] late_wb_pkt,iwb_pkt,fwb_pkt;
  wire [32:0] trans_info_lo;

  bp_be_director_00
  director
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .cfg_bus_i(cfg_bus_i),
    .issue_pkt_i(issue_pkt),
    .expected_npc_o(expected_npc_lo),
    .poison_isd_o(poison_isd_lo),
    .clear_iss_o(clear_iss_lo),
    .suppress_iss_o(suppress_iss_lo),
    .resume_o(resume_lo),
    .irq_waiting_i(irq_waiting_lo),
    .mem_busy_i(mem_busy_lo),
    .cmd_full_n_o(cmd_full_n_lo),
    .cmd_full_r_o(cmd_full_r_lo),
    .fe_cmd_o(fe_cmd_o),
    .fe_cmd_v_o(fe_cmd_v_o),
    .fe_cmd_yumi_i(fe_cmd_yumi_i),
    .br_pkt_i(br_pkt),
    .commit_pkt_i(commit_pkt)
  );


  bp_be_detector_00
  detector
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .issue_pkt_i(issue_pkt),
    .cmd_full_i(cmd_full_r_lo),
    .credits_full_i(cache_req_credits_full_i),
    .credits_empty_i(cache_req_credits_empty_i),
    .idiv_busy_i(idiv_busy_lo),
    .fdiv_busy_i(fdiv_busy_lo),
    .mem_busy_i(mem_busy_lo),
    .mem_ordered_i(mem_ordered_lo),
    .hazard_v_o(hazard_v),
    .ordered_v_o(ordered_v),
    .dispatch_pkt_i(dispatch_pkt),
    .commit_pkt_i(commit_pkt),
    .late_wb_pkt_i(late_wb_pkt),
    .late_wb_yumi_i(late_wb_yumi_li),
    .ispec_v_o(ispec_v)
  );


  bp_be_scheduler_00
  scheduler
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .issue_pkt_o(issue_pkt),
    .expected_npc_i(expected_npc_lo),
    .clear_iss_i(clear_iss_lo),
    .suppress_iss_i(suppress_iss_lo),
    .resume_i(resume_lo),
    .decode_info_i({ decode_info_lo_u_mode_, decode_info_lo_s_mode_, decode_info_lo_m_mode_, decode_info_lo_debug_mode_, decode_info_lo_tsr_, decode_info_lo_tw_, decode_info_lo_tvm_, decode_info_lo_ebreakm_, decode_info_lo_ebreaks_, decode_info_lo_ebreaku_, decode_info_lo_fpu_en_, decode_info_lo_cycle_en_, decode_info_lo_instret_en_ }),
    .hazard_v_i(hazard_v),
    .irq_pending_i(irq_pending_lo),
    .ispec_v_i(ispec_v),
    .poison_isd_i(poison_isd_lo),
    .ordered_v_i(ordered_v),
    .trans_info_i(trans_info_lo),
    .fe_queue_i(fe_queue_i),
    .fe_queue_v_i(fe_queue_v_i),
    .fe_queue_ready_and_o(fe_queue_ready_and_o),
    .dispatch_pkt_o(dispatch_pkt),
    .commit_pkt_i(commit_pkt),
    .iwb_pkt_i(iwb_pkt),
    .fwb_pkt_i(fwb_pkt),
    .late_wb_pkt_i(late_wb_pkt),
    .late_wb_v_i(late_wb_v_lo),
    .late_wb_force_i(late_wb_force_lo),
    .late_wb_yumi_o(late_wb_yumi_li)
  );


  bp_be_calculator_top_00
  calculator
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .cfg_bus_i(cfg_bus_i),
    .dispatch_pkt_i(dispatch_pkt),
    .idiv_busy_o(idiv_busy_lo),
    .fdiv_busy_o(fdiv_busy_lo),
    .mem_busy_o(mem_busy_lo),
    .mem_ordered_o(mem_ordered_lo),
    .decode_info_o({ decode_info_lo_u_mode_, decode_info_lo_s_mode_, decode_info_lo_m_mode_, decode_info_lo_debug_mode_, decode_info_lo_tsr_, decode_info_lo_tw_, decode_info_lo_tvm_, decode_info_lo_ebreakm_, decode_info_lo_ebreaks_, decode_info_lo_ebreaku_, decode_info_lo_fpu_en_, decode_info_lo_cycle_en_, decode_info_lo_instret_en_ }),
    .trans_info_o(trans_info_lo),
    .cmd_full_n_i(cmd_full_n_lo),
    .commit_pkt_o(commit_pkt),
    .br_pkt_o(br_pkt),
    .iwb_pkt_o(iwb_pkt),
    .fwb_pkt_o(fwb_pkt),
    .late_wb_pkt_o(late_wb_pkt),
    .late_wb_v_o(late_wb_v_lo),
    .late_wb_force_o(late_wb_force_lo),
    .late_wb_yumi_i(late_wb_yumi_li),
    .debug_irq_i(debug_irq_i),
    .timer_irq_i(timer_irq_i),
    .software_irq_i(software_irq_i),
    .m_external_irq_i(m_external_irq_i),
    .s_external_irq_i(s_external_irq_i),
    .irq_waiting_o(irq_waiting_lo),
    .irq_pending_o(irq_pending_lo),
    .cache_req_o(cache_req_o),
    .cache_req_v_o(cache_req_v_o),
    .cache_req_yumi_i(cache_req_yumi_i),
    .cache_req_lock_i(cache_req_lock_i),
    .cache_req_metadata_o(cache_req_metadata_o),
    .cache_req_metadata_v_o(cache_req_metadata_v_o),
    .cache_req_id_i(cache_req_id_i[0]),
    .cache_req_critical_i(cache_req_critical_i),
    .cache_req_last_i(cache_req_last_i),
    .cache_req_credits_full_i(cache_req_credits_full_i),
    .cache_req_credits_empty_i(cache_req_credits_empty_i),
    .data_mem_pkt_v_i(data_mem_pkt_v_i),
    .data_mem_pkt_i(data_mem_pkt_i),
    .data_mem_pkt_yumi_o(data_mem_pkt_yumi_o),
    .data_mem_o(data_mem_o),
    .tag_mem_pkt_v_i(tag_mem_pkt_v_i),
    .tag_mem_pkt_i(tag_mem_pkt_i),
    .tag_mem_pkt_yumi_o(tag_mem_pkt_yumi_o),
    .tag_mem_o(tag_mem_o),
    .stat_mem_pkt_v_i(stat_mem_pkt_v_i),
    .stat_mem_pkt_i(stat_mem_pkt_i),
    .stat_mem_pkt_yumi_o(stat_mem_pkt_yumi_o),
    .stat_mem_o(stat_mem_o)
  );


endmodule

