

module bsg_circular_ptr_00000004_1
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [0:0] add_i;
  output [1:0] o;
  output [1:0] n_o;
  input clk;
  input reset_i;
  wire [1:0] o,n_o,\genblk1.genblk1.ptr_r_p1 ;
  wire N0,N1,N2;
  reg o_1_sv2v_reg,o_0_sv2v_reg;
  assign o[1] = o_1_sv2v_reg;
  assign o[0] = o_0_sv2v_reg;
  assign \genblk1.genblk1.ptr_r_p1  = o + 1'b1;
  assign n_o = (N0)? \genblk1.genblk1.ptr_r_p1  : 
               (N1)? o : 1'b0;
  assign N0 = add_i[0];
  assign N1 = N2;
  assign N2 = ~add_i[0];

  always @(posedge clk) begin
    if(reset_i) begin
      o_1_sv2v_reg <= 1'b0;
      o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      o_1_sv2v_reg <= n_o[1];
      o_0_sv2v_reg <= n_o[0];
    end 
  end


endmodule



module bsg_fifo_tracker_00000004
(
  clk_i,
  reset_i,
  enq_i,
  deq_i,
  wptr_r_o,
  rptr_r_o,
  rptr_n_o,
  full_o,
  empty_o
);

  output [1:0] wptr_r_o;
  output [1:0] rptr_r_o;
  output [1:0] rptr_n_o;
  input clk_i;
  input reset_i;
  input enq_i;
  input deq_i;
  output full_o;
  output empty_o;
  wire [1:0] wptr_r_o,rptr_r_o,rptr_n_o;
  wire full_o,empty_o,enq_r,deq_r,N0,equal_ptrs,sv2v_dc_1,sv2v_dc_2;
  reg deq_r_sv2v_reg,enq_r_sv2v_reg;
  assign deq_r = deq_r_sv2v_reg;
  assign enq_r = enq_r_sv2v_reg;

  bsg_circular_ptr_00000004_1
  rptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(deq_i),
    .o(rptr_r_o),
    .n_o(rptr_n_o)
  );


  bsg_circular_ptr_00000004_1
  wptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(enq_i),
    .o(wptr_r_o),
    .n_o({ sv2v_dc_1, sv2v_dc_2 })
  );

  assign equal_ptrs = rptr_r_o == wptr_r_o;
  assign N0 = enq_i | deq_i;
  assign empty_o = equal_ptrs & deq_r;
  assign full_o = equal_ptrs & enq_r;

  always @(posedge clk_i) begin
    if(reset_i) begin
      deq_r_sv2v_reg <= 1'b1;
      enq_r_sv2v_reg <= 1'b0;
    end else if(N0) begin
      deq_r_sv2v_reg <= deq_i;
      enq_r_sv2v_reg <= enq_i;
    end 
  end


endmodule



module bsg_fifo_1r1w_small_unhardened_000000c1_00000004_0
(
  clk_i,
  reset_i,
  v_i,
  ready_param_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [192:0] data_i;
  output [192:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_param_o;
  output v_o;
  wire [192:0] data_o;
  wire ready_param_o,v_o,enque,full,empty,sv2v_dc_1,sv2v_dc_2;
  wire [1:0] wptr_r,rptr_r;

  bsg_fifo_tracker_00000004
  ft
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .enq_i(enque),
    .deq_i(yumi_i),
    .wptr_r_o(wptr_r),
    .rptr_r_o(rptr_r),
    .rptr_n_o({ sv2v_dc_1, sv2v_dc_2 }),
    .full_o(full),
    .empty_o(empty)
  );


  bsg_mem_1r1w
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enque),
    .w_addr_i(wptr_r),
    .w_data_i(data_i),
    .r_v_i(v_o),
    .r_addr_i(rptr_r),
    .r_data_o(data_o)
  );

  assign enque = v_i & ready_param_o;
  assign ready_param_o = ~full;
  assign v_o = ~empty;

endmodule



module bsg_fifo_1r1w_small_000000c1_00000004
(
  clk_i,
  reset_i,
  v_i,
  ready_param_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [192:0] data_i;
  output [192:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_param_o;
  output v_o;
  wire [192:0] data_o;
  wire ready_param_o,v_o;

  bsg_fifo_1r1w_small_unhardened_000000c1_00000004_0
  \unhardened.un.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_param_o(ready_param_o),
    .data_i(data_i),
    .v_o(v_o),
    .data_o(data_o),
    .yumi_i(yumi_i)
  );


endmodule



module bsg_circular_ptr_slots_p3_max_add_p1
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [0:0] add_i;
  output [1:0] o;
  output [1:0] n_o;
  input clk;
  input reset_i;
  wire [1:0] o,n_o,ptr_nowrap;
  wire N0,N1,N2,N3,N4,N5;
  wire [2:0] ptr_wrap;
  reg o_1_sv2v_reg,o_0_sv2v_reg;
  assign o[1] = o_1_sv2v_reg;
  assign o[0] = o_0_sv2v_reg;
  assign ptr_nowrap = o + add_i[0];
  assign { N4, N3, N2 } = o - { 1'b1, 1'b1 };
  assign ptr_wrap = { N4, N3, N2 } + add_i[0];
  assign n_o = (N0)? ptr_wrap[1:0] : 
               (N1)? ptr_nowrap : 1'b0;
  assign N0 = N5;
  assign N1 = ptr_wrap[2];
  assign N5 = ~ptr_wrap[2];

  always @(posedge clk) begin
    if(reset_i) begin
      o_1_sv2v_reg <= 1'b0;
      o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      o_1_sv2v_reg <= n_o[1];
      o_0_sv2v_reg <= n_o[0];
    end 
  end


endmodule



module bsg_fifo_tracker_els_p3
(
  clk_i,
  reset_i,
  enq_i,
  deq_i,
  wptr_r_o,
  rptr_r_o,
  rptr_n_o,
  full_o,
  empty_o
);

  output [1:0] wptr_r_o;
  output [1:0] rptr_r_o;
  output [1:0] rptr_n_o;
  input clk_i;
  input reset_i;
  input enq_i;
  input deq_i;
  output full_o;
  output empty_o;
  wire [1:0] wptr_r_o,rptr_r_o,rptr_n_o;
  wire full_o,empty_o,enq_r,deq_r,N0,equal_ptrs,sv2v_dc_1,sv2v_dc_2;
  reg deq_r_sv2v_reg,enq_r_sv2v_reg;
  assign deq_r = deq_r_sv2v_reg;
  assign enq_r = enq_r_sv2v_reg;

  bsg_circular_ptr_slots_p3_max_add_p1
  rptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(deq_i),
    .o(rptr_r_o),
    .n_o(rptr_n_o)
  );


  bsg_circular_ptr_slots_p3_max_add_p1
  wptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(enq_i),
    .o(wptr_r_o),
    .n_o({ sv2v_dc_1, sv2v_dc_2 })
  );

  assign equal_ptrs = rptr_r_o == wptr_r_o;
  assign N0 = enq_i | deq_i;
  assign empty_o = equal_ptrs & deq_r;
  assign full_o = equal_ptrs & enq_r;

  always @(posedge clk_i) begin
    if(reset_i) begin
      deq_r_sv2v_reg <= 1'b1;
      enq_r_sv2v_reg <= 1'b0;
    end else if(N0) begin
      deq_r_sv2v_reg <= deq_i;
      enq_r_sv2v_reg <= enq_i;
    end 
  end


endmodule



module bsg_fifo_1r1w_small_unhardened_width_p1_els_p3_ready_THEN_valid_p1
(
  clk_i,
  reset_i,
  v_i,
  ready_param_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_param_o;
  output v_o;
  wire [0:0] data_o;
  wire ready_param_o,v_o,full,empty,sv2v_dc_1,sv2v_dc_2;
  wire [1:0] wptr_r,rptr_r;

  bsg_fifo_tracker_els_p3
  ft
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .enq_i(v_i),
    .deq_i(yumi_i),
    .wptr_r_o(wptr_r),
    .rptr_r_o(rptr_r),
    .rptr_n_o({ sv2v_dc_1, sv2v_dc_2 }),
    .full_o(full),
    .empty_o(empty)
  );


  bsg_mem_1r1w
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(v_i),
    .w_addr_i(wptr_r),
    .w_data_i(data_i[0]),
    .r_v_i(v_o),
    .r_addr_i(rptr_r),
    .r_data_o(data_o[0])
  );

  assign ready_param_o = ~full;
  assign v_o = ~empty;

endmodule



module bsg_fifo_1r1w_small_width_p1_els_p3_ready_THEN_valid_p1
(
  clk_i,
  reset_i,
  v_i,
  ready_param_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_param_o;
  output v_o;
  wire [0:0] data_o;
  wire ready_param_o,v_o;

  bsg_fifo_1r1w_small_unhardened_width_p1_els_p3_ready_THEN_valid_p1
  \unhardened.un.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_param_o(ready_param_o),
    .data_i(data_i[0]),
    .v_o(v_o),
    .data_o(data_o[0]),
    .yumi_i(yumi_i)
  );


endmodule



module bsg_two_fifo_000000c1
(
  clk_i,
  reset_i,
  ready_param_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [192:0] data_i;
  output [192:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_param_o;
  output v_o;
  wire [192:0] data_o;
  wire ready_param_o,v_o,enq_i,tail_r,_0_net_,head_r,empty_r,full_r,N0,N1,N2,N3,N4,N5,
  N6,N7,N8,N9,N10,N11,N12,N13,N14;
  reg full_r_sv2v_reg,tail_r_sv2v_reg,head_r_sv2v_reg,empty_r_sv2v_reg;
  assign full_r = full_r_sv2v_reg;
  assign tail_r = tail_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign empty_r = empty_r_sv2v_reg;

  bsg_mem_1r1w
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign _0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_param_o = ~full_r;
  assign enq_i = v_i & N5;
  assign N5 = ~full_r;
  assign N1 = enq_i;
  assign N0 = ~tail_r;
  assign N2 = ~head_r;
  assign N3 = N7 | N9;
  assign N7 = empty_r & N6;
  assign N6 = ~enq_i;
  assign N9 = N8 & N6;
  assign N8 = N5 & yumi_i;
  assign N4 = N13 | N14;
  assign N13 = N11 & N12;
  assign N11 = N10 & enq_i;
  assign N10 = ~empty_r;
  assign N12 = ~yumi_i;
  assign N14 = full_r & N12;

  always @(posedge clk_i) begin
    if(reset_i) begin
      full_r_sv2v_reg <= 1'b0;
      empty_r_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      full_r_sv2v_reg <= N4;
      empty_r_sv2v_reg <= N3;
    end 
    if(reset_i) begin
      tail_r_sv2v_reg <= 1'b0;
    end else if(N1) begin
      tail_r_sv2v_reg <= N0;
    end 
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bp_me_stream_gearbox_00_00000080_00000080_0000000e_6
(
  clk_i,
  reset_i,
  msg_header_i,
  msg_data_i,
  msg_v_i,
  msg_ready_and_o,
  msg_header_o,
  msg_data_o,
  msg_v_o,
  msg_ready_param_i
);

  input [64:0] msg_header_i;
  input [127:0] msg_data_i;
  output [64:0] msg_header_o;
  output [127:0] msg_data_o;
  input clk_i;
  input reset_i;
  input msg_v_i;
  input msg_ready_param_i;
  output msg_ready_and_o;
  output msg_v_o;
  wire [64:0] msg_header_o;
  wire [127:0] msg_data_o;
  wire msg_ready_and_o,msg_v_o,_2_net_;

  bsg_two_fifo_000000c1
  fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_param_o(msg_ready_and_o),
    .data_i({ msg_header_i, msg_data_i }),
    .v_i(msg_v_i),
    .v_o(msg_v_o),
    .data_o({ msg_header_o, msg_data_o }),
    .yumi_i(_2_net_)
  );

  assign _2_net_ = msg_ready_param_i & msg_v_o;

endmodule



module bsg_counter_set_en_3_0
(
  clk_i,
  reset_i,
  set_i,
  en_i,
  val_i,
  count_o
);

  input [1:0] val_i;
  output [1:0] count_o;
  input clk_i;
  input reset_i;
  input set_i;
  input en_i;
  wire [1:0] count_o;
  wire N0,N1,N4,N5,N6,N8,N9,N10,N11,N12,N13,N2,N3,N7;
  reg count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign { N5, N4 } = count_o + 1'b1;
  assign N8 = (N0)? 1'b1 : 
              (N7)? 1'b1 : 
              (N3)? 1'b0 : 1'b0;
  assign N0 = set_i;
  assign { N9, N6 } = (N0)? val_i : 
                      (N7)? { N5, N4 } : 1'b0;
  assign N1 = N13;
  assign N10 = ~reset_i;
  assign N11 = ~set_i;
  assign N12 = N10 & N11;
  assign N13 = en_i & N12;
  assign N2 = en_i | set_i;
  assign N3 = ~N2;
  assign N7 = en_i & N11;

  always @(posedge clk_i) begin
    if(reset_i) begin
      count_o_1_sv2v_reg <= 1'b0;
      count_o_0_sv2v_reg <= 1'b0;
    end else if(N8) begin
      count_o_1_sv2v_reg <= N9;
      count_o_0_sv2v_reg <= N6;
    end 
  end


endmodule



module bsg_mux_segmented_00000002_1
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [1:0] data0_i;
  input [1:0] data1_i;
  input [1:0] sel_i;
  output [1:0] data_o;
  wire [1:0] data_o;
  wire N0,N1,N2,N3;
  assign data_o[0] = (N0)? data1_i[0] : 
                     (N2)? data0_i[0] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[1] = (N1)? data1_i[1] : 
                     (N3)? data0_i[1] : 1'b0;
  assign N1 = sel_i[1];
  assign N2 = ~sel_i[0];
  assign N3 = ~sel_i[1];

endmodule



module bsg_mux_bitwise_00000002
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [1:0] data0_i;
  input [1:0] data1_i;
  input [1:0] sel_i;
  output [1:0] data_o;
  wire [1:0] data_o;

  bsg_mux_segmented_00000002_1
  mux_segmented
  (
    .data0_i(data0_i),
    .data1_i(data1_i),
    .sel_i(sel_i),
    .data_o(data_o)
  );


endmodule



module bp_me_stream_pump_control_00_0000000e_00000080_7_00000006
(
  clk_i,
  reset_i,
  header_i,
  ack_i,
  addr_o,
  first_o,
  critical_o,
  last_o
);

  input [64:0] header_i;
  output [39:0] addr_o;
  input clk_i;
  input reset_i;
  input ack_i;
  output first_o;
  output critical_o;
  output last_o;
  wire [39:0] addr_o,\nz.req_mask ,\nz.addr_mask ,\nz.beat_mask ,\nz.final_mask ;
  wire first_o,critical_o,last_o,N0,N1,N2,N3,N4,N5,N10,N11,N12,N13,N14,\nz.state_r ,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,\nz.stream ,N25,N26,N27,N28,N29,N30,N31,
  N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,\nz.state_n ,N43,N44,N6,N7,N8,N9,N46,
  N47,N48,N49,N50,N51,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4;
  wire [1:0] \nz.stream_size ,\nz.size_li ,\nz.last_cnt ,\nz.cnt_val_li ,\nz.cnt_r ,
  \nz.cnt_lo ,\nz.wrap_lo ,\nz.wrap_cnt ;
  wire [5:4] \nz.base_addr ,\nz.critical_addr ;
  wire [0:0] \nz.wrap_sel_li ;
  reg \nz.state_r_sv2v_reg ;
  assign \nz.state_r  = \nz.state_r_sv2v_reg ;
  assign N19 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N18, N17, N16, N15 } > 1'b1;
  assign N35 = \nz.req_mask  > { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign N37 = \nz.addr_mask  > \nz.beat_mask ;

  bsg_counter_set_en_3_0
  \nz.counter 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .set_i(first_o),
    .en_i(ack_i),
    .val_i(\nz.cnt_val_li ),
    .count_o(\nz.cnt_r )
  );

  assign critical_o = \nz.critical_addr  == \nz.cnt_lo ;
  assign last_o = \nz.last_cnt  == \nz.cnt_lo ;

  bsg_mux_bitwise_00000002
  \nz.wrap_mux 
  (
    .data0_i(\nz.base_addr ),
    .data1_i(\nz.cnt_lo ),
    .sel_i({ \nz.size_li [1:1], \nz.wrap_sel_li [0:0] }),
    .data_o(\nz.wrap_lo )
  );

  assign first_o = ~\nz.state_r ;
  assign { N22, N21, sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << header_i[50:48];
  assign { N18, N17, N16, N15, N9, N8, N7, N6 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << header_i[50:48];
  assign { N34, N33, N32, N31, N30, N29, N28, N27, N26 } = { N18, N17, N16, N15, N9, N8, N7, N6 } - 1'b1;
  assign \nz.stream_size  = { N24, N23 } - 1'b1;
  assign \nz.last_cnt  = \nz.base_addr  + \nz.size_li ;
  assign \nz.cnt_val_li  = \nz.base_addr  + ack_i;
  assign { N24, N23 } = (N0)? { N22, N21 } : 
                        (N20)? { 1'b0, 1'b1 } : 1'b0;
  assign N0 = N19;
  assign \nz.size_li  = (N1)? \nz.stream_size  : 
                        (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = \nz.stream ;
  assign N2 = N25;
  assign \nz.addr_mask  = (N3)? \nz.req_mask  : 
                          (N36)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N3 = N35;
  assign \nz.final_mask  = (N4)? \nz.addr_mask  : 
                           (N38)? \nz.beat_mask  : 1'b0;
  assign N4 = N37;
  assign \nz.cnt_lo  = (N5)? \nz.base_addr  : 
                       (N10)? \nz.cnt_r  : 1'b0;
  assign N5 = N40;
  assign N10 = N39;
  assign \nz.wrap_cnt  = (N5)? \nz.base_addr  : 
                         (N10)? \nz.wrap_lo  : 1'b0;
  assign N43 = ~N42;
  assign \nz.state_n  = (N11)? N43 : 
                        (N12)? N44 : 1'b0;
  assign N11 = \nz.state_r ;
  assign N12 = N41;
  assign N46 = ~header_i[0];
  assign N47 = ~header_i[1];
  assign N48 = header_i[1] & N46;
  assign N49 = N47 | N48;
  assign N50 = N13 & N49;
  assign N13 = ~header_i[2];
  assign \nz.stream  = N14 & N50;
  assign N14 = ~header_i[3];
  assign N20 = ~N19;
  assign N25 = ~\nz.stream ;
  assign \nz.req_mask [39] = ~N34;
  assign \nz.req_mask [38] = ~N34;
  assign \nz.req_mask [37] = ~N34;
  assign \nz.req_mask [36] = ~N34;
  assign \nz.req_mask [35] = ~N34;
  assign \nz.req_mask [34] = ~N34;
  assign \nz.req_mask [33] = ~N34;
  assign \nz.req_mask [32] = ~N34;
  assign \nz.req_mask [31] = ~N34;
  assign \nz.req_mask [30] = ~N34;
  assign \nz.req_mask [29] = ~N34;
  assign \nz.req_mask [28] = ~N34;
  assign \nz.req_mask [27] = ~N34;
  assign \nz.req_mask [26] = ~N34;
  assign \nz.req_mask [25] = ~N34;
  assign \nz.req_mask [24] = ~N34;
  assign \nz.req_mask [23] = ~N34;
  assign \nz.req_mask [22] = ~N34;
  assign \nz.req_mask [21] = ~N34;
  assign \nz.req_mask [20] = ~N34;
  assign \nz.req_mask [19] = ~N34;
  assign \nz.req_mask [18] = ~N34;
  assign \nz.req_mask [17] = ~N34;
  assign \nz.req_mask [16] = ~N34;
  assign \nz.req_mask [15] = ~N34;
  assign \nz.req_mask [14] = ~N34;
  assign \nz.req_mask [13] = ~N34;
  assign \nz.req_mask [12] = ~N34;
  assign \nz.req_mask [11] = ~N34;
  assign \nz.req_mask [10] = ~N34;
  assign \nz.req_mask [9] = ~N34;
  assign \nz.req_mask [8] = ~N34;
  assign \nz.req_mask [7] = ~N33;
  assign \nz.req_mask [6] = ~N32;
  assign \nz.req_mask [5] = ~N31;
  assign \nz.req_mask [4] = ~N30;
  assign \nz.req_mask [3] = ~N29;
  assign \nz.req_mask [2] = ~N28;
  assign \nz.req_mask [1] = ~N27;
  assign \nz.req_mask [0] = ~N26;
  assign N36 = ~N35;
  assign \nz.beat_mask [39] = ~1'b0;
  assign \nz.beat_mask [38] = ~1'b0;
  assign \nz.beat_mask [37] = ~1'b0;
  assign \nz.beat_mask [36] = ~1'b0;
  assign \nz.beat_mask [35] = ~1'b0;
  assign \nz.beat_mask [34] = ~1'b0;
  assign \nz.beat_mask [33] = ~1'b0;
  assign \nz.beat_mask [32] = ~1'b0;
  assign \nz.beat_mask [31] = ~1'b0;
  assign \nz.beat_mask [30] = ~1'b0;
  assign \nz.beat_mask [29] = ~1'b0;
  assign \nz.beat_mask [28] = ~1'b0;
  assign \nz.beat_mask [27] = ~1'b0;
  assign \nz.beat_mask [26] = ~1'b0;
  assign \nz.beat_mask [25] = ~1'b0;
  assign \nz.beat_mask [24] = ~1'b0;
  assign \nz.beat_mask [23] = ~1'b0;
  assign \nz.beat_mask [22] = ~1'b0;
  assign \nz.beat_mask [21] = ~1'b0;
  assign \nz.beat_mask [20] = ~1'b0;
  assign \nz.beat_mask [19] = ~1'b0;
  assign \nz.beat_mask [18] = ~1'b0;
  assign \nz.beat_mask [17] = ~1'b0;
  assign \nz.beat_mask [16] = ~1'b0;
  assign \nz.beat_mask [15] = ~1'b0;
  assign \nz.beat_mask [14] = ~1'b0;
  assign \nz.beat_mask [13] = ~1'b0;
  assign \nz.beat_mask [12] = ~1'b0;
  assign \nz.beat_mask [11] = ~1'b0;
  assign \nz.beat_mask [10] = ~1'b0;
  assign \nz.beat_mask [9] = ~1'b0;
  assign \nz.beat_mask [8] = ~1'b0;
  assign \nz.beat_mask [7] = ~1'b0;
  assign \nz.beat_mask [6] = ~1'b0;
  assign \nz.beat_mask [5] = ~1'b0;
  assign \nz.beat_mask [4] = ~1'b0;
  assign \nz.beat_mask [3] = ~1'b1;
  assign \nz.beat_mask [2] = ~1'b1;
  assign \nz.beat_mask [1] = ~1'b1;
  assign \nz.beat_mask [0] = ~1'b1;
  assign N38 = ~N37;
  assign \nz.base_addr [5] = header_i[13] & \nz.addr_mask [5];
  assign \nz.base_addr [4] = header_i[12] & \nz.addr_mask [4];
  assign \nz.critical_addr [5] = header_i[13] & \nz.beat_mask [5];
  assign \nz.critical_addr [4] = header_i[12] & \nz.beat_mask [4];
  assign N39 = ~first_o;
  assign N40 = first_o;
  assign \nz.wrap_sel_li [0] = \nz.size_li [1] | \nz.size_li [0];
  assign addr_o[39] = header_i[47] & \nz.final_mask [39];
  assign addr_o[38] = header_i[46] & \nz.final_mask [38];
  assign addr_o[37] = header_i[45] & \nz.final_mask [37];
  assign addr_o[36] = header_i[44] & \nz.final_mask [36];
  assign addr_o[35] = header_i[43] & \nz.final_mask [35];
  assign addr_o[34] = header_i[42] & \nz.final_mask [34];
  assign addr_o[33] = header_i[41] & \nz.final_mask [33];
  assign addr_o[32] = header_i[40] & \nz.final_mask [32];
  assign addr_o[31] = header_i[39] & \nz.final_mask [31];
  assign addr_o[30] = header_i[38] & \nz.final_mask [30];
  assign addr_o[29] = header_i[37] & \nz.final_mask [29];
  assign addr_o[28] = header_i[36] & \nz.final_mask [28];
  assign addr_o[27] = header_i[35] & \nz.final_mask [27];
  assign addr_o[26] = header_i[34] & \nz.final_mask [26];
  assign addr_o[25] = header_i[33] & \nz.final_mask [25];
  assign addr_o[24] = header_i[32] & \nz.final_mask [24];
  assign addr_o[23] = header_i[31] & \nz.final_mask [23];
  assign addr_o[22] = header_i[30] & \nz.final_mask [22];
  assign addr_o[21] = header_i[29] & \nz.final_mask [21];
  assign addr_o[20] = header_i[28] & \nz.final_mask [20];
  assign addr_o[19] = header_i[27] & \nz.final_mask [19];
  assign addr_o[18] = header_i[26] & \nz.final_mask [18];
  assign addr_o[17] = header_i[25] & \nz.final_mask [17];
  assign addr_o[16] = header_i[24] & \nz.final_mask [16];
  assign addr_o[15] = header_i[23] & \nz.final_mask [15];
  assign addr_o[14] = header_i[22] & \nz.final_mask [14];
  assign addr_o[13] = header_i[21] & \nz.final_mask [13];
  assign addr_o[12] = header_i[20] & \nz.final_mask [12];
  assign addr_o[11] = header_i[19] & \nz.final_mask [11];
  assign addr_o[10] = header_i[18] & \nz.final_mask [10];
  assign addr_o[9] = header_i[17] & \nz.final_mask [9];
  assign addr_o[8] = header_i[16] & \nz.final_mask [8];
  assign addr_o[7] = header_i[15] & \nz.final_mask [7];
  assign addr_o[6] = header_i[14] & \nz.final_mask [6];
  assign addr_o[5] = \nz.wrap_cnt [1] & \nz.final_mask [5];
  assign addr_o[4] = \nz.wrap_cnt [0] & \nz.final_mask [4];
  assign addr_o[3] = header_i[11] & \nz.final_mask [3];
  assign addr_o[2] = header_i[10] & \nz.final_mask [2];
  assign addr_o[1] = header_i[9] & \nz.final_mask [1];
  assign addr_o[0] = header_i[8] & \nz.final_mask [0];
  assign N41 = first_o;
  assign N42 = ack_i & last_o;
  assign N44 = ack_i & N51;
  assign N51 = ~last_o;

  always @(posedge clk_i) begin
    if(reset_i) begin
      \nz.state_r_sv2v_reg  <= 1'b0;
    end else if(1'b1) begin
      \nz.state_r_sv2v_reg  <= \nz.state_n ;
    end 
  end


endmodule



module bp_me_stream_pump_in_00_00000080_0000000e_6_7
(
  clk_i,
  reset_i,
  msg_header_i,
  msg_data_i,
  msg_v_i,
  msg_ready_and_o,
  fsm_header_o,
  fsm_data_o,
  fsm_v_o,
  fsm_yumi_i,
  fsm_addr_o,
  fsm_new_o,
  fsm_critical_o,
  fsm_last_o
);

  input [64:0] msg_header_i;
  input [127:0] msg_data_i;
  output [64:0] fsm_header_o;
  output [127:0] fsm_data_o;
  output [39:0] fsm_addr_o;
  input clk_i;
  input reset_i;
  input msg_v_i;
  input fsm_yumi_i;
  output msg_ready_and_o;
  output fsm_v_o;
  output fsm_new_o;
  output fsm_critical_o;
  output fsm_last_o;
  wire [64:0] fsm_header_o;
  wire [127:0] fsm_data_o;
  wire [39:0] fsm_addr_o;
  wire msg_ready_and_o,fsm_v_o,fsm_new_o,fsm_critical_o,fsm_last_o,N0,N1,msg_yumi_lo,
  N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,nz_stream,fsm_stream,msg_stream,N12,N13,N14,N15,
  N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,
  N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,
  sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8;
  wire [1:0] stream_size;

  bp_me_stream_gearbox_00_00000080_00000080_0000000e_6
  gearbox
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .msg_header_i(msg_header_i),
    .msg_data_i(msg_data_i),
    .msg_v_i(msg_v_i),
    .msg_ready_and_o(msg_ready_and_o),
    .msg_header_o(fsm_header_o),
    .msg_data_o(fsm_data_o),
    .msg_v_o(fsm_v_o),
    .msg_ready_param_i(msg_yumi_lo)
  );

  assign N6 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N5, N4, N3, N2 } > 1'b1;
  assign nz_stream = stream_size > 1'b0;

  bp_me_stream_pump_control_00_0000000e_00000080_7_00000006
  pump_control
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .header_i(fsm_header_o),
    .ack_i(fsm_yumi_i),
    .addr_o(fsm_addr_o),
    .first_o(fsm_new_o),
    .critical_o(fsm_critical_o),
    .last_o(fsm_last_o)
  );

  assign { N9, N8, sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fsm_header_o[50:48];
  assign { N5, N4, N3, N2, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fsm_header_o[50:48];
  assign stream_size = { N11, N10 } - 1'b1;
  assign { N11, N10 } = (N0)? { N9, N8 } : 
                        (N7)? { 1'b0, 1'b1 } : 1'b0;
  assign N0 = N6;
  assign msg_yumi_lo = (N1)? N14 : 
                       (N13)? fsm_yumi_i : 1'b0;
  assign N1 = N12;
  assign msg_stream = (N31)? 1'b0 : 
                      (N33)? 1'b1 : 
                      (N35)? 1'b1 : 
                      (N37)? 1'b0 : 
                      (N39)? 1'b0 : 
                      (N41)? 1'b0 : 
                      (N43)? 1'b0 : 
                      (N45)? 1'b0 : 
                      (N32)? 1'b0 : 
                      (N34)? 1'b0 : 
                      (N36)? 1'b0 : 
                      (N38)? 1'b0 : 
                      (N40)? 1'b0 : 
                      (N42)? 1'b0 : 
                      (N44)? 1'b0 : 
                      (N46)? 1'b0 : 1'b0;
  assign fsm_stream = (N31)? 1'b1 : 
                      (N33)? 1'b1 : 
                      (N35)? 1'b1 : 
                      (N37)? 1'b0 : 
                      (N39)? 1'b0 : 
                      (N41)? 1'b0 : 
                      (N43)? 1'b0 : 
                      (N45)? 1'b0 : 
                      (N32)? 1'b0 : 
                      (N34)? 1'b0 : 
                      (N36)? 1'b0 : 
                      (N38)? 1'b0 : 
                      (N40)? 1'b0 : 
                      (N42)? 1'b0 : 
                      (N44)? 1'b0 : 
                      (N46)? 1'b0 : 1'b0;
  assign N7 = ~N6;
  assign N12 = N48 & nz_stream;
  assign N48 = N47 & fsm_stream;
  assign N47 = ~msg_stream;
  assign N13 = ~N12;
  assign N14 = fsm_last_o & fsm_yumi_i;
  assign N15 = ~fsm_header_o[0];
  assign N16 = ~fsm_header_o[1];
  assign N17 = N15 & N16;
  assign N18 = N15 & fsm_header_o[1];
  assign N19 = fsm_header_o[0] & N16;
  assign N20 = fsm_header_o[0] & fsm_header_o[1];
  assign N21 = ~fsm_header_o[2];
  assign N22 = N17 & N21;
  assign N23 = N17 & fsm_header_o[2];
  assign N24 = N19 & N21;
  assign N25 = N19 & fsm_header_o[2];
  assign N26 = N18 & N21;
  assign N27 = N18 & fsm_header_o[2];
  assign N28 = N20 & N21;
  assign N29 = N20 & fsm_header_o[2];
  assign N30 = ~fsm_header_o[3];
  assign N31 = N22 & N30;
  assign N32 = N22 & fsm_header_o[3];
  assign N33 = N24 & N30;
  assign N34 = N24 & fsm_header_o[3];
  assign N35 = N26 & N30;
  assign N36 = N26 & fsm_header_o[3];
  assign N37 = N28 & N30;
  assign N38 = N28 & fsm_header_o[3];
  assign N39 = N23 & N30;
  assign N40 = N23 & fsm_header_o[3];
  assign N41 = N25 & N30;
  assign N42 = N25 & fsm_header_o[3];
  assign N43 = N27 & N30;
  assign N44 = N27 & fsm_header_o[3];
  assign N45 = N29 & N30;
  assign N46 = N29 & fsm_header_o[3];

endmodule



module bp_me_stream_gearbox_00_00000080_00000080_0000000e_5
(
  clk_i,
  reset_i,
  msg_header_i,
  msg_data_i,
  msg_v_i,
  msg_ready_and_o,
  msg_header_o,
  msg_data_o,
  msg_v_o,
  msg_ready_param_i
);

  input [64:0] msg_header_i;
  input [127:0] msg_data_i;
  output [64:0] msg_header_o;
  output [127:0] msg_data_o;
  input clk_i;
  input reset_i;
  input msg_v_i;
  input msg_ready_param_i;
  output msg_ready_and_o;
  output msg_v_o;
  wire [64:0] msg_header_o;
  wire [127:0] msg_data_o;
  wire msg_ready_and_o,msg_v_o,_2_net_;

  bsg_two_fifo_000000c1
  fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_param_o(msg_ready_and_o),
    .data_i({ msg_header_i, msg_data_i }),
    .v_i(msg_v_i),
    .v_o(msg_v_o),
    .data_o({ msg_header_o, msg_data_o }),
    .yumi_i(_2_net_)
  );

  assign _2_net_ = msg_ready_param_i & msg_v_o;

endmodule



module bp_me_stream_pump_out_00_00000080_0000000e_5_7
(
  clk_i,
  reset_i,
  msg_header_o,
  msg_data_o,
  msg_v_o,
  msg_ready_and_i,
  fsm_header_i,
  fsm_data_i,
  fsm_v_i,
  fsm_ready_then_o,
  fsm_addr_o,
  fsm_new_o,
  fsm_last_o,
  fsm_critical_o
);

  output [64:0] msg_header_o;
  output [127:0] msg_data_o;
  input [64:0] fsm_header_i;
  input [127:0] fsm_data_i;
  output [39:0] fsm_addr_o;
  input clk_i;
  input reset_i;
  input msg_ready_and_i;
  input fsm_v_i;
  output msg_v_o;
  output fsm_ready_then_o;
  output fsm_new_o;
  output fsm_last_o;
  output fsm_critical_o;
  wire [64:0] msg_header_o;
  wire [127:0] msg_data_o;
  wire [39:0] fsm_addr_o;
  wire msg_v_o,fsm_ready_then_o,fsm_new_o,fsm_last_o,fsm_critical_o,N0,N1,N2,N3,N4,N5,
  N6,N7,msg_v_lo,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,nz_stream,fsm_stream,
  msg_stream,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,sv2v_dc_1,sv2v_dc_2,
  sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8;
  wire [1:0] stream_size;

  bp_me_stream_gearbox_00_00000080_00000080_0000000e_5
  gearbox
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .msg_header_i(fsm_header_i),
    .msg_data_i(fsm_data_i),
    .msg_v_i(msg_v_lo),
    .msg_ready_and_o(fsm_ready_then_o),
    .msg_header_o(msg_header_o),
    .msg_data_o(msg_data_o),
    .msg_v_o(msg_v_o),
    .msg_ready_param_i(msg_ready_and_i)
  );

  assign N12 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N11, N10, N9, N8 } > 1'b1;
  assign nz_stream = stream_size > 1'b0;

  bp_me_stream_pump_control_00_0000000e_00000080_7_00000006
  pump_control
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .header_i(fsm_header_i),
    .ack_i(fsm_v_i),
    .addr_o(fsm_addr_o),
    .first_o(fsm_new_o),
    .critical_o(fsm_critical_o),
    .last_o(fsm_last_o)
  );

  assign { N15, N14, sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fsm_header_i[50:48];
  assign { N11, N10, N9, N8, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fsm_header_i[50:48];
  assign stream_size = { N17, N16 } - 1'b1;
  assign { N17, N16 } = (N0)? { N15, N14 } : 
                        (N13)? { 1'b0, 1'b1 } : 1'b0;
  assign N0 = N12;
  assign msg_v_lo = (N1)? N20 : 
                    (N19)? fsm_v_i : 1'b0;
  assign N1 = N18;
  assign N21 = ~fsm_header_i[0];
  assign N22 = N2 & N21;
  assign N2 = ~fsm_header_i[2];
  assign msg_stream = N3 & N22;
  assign N3 = ~fsm_header_i[3];
  assign N23 = ~fsm_header_i[1];
  assign N24 = N4 & N23;
  assign N4 = ~fsm_header_i[2];
  assign N25 = N5 & N24;
  assign N5 = ~fsm_header_i[3];
  assign N26 = ~fsm_header_i[0];
  assign N27 = N6 & N26;
  assign N6 = ~fsm_header_i[2];
  assign N28 = N7 & N27;
  assign N7 = ~fsm_header_i[3];
  assign fsm_stream = N25 | N28;
  assign N13 = ~N12;
  assign N18 = N30 & nz_stream;
  assign N30 = fsm_stream & N29;
  assign N29 = ~msg_stream;
  assign N19 = ~N18;
  assign N20 = fsm_v_i & fsm_new_o;

endmodule



module bsg_circular_ptr_00000006_1
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [0:0] add_i;
  output [2:0] o;
  output [2:0] n_o;
  input clk;
  input reset_i;
  wire [2:0] o,n_o,ptr_nowrap;
  wire N0,N1,N2,N3,N4,N5,N6;
  wire [3:0] ptr_wrap;
  reg o_2_sv2v_reg,o_1_sv2v_reg,o_0_sv2v_reg;
  assign o[2] = o_2_sv2v_reg;
  assign o[1] = o_1_sv2v_reg;
  assign o[0] = o_0_sv2v_reg;
  assign ptr_nowrap = o + add_i[0];
  assign { N5, N4, N3, N2 } = o - { 1'b1, 1'b1, 1'b0 };
  assign ptr_wrap = { N5, N4, N3, N2 } + add_i[0];
  assign n_o = (N0)? ptr_wrap[2:0] : 
               (N1)? ptr_nowrap : 1'b0;
  assign N0 = N6;
  assign N1 = ptr_wrap[3];
  assign N6 = ~ptr_wrap[3];

  always @(posedge clk) begin
    if(reset_i) begin
      o_2_sv2v_reg <= 1'b0;
      o_1_sv2v_reg <= 1'b0;
      o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      o_2_sv2v_reg <= n_o[2];
      o_1_sv2v_reg <= n_o[1];
      o_0_sv2v_reg <= n_o[0];
    end 
  end


endmodule



module bsg_fifo_tracker_00000006
(
  clk_i,
  reset_i,
  enq_i,
  deq_i,
  wptr_r_o,
  rptr_r_o,
  rptr_n_o,
  full_o,
  empty_o
);

  output [2:0] wptr_r_o;
  output [2:0] rptr_r_o;
  output [2:0] rptr_n_o;
  input clk_i;
  input reset_i;
  input enq_i;
  input deq_i;
  output full_o;
  output empty_o;
  wire [2:0] wptr_r_o,rptr_r_o,rptr_n_o;
  wire full_o,empty_o,enq_r,deq_r,N0,equal_ptrs,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3;
  reg deq_r_sv2v_reg,enq_r_sv2v_reg;
  assign deq_r = deq_r_sv2v_reg;
  assign enq_r = enq_r_sv2v_reg;

  bsg_circular_ptr_00000006_1
  rptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(deq_i),
    .o(rptr_r_o),
    .n_o(rptr_n_o)
  );


  bsg_circular_ptr_00000006_1
  wptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(enq_i),
    .o(wptr_r_o),
    .n_o({ sv2v_dc_1, sv2v_dc_2, sv2v_dc_3 })
  );

  assign equal_ptrs = rptr_r_o == wptr_r_o;
  assign N0 = enq_i | deq_i;
  assign empty_o = equal_ptrs & deq_r;
  assign full_o = equal_ptrs & enq_r;

  always @(posedge clk_i) begin
    if(reset_i) begin
      deq_r_sv2v_reg <= 1'b1;
      enq_r_sv2v_reg <= 1'b0;
    end else if(N0) begin
      deq_r_sv2v_reg <= deq_i;
      enq_r_sv2v_reg <= enq_i;
    end 
  end


endmodule



module bsg_fifo_1r1w_small_unhardened_00000042_00000006_1
(
  clk_i,
  reset_i,
  v_i,
  ready_param_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [65:0] data_i;
  output [65:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_param_o;
  output v_o;
  wire [65:0] data_o;
  wire ready_param_o,v_o,full,empty,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3;
  wire [2:0] wptr_r,rptr_r;

  bsg_fifo_tracker_00000006
  ft
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .enq_i(v_i),
    .deq_i(yumi_i),
    .wptr_r_o(wptr_r),
    .rptr_r_o(rptr_r),
    .rptr_n_o({ sv2v_dc_1, sv2v_dc_2, sv2v_dc_3 }),
    .full_o(full),
    .empty_o(empty)
  );


  bsg_mem_1r1w
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(v_i),
    .w_addr_i(wptr_r),
    .w_data_i(data_i),
    .r_v_i(v_o),
    .r_addr_i(rptr_r),
    .r_data_o(data_o)
  );

  assign ready_param_o = ~full;
  assign v_o = ~empty;

endmodule



module bsg_fifo_1r1w_small_00000042_00000006_1
(
  clk_i,
  reset_i,
  v_i,
  ready_param_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [65:0] data_i;
  output [65:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_param_o;
  output v_o;
  wire [65:0] data_o;
  wire ready_param_o,v_o;

  bsg_fifo_1r1w_small_unhardened_00000042_00000006_1
  \unhardened.un.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_param_o(ready_param_o),
    .data_i(data_i),
    .v_o(v_o),
    .data_o(data_o),
    .yumi_i(yumi_i)
  );


endmodule



module bp_me_stream_pump_00_00000080_0000000e_6_7_00000080_0000000e_5_7_00000042_00000006
(
  clk_i,
  reset_i,
  in_msg_header_i,
  in_msg_data_i,
  in_msg_v_i,
  in_msg_ready_and_o,
  in_fsm_header_o,
  in_fsm_data_o,
  in_fsm_v_o,
  in_fsm_yumi_i,
  in_fsm_metadata_i,
  in_fsm_addr_o,
  in_fsm_new_o,
  in_fsm_critical_o,
  in_fsm_last_o,
  out_msg_header_o,
  out_msg_data_o,
  out_msg_v_o,
  out_msg_ready_and_i,
  out_fsm_header_i,
  out_fsm_data_i,
  out_fsm_v_i,
  out_fsm_ready_then_o,
  out_fsm_metadata_o,
  out_fsm_addr_o,
  out_fsm_new_o,
  out_fsm_last_o,
  out_fsm_critical_o
);

  input [64:0] in_msg_header_i;
  input [127:0] in_msg_data_i;
  output [64:0] in_fsm_header_o;
  output [127:0] in_fsm_data_o;
  input [65:0] in_fsm_metadata_i;
  output [39:0] in_fsm_addr_o;
  output [64:0] out_msg_header_o;
  output [127:0] out_msg_data_o;
  input [64:0] out_fsm_header_i;
  input [127:0] out_fsm_data_i;
  output [65:0] out_fsm_metadata_o;
  output [39:0] out_fsm_addr_o;
  input clk_i;
  input reset_i;
  input in_msg_v_i;
  input in_fsm_yumi_i;
  input out_msg_ready_and_i;
  input out_fsm_v_i;
  output in_msg_ready_and_o;
  output in_fsm_v_o;
  output in_fsm_new_o;
  output in_fsm_critical_o;
  output in_fsm_last_o;
  output out_msg_v_o;
  output out_fsm_ready_then_o;
  output out_fsm_new_o;
  output out_fsm_last_o;
  output out_fsm_critical_o;
  wire [64:0] in_fsm_header_o,out_msg_header_o;
  wire [127:0] in_fsm_data_o,out_msg_data_o;
  wire [39:0] in_fsm_addr_o,out_fsm_addr_o;
  wire [65:0] out_fsm_metadata_o;
  wire in_msg_ready_and_o,in_fsm_v_o,in_fsm_new_o,in_fsm_critical_o,in_fsm_last_o,
  out_msg_v_o,out_fsm_ready_then_o,out_fsm_new_o,out_fsm_last_o,out_fsm_critical_o,
  in_fsm_v_lo,out_fsm_ready_then_lo,stream_fifo_v_li,stream_fifo_ready_then_lo,
  stream_fifo_v_lo,stream_fifo_yumi_li;

  bp_me_stream_pump_in_00_00000080_0000000e_6_7
  in
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .msg_header_i(in_msg_header_i),
    .msg_data_i(in_msg_data_i),
    .msg_v_i(in_msg_v_i),
    .msg_ready_and_o(in_msg_ready_and_o),
    .fsm_header_o(in_fsm_header_o),
    .fsm_data_o(in_fsm_data_o),
    .fsm_v_o(in_fsm_v_lo),
    .fsm_yumi_i(in_fsm_yumi_i),
    .fsm_addr_o(in_fsm_addr_o),
    .fsm_new_o(in_fsm_new_o),
    .fsm_critical_o(in_fsm_critical_o),
    .fsm_last_o(in_fsm_last_o)
  );


  bp_me_stream_pump_out_00_00000080_0000000e_5_7
  out
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .msg_header_o(out_msg_header_o),
    .msg_data_o(out_msg_data_o),
    .msg_v_o(out_msg_v_o),
    .msg_ready_and_i(out_msg_ready_and_i),
    .fsm_header_i(out_fsm_header_i),
    .fsm_data_i(out_fsm_data_i),
    .fsm_v_i(out_fsm_v_i),
    .fsm_ready_then_o(out_fsm_ready_then_lo),
    .fsm_addr_o(out_fsm_addr_o),
    .fsm_new_o(out_fsm_new_o),
    .fsm_last_o(out_fsm_last_o),
    .fsm_critical_o(out_fsm_critical_o)
  );


  bsg_fifo_1r1w_small_00000042_00000006_1
  stream_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(stream_fifo_v_li),
    .ready_param_o(stream_fifo_ready_then_lo),
    .data_i(in_fsm_metadata_i),
    .v_o(stream_fifo_v_lo),
    .data_o(out_fsm_metadata_o),
    .yumi_i(stream_fifo_yumi_li)
  );

  assign in_fsm_v_o = in_fsm_v_lo & stream_fifo_ready_then_lo;
  assign stream_fifo_v_li = in_fsm_yumi_i & in_fsm_new_o;
  assign out_fsm_ready_then_o = out_fsm_ready_then_lo & stream_fifo_v_lo;
  assign stream_fifo_yumi_li = out_fsm_v_i & out_fsm_last_o;

endmodule



module bsg_counter_clear_up_000007ff_0
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [10:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire [10:0] count_o;
  wire N0,N1,N4,N5,N6,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N2,
  N3,N7,N30,N24;
  reg count_o_10_sv2v_reg,count_o_9_sv2v_reg,count_o_8_sv2v_reg,count_o_7_sv2v_reg,
  count_o_6_sv2v_reg,count_o_5_sv2v_reg,count_o_4_sv2v_reg,count_o_3_sv2v_reg,
  count_o_2_sv2v_reg,count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[10] = count_o_10_sv2v_reg;
  assign count_o[9] = count_o_9_sv2v_reg;
  assign count_o[8] = count_o_8_sv2v_reg;
  assign count_o[7] = count_o_7_sv2v_reg;
  assign count_o[6] = count_o_6_sv2v_reg;
  assign count_o[5] = count_o_5_sv2v_reg;
  assign count_o[4] = count_o_4_sv2v_reg;
  assign count_o[3] = count_o_3_sv2v_reg;
  assign count_o[2] = count_o_2_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign N24 = reset_i | clear_i;
  assign { N16, N15, N14, N13, N12, N11, N10, N9, N8, N6, N5 } = count_o + 1'b1;
  assign N17 = (N0)? 1'b1 : 
               (N7)? 1'b1 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = clear_i;
  assign N19 = (N1)? 1'b1 : 
               (N30)? 1'b0 : 1'b0;
  assign N1 = up_i;
  assign N18 = (N0)? up_i : 
               (N7)? N5 : 1'b0;
  assign N4 = N23;
  assign N20 = ~reset_i;
  assign N21 = ~clear_i;
  assign N22 = N20 & N21;
  assign N23 = up_i & N22;
  assign N2 = up_i | clear_i;
  assign N3 = ~N2;
  assign N7 = up_i & N21;
  assign N30 = ~up_i;

  always @(posedge clk_i) begin
    if(N24) begin
      count_o_10_sv2v_reg <= 1'b0;
      count_o_9_sv2v_reg <= 1'b0;
      count_o_8_sv2v_reg <= 1'b0;
      count_o_7_sv2v_reg <= 1'b0;
      count_o_6_sv2v_reg <= 1'b0;
      count_o_5_sv2v_reg <= 1'b0;
      count_o_4_sv2v_reg <= 1'b0;
      count_o_3_sv2v_reg <= 1'b0;
      count_o_2_sv2v_reg <= 1'b0;
      count_o_1_sv2v_reg <= 1'b0;
    end else if(N19) begin
      count_o_10_sv2v_reg <= N16;
      count_o_9_sv2v_reg <= N15;
      count_o_8_sv2v_reg <= N14;
      count_o_7_sv2v_reg <= N13;
      count_o_6_sv2v_reg <= N12;
      count_o_5_sv2v_reg <= N11;
      count_o_4_sv2v_reg <= N10;
      count_o_3_sv2v_reg <= N9;
      count_o_2_sv2v_reg <= N8;
      count_o_1_sv2v_reg <= N6;
    end 
    if(reset_i) begin
      count_o_0_sv2v_reg <= 1'b0;
    end else if(N17) begin
      count_o_0_sv2v_reg <= N18;
    end 
  end


endmodule



module bsg_expand_bitmask_00000010_1
(
  i,
  o
);

  input [15:0] i;
  output [15:0] o;
  wire [15:0] o;
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_expand_bitmask_00000008_2
(
  i,
  o
);

  input [7:0] i;
  output [15:0] o;
  wire [15:0] o;
  wire o_15_,o_13_,o_11_,o_9_,o_7_,o_5_,o_3_,o_1_;
  assign o_15_ = i[7];
  assign o[14] = o_15_;
  assign o[15] = o_15_;
  assign o_13_ = i[6];
  assign o[12] = o_13_;
  assign o[13] = o_13_;
  assign o_11_ = i[5];
  assign o[10] = o_11_;
  assign o[11] = o_11_;
  assign o_9_ = i[4];
  assign o[8] = o_9_;
  assign o[9] = o_9_;
  assign o_7_ = i[3];
  assign o[6] = o_7_;
  assign o[7] = o_7_;
  assign o_5_ = i[2];
  assign o[4] = o_5_;
  assign o[5] = o_5_;
  assign o_3_ = i[1];
  assign o[2] = o_3_;
  assign o[3] = o_3_;
  assign o_1_ = i[0];
  assign o[0] = o_1_;
  assign o[1] = o_1_;

endmodule



module bsg_expand_bitmask_00000004_4
(
  i,
  o
);

  input [3:0] i;
  output [15:0] o;
  wire [15:0] o;
  wire o_15_,o_11_,o_7_,o_3_;
  assign o_15_ = i[3];
  assign o[12] = o_15_;
  assign o[13] = o_15_;
  assign o[14] = o_15_;
  assign o[15] = o_15_;
  assign o_11_ = i[2];
  assign o[8] = o_11_;
  assign o[9] = o_11_;
  assign o[10] = o_11_;
  assign o[11] = o_11_;
  assign o_7_ = i[1];
  assign o[4] = o_7_;
  assign o[5] = o_7_;
  assign o[6] = o_7_;
  assign o[7] = o_7_;
  assign o_3_ = i[0];
  assign o[0] = o_3_;
  assign o[1] = o_3_;
  assign o[2] = o_3_;
  assign o[3] = o_3_;

endmodule



module bsg_expand_bitmask_00000002_8
(
  i,
  o
);

  input [1:0] i;
  output [15:0] o;
  wire [15:0] o;
  wire o_15_,o_7_;
  assign o_15_ = i[1];
  assign o[8] = o_15_;
  assign o[9] = o_15_;
  assign o[10] = o_15_;
  assign o[11] = o_15_;
  assign o[12] = o_15_;
  assign o[13] = o_15_;
  assign o[14] = o_15_;
  assign o[15] = o_15_;
  assign o_7_ = i[0];
  assign o[0] = o_7_;
  assign o[1] = o_7_;
  assign o[2] = o_7_;
  assign o[3] = o_7_;
  assign o[4] = o_7_;
  assign o[5] = o_7_;
  assign o[6] = o_7_;
  assign o[7] = o_7_;

endmodule



module bsg_mux_00000010_00000005
(
  data_i,
  sel_i,
  data_o
);

  input [79:0] data_i;
  input [2:0] sel_i;
  output [15:0] data_o;
  wire [15:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;
  assign N10 = N0 & N1 & N2;
  assign N0 = ~sel_i[2];
  assign N1 = ~sel_i[0];
  assign N2 = ~sel_i[1];
  assign N11 = sel_i[0] & N3;
  assign N3 = ~sel_i[1];
  assign N12 = N4 & sel_i[1];
  assign N4 = ~sel_i[0];
  assign N13 = sel_i[0] & sel_i[1];
  assign data_o[15] = (N5)? data_i[15] : 
                      (N6)? data_i[31] : 
                      (N7)? data_i[47] : 
                      (N8)? data_i[63] : 
                      (N9)? data_i[79] : 1'b0;
  assign N5 = N10;
  assign N6 = N11;
  assign N7 = N12;
  assign N8 = N13;
  assign N9 = sel_i[2];
  assign data_o[14] = (N5)? data_i[14] : 
                      (N6)? data_i[30] : 
                      (N7)? data_i[46] : 
                      (N8)? data_i[62] : 
                      (N9)? data_i[78] : 1'b0;
  assign data_o[13] = (N5)? data_i[13] : 
                      (N6)? data_i[29] : 
                      (N7)? data_i[45] : 
                      (N8)? data_i[61] : 
                      (N9)? data_i[77] : 1'b0;
  assign data_o[12] = (N5)? data_i[12] : 
                      (N6)? data_i[28] : 
                      (N7)? data_i[44] : 
                      (N8)? data_i[60] : 
                      (N9)? data_i[76] : 1'b0;
  assign data_o[11] = (N5)? data_i[11] : 
                      (N6)? data_i[27] : 
                      (N7)? data_i[43] : 
                      (N8)? data_i[59] : 
                      (N9)? data_i[75] : 1'b0;
  assign data_o[10] = (N5)? data_i[10] : 
                      (N6)? data_i[26] : 
                      (N7)? data_i[42] : 
                      (N8)? data_i[58] : 
                      (N9)? data_i[74] : 1'b0;
  assign data_o[9] = (N5)? data_i[9] : 
                     (N6)? data_i[25] : 
                     (N7)? data_i[41] : 
                     (N8)? data_i[57] : 
                     (N9)? data_i[73] : 1'b0;
  assign data_o[8] = (N5)? data_i[8] : 
                     (N6)? data_i[24] : 
                     (N7)? data_i[40] : 
                     (N8)? data_i[56] : 
                     (N9)? data_i[72] : 1'b0;
  assign data_o[7] = (N5)? data_i[7] : 
                     (N6)? data_i[23] : 
                     (N7)? data_i[39] : 
                     (N8)? data_i[55] : 
                     (N9)? data_i[71] : 1'b0;
  assign data_o[6] = (N5)? data_i[6] : 
                     (N6)? data_i[22] : 
                     (N7)? data_i[38] : 
                     (N8)? data_i[54] : 
                     (N9)? data_i[70] : 1'b0;
  assign data_o[5] = (N5)? data_i[5] : 
                     (N6)? data_i[21] : 
                     (N7)? data_i[37] : 
                     (N8)? data_i[53] : 
                     (N9)? data_i[69] : 1'b0;
  assign data_o[4] = (N5)? data_i[4] : 
                     (N6)? data_i[20] : 
                     (N7)? data_i[36] : 
                     (N8)? data_i[52] : 
                     (N9)? data_i[68] : 1'b0;
  assign data_o[3] = (N5)? data_i[3] : 
                     (N6)? data_i[19] : 
                     (N7)? data_i[35] : 
                     (N8)? data_i[51] : 
                     (N9)? data_i[67] : 1'b0;
  assign data_o[2] = (N5)? data_i[2] : 
                     (N6)? data_i[18] : 
                     (N7)? data_i[34] : 
                     (N8)? data_i[50] : 
                     (N9)? data_i[66] : 1'b0;
  assign data_o[1] = (N5)? data_i[1] : 
                     (N6)? data_i[17] : 
                     (N7)? data_i[33] : 
                     (N8)? data_i[49] : 
                     (N9)? data_i[65] : 1'b0;
  assign data_o[0] = (N5)? data_i[0] : 
                     (N6)? data_i[16] : 
                     (N7)? data_i[32] : 
                     (N8)? data_i[48] : 
                     (N9)? data_i[64] : 1'b0;

endmodule



module bp_me_dram_hash_encode_00
(
  paddr_i,
  data_i,
  dram_o,
  daddr_o,
  slice_o,
  bank_o,
  data_o
);

  input [39:0] paddr_i;
  input [127:0] data_i;
  output [32:0] daddr_o;
  output [0:0] slice_o;
  output [0:0] bank_o;
  output [127:0] data_o;
  output dram_o;
  wire [32:0] daddr_o,daddr;
  wire [0:0] slice_o,bank_o,tag_slice;
  wire [127:0] data_o;
  wire dram_o,N0,N1,is_csr_addr,is_tag_op,N2,is_addr_op,N3,N4,N5,N6,N7;
  assign data_o[127] = data_i[127];
  assign data_o[126] = data_i[126];
  assign data_o[125] = data_i[125];
  assign data_o[124] = data_i[124];
  assign data_o[123] = data_i[123];
  assign data_o[122] = data_i[122];
  assign data_o[121] = data_i[121];
  assign data_o[120] = data_i[120];
  assign data_o[119] = data_i[119];
  assign data_o[118] = data_i[118];
  assign data_o[117] = data_i[117];
  assign data_o[116] = data_i[116];
  assign data_o[115] = data_i[115];
  assign data_o[114] = data_i[114];
  assign data_o[113] = data_i[113];
  assign data_o[112] = data_i[112];
  assign data_o[111] = data_i[111];
  assign data_o[110] = data_i[110];
  assign data_o[109] = data_i[109];
  assign data_o[108] = data_i[108];
  assign data_o[107] = data_i[107];
  assign data_o[106] = data_i[106];
  assign data_o[105] = data_i[105];
  assign data_o[104] = data_i[104];
  assign data_o[103] = data_i[103];
  assign data_o[102] = data_i[102];
  assign data_o[101] = data_i[101];
  assign data_o[100] = data_i[100];
  assign data_o[99] = data_i[99];
  assign data_o[98] = data_i[98];
  assign data_o[97] = data_i[97];
  assign data_o[96] = data_i[96];
  assign data_o[95] = data_i[95];
  assign data_o[94] = data_i[94];
  assign data_o[93] = data_i[93];
  assign data_o[92] = data_i[92];
  assign data_o[91] = data_i[91];
  assign data_o[90] = data_i[90];
  assign data_o[89] = data_i[89];
  assign data_o[88] = data_i[88];
  assign data_o[87] = data_i[87];
  assign data_o[86] = data_i[86];
  assign data_o[85] = data_i[85];
  assign data_o[84] = data_i[84];
  assign data_o[83] = data_i[83];
  assign data_o[82] = data_i[82];
  assign data_o[81] = data_i[81];
  assign data_o[80] = data_i[80];
  assign data_o[79] = data_i[79];
  assign data_o[78] = data_i[78];
  assign data_o[77] = data_i[77];
  assign data_o[76] = data_i[76];
  assign data_o[75] = data_i[75];
  assign data_o[74] = data_i[74];
  assign data_o[73] = data_i[73];
  assign data_o[72] = data_i[72];
  assign data_o[71] = data_i[71];
  assign data_o[70] = data_i[70];
  assign data_o[69] = data_i[69];
  assign data_o[68] = data_i[68];
  assign data_o[67] = data_i[67];
  assign data_o[66] = data_i[66];
  assign data_o[65] = data_i[65];
  assign data_o[64] = data_i[64];
  assign data_o[63] = data_i[63];
  assign data_o[62] = data_i[62];
  assign data_o[61] = data_i[61];
  assign data_o[60] = data_i[60];
  assign data_o[59] = data_i[59];
  assign data_o[58] = data_i[58];
  assign data_o[57] = data_i[57];
  assign data_o[56] = data_i[56];
  assign data_o[55] = data_i[55];
  assign data_o[54] = data_i[54];
  assign data_o[53] = data_i[53];
  assign data_o[52] = data_i[52];
  assign data_o[51] = data_i[51];
  assign data_o[50] = data_i[50];
  assign data_o[49] = data_i[49];
  assign data_o[48] = data_i[48];
  assign data_o[47] = data_i[47];
  assign data_o[46] = data_i[46];
  assign data_o[45] = data_i[45];
  assign data_o[44] = data_i[44];
  assign data_o[43] = data_i[43];
  assign data_o[42] = data_i[42];
  assign data_o[41] = data_i[41];
  assign data_o[40] = data_i[40];
  assign data_o[39] = data_i[39];
  assign data_o[38] = data_i[38];
  assign data_o[37] = data_i[37];
  assign data_o[36] = data_i[36];
  assign data_o[35] = data_i[35];
  assign data_o[34] = data_i[34];
  assign data_o[33] = data_i[33];
  assign data_o[32] = data_i[32];
  assign data_o[31] = data_i[31];
  assign data_o[30] = data_i[30];
  assign data_o[29] = data_i[29];
  assign data_o[28] = data_i[28];
  assign data_o[27] = data_i[27];
  assign data_o[26] = data_i[26];
  assign data_o[25] = data_i[25];
  assign data_o[24] = data_i[24];
  assign data_o[23] = data_i[23];
  assign data_o[22] = data_i[22];
  assign data_o[21] = data_i[21];
  assign data_o[20] = data_i[20];
  assign data_o[19] = data_i[19];
  assign data_o[18] = data_i[18];
  assign data_o[17] = data_i[17];
  assign data_o[16] = data_i[16];
  assign data_o[15] = data_i[15];
  assign data_o[14] = data_i[14];
  assign data_o[13] = data_i[13];
  assign data_o[12] = data_i[12];
  assign data_o[11] = data_i[11];
  assign data_o[10] = data_i[10];
  assign data_o[9] = data_i[9];
  assign data_o[8] = data_i[8];
  assign data_o[7] = data_i[7];
  assign data_o[6] = data_i[6];
  assign data_o[5] = data_i[5];
  assign data_o[4] = data_i[4];
  assign data_o[3] = data_i[3];
  assign data_o[2] = data_i[2];
  assign data_o[1] = data_i[1];
  assign data_o[0] = data_i[0];
  assign dram_o = paddr_i >= { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign is_csr_addr = paddr_i < { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign N2 = ~paddr_i[5];
  assign tag_slice[0] = paddr_i[20] ^ 1'b0;
  assign daddr = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, paddr_i[16:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                 (N6)? data_o[32:0] : 
                 (N4)? paddr_i[32:0] : 1'b0;
  assign N0 = is_tag_op;
  assign daddr_o = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, paddr_i[16:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                   (N1)? daddr : 1'b0;
  assign N1 = N7;
  assign slice_o[0] = (N0)? tag_slice[0] : 
                      (N1)? daddr[6] : 1'b0;
  assign bank_o[0] = (N0)? paddr_i[17] : 
                     (N1)? daddr[7] : 1'b0;
  assign is_tag_op = is_csr_addr & paddr_i[5];
  assign is_addr_op = is_csr_addr & N2;
  assign N3 = is_addr_op | is_tag_op;
  assign N4 = ~N3;
  assign N5 = ~is_tag_op;
  assign N6 = is_addr_op & N5;
  assign N7 = ~is_tag_op;

endmodule



module bsg_decode_00000002
(
  i,
  o
);

  input [0:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o = { 1'b0, 1'b1 } << i[0];

endmodule



module bsg_decode_with_v_00000002
(
  i,
  v_i,
  o
);

  input [0:0] i;
  output [1:0] o;
  input v_i;
  wire [1:0] o,lo;

  bsg_decode_00000002
  bd
  (
    .i(i[0]),
    .o(lo)
  );

  assign o[1] = v_i & lo[1];
  assign o[0] = v_i & lo[0];

endmodule



module bsg_mux_00000080_00000002
(
  data_i,
  sel_i,
  data_o
);

  input [255:0] data_i;
  input [0:0] sel_i;
  output [127:0] data_o;
  wire [127:0] data_o;
  wire N0,N1;
  assign data_o[127] = (N1)? data_i[127] : 
                       (N0)? data_i[255] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[126] = (N1)? data_i[126] : 
                       (N0)? data_i[254] : 1'b0;
  assign data_o[125] = (N1)? data_i[125] : 
                       (N0)? data_i[253] : 1'b0;
  assign data_o[124] = (N1)? data_i[124] : 
                       (N0)? data_i[252] : 1'b0;
  assign data_o[123] = (N1)? data_i[123] : 
                       (N0)? data_i[251] : 1'b0;
  assign data_o[122] = (N1)? data_i[122] : 
                       (N0)? data_i[250] : 1'b0;
  assign data_o[121] = (N1)? data_i[121] : 
                       (N0)? data_i[249] : 1'b0;
  assign data_o[120] = (N1)? data_i[120] : 
                       (N0)? data_i[248] : 1'b0;
  assign data_o[119] = (N1)? data_i[119] : 
                       (N0)? data_i[247] : 1'b0;
  assign data_o[118] = (N1)? data_i[118] : 
                       (N0)? data_i[246] : 1'b0;
  assign data_o[117] = (N1)? data_i[117] : 
                       (N0)? data_i[245] : 1'b0;
  assign data_o[116] = (N1)? data_i[116] : 
                       (N0)? data_i[244] : 1'b0;
  assign data_o[115] = (N1)? data_i[115] : 
                       (N0)? data_i[243] : 1'b0;
  assign data_o[114] = (N1)? data_i[114] : 
                       (N0)? data_i[242] : 1'b0;
  assign data_o[113] = (N1)? data_i[113] : 
                       (N0)? data_i[241] : 1'b0;
  assign data_o[112] = (N1)? data_i[112] : 
                       (N0)? data_i[240] : 1'b0;
  assign data_o[111] = (N1)? data_i[111] : 
                       (N0)? data_i[239] : 1'b0;
  assign data_o[110] = (N1)? data_i[110] : 
                       (N0)? data_i[238] : 1'b0;
  assign data_o[109] = (N1)? data_i[109] : 
                       (N0)? data_i[237] : 1'b0;
  assign data_o[108] = (N1)? data_i[108] : 
                       (N0)? data_i[236] : 1'b0;
  assign data_o[107] = (N1)? data_i[107] : 
                       (N0)? data_i[235] : 1'b0;
  assign data_o[106] = (N1)? data_i[106] : 
                       (N0)? data_i[234] : 1'b0;
  assign data_o[105] = (N1)? data_i[105] : 
                       (N0)? data_i[233] : 1'b0;
  assign data_o[104] = (N1)? data_i[104] : 
                       (N0)? data_i[232] : 1'b0;
  assign data_o[103] = (N1)? data_i[103] : 
                       (N0)? data_i[231] : 1'b0;
  assign data_o[102] = (N1)? data_i[102] : 
                       (N0)? data_i[230] : 1'b0;
  assign data_o[101] = (N1)? data_i[101] : 
                       (N0)? data_i[229] : 1'b0;
  assign data_o[100] = (N1)? data_i[100] : 
                       (N0)? data_i[228] : 1'b0;
  assign data_o[99] = (N1)? data_i[99] : 
                      (N0)? data_i[227] : 1'b0;
  assign data_o[98] = (N1)? data_i[98] : 
                      (N0)? data_i[226] : 1'b0;
  assign data_o[97] = (N1)? data_i[97] : 
                      (N0)? data_i[225] : 1'b0;
  assign data_o[96] = (N1)? data_i[96] : 
                      (N0)? data_i[224] : 1'b0;
  assign data_o[95] = (N1)? data_i[95] : 
                      (N0)? data_i[223] : 1'b0;
  assign data_o[94] = (N1)? data_i[94] : 
                      (N0)? data_i[222] : 1'b0;
  assign data_o[93] = (N1)? data_i[93] : 
                      (N0)? data_i[221] : 1'b0;
  assign data_o[92] = (N1)? data_i[92] : 
                      (N0)? data_i[220] : 1'b0;
  assign data_o[91] = (N1)? data_i[91] : 
                      (N0)? data_i[219] : 1'b0;
  assign data_o[90] = (N1)? data_i[90] : 
                      (N0)? data_i[218] : 1'b0;
  assign data_o[89] = (N1)? data_i[89] : 
                      (N0)? data_i[217] : 1'b0;
  assign data_o[88] = (N1)? data_i[88] : 
                      (N0)? data_i[216] : 1'b0;
  assign data_o[87] = (N1)? data_i[87] : 
                      (N0)? data_i[215] : 1'b0;
  assign data_o[86] = (N1)? data_i[86] : 
                      (N0)? data_i[214] : 1'b0;
  assign data_o[85] = (N1)? data_i[85] : 
                      (N0)? data_i[213] : 1'b0;
  assign data_o[84] = (N1)? data_i[84] : 
                      (N0)? data_i[212] : 1'b0;
  assign data_o[83] = (N1)? data_i[83] : 
                      (N0)? data_i[211] : 1'b0;
  assign data_o[82] = (N1)? data_i[82] : 
                      (N0)? data_i[210] : 1'b0;
  assign data_o[81] = (N1)? data_i[81] : 
                      (N0)? data_i[209] : 1'b0;
  assign data_o[80] = (N1)? data_i[80] : 
                      (N0)? data_i[208] : 1'b0;
  assign data_o[79] = (N1)? data_i[79] : 
                      (N0)? data_i[207] : 1'b0;
  assign data_o[78] = (N1)? data_i[78] : 
                      (N0)? data_i[206] : 1'b0;
  assign data_o[77] = (N1)? data_i[77] : 
                      (N0)? data_i[205] : 1'b0;
  assign data_o[76] = (N1)? data_i[76] : 
                      (N0)? data_i[204] : 1'b0;
  assign data_o[75] = (N1)? data_i[75] : 
                      (N0)? data_i[203] : 1'b0;
  assign data_o[74] = (N1)? data_i[74] : 
                      (N0)? data_i[202] : 1'b0;
  assign data_o[73] = (N1)? data_i[73] : 
                      (N0)? data_i[201] : 1'b0;
  assign data_o[72] = (N1)? data_i[72] : 
                      (N0)? data_i[200] : 1'b0;
  assign data_o[71] = (N1)? data_i[71] : 
                      (N0)? data_i[199] : 1'b0;
  assign data_o[70] = (N1)? data_i[70] : 
                      (N0)? data_i[198] : 1'b0;
  assign data_o[69] = (N1)? data_i[69] : 
                      (N0)? data_i[197] : 1'b0;
  assign data_o[68] = (N1)? data_i[68] : 
                      (N0)? data_i[196] : 1'b0;
  assign data_o[67] = (N1)? data_i[67] : 
                      (N0)? data_i[195] : 1'b0;
  assign data_o[66] = (N1)? data_i[66] : 
                      (N0)? data_i[194] : 1'b0;
  assign data_o[65] = (N1)? data_i[65] : 
                      (N0)? data_i[193] : 1'b0;
  assign data_o[64] = (N1)? data_i[64] : 
                      (N0)? data_i[192] : 1'b0;
  assign data_o[63] = (N1)? data_i[63] : 
                      (N0)? data_i[191] : 1'b0;
  assign data_o[62] = (N1)? data_i[62] : 
                      (N0)? data_i[190] : 1'b0;
  assign data_o[61] = (N1)? data_i[61] : 
                      (N0)? data_i[189] : 1'b0;
  assign data_o[60] = (N1)? data_i[60] : 
                      (N0)? data_i[188] : 1'b0;
  assign data_o[59] = (N1)? data_i[59] : 
                      (N0)? data_i[187] : 1'b0;
  assign data_o[58] = (N1)? data_i[58] : 
                      (N0)? data_i[186] : 1'b0;
  assign data_o[57] = (N1)? data_i[57] : 
                      (N0)? data_i[185] : 1'b0;
  assign data_o[56] = (N1)? data_i[56] : 
                      (N0)? data_i[184] : 1'b0;
  assign data_o[55] = (N1)? data_i[55] : 
                      (N0)? data_i[183] : 1'b0;
  assign data_o[54] = (N1)? data_i[54] : 
                      (N0)? data_i[182] : 1'b0;
  assign data_o[53] = (N1)? data_i[53] : 
                      (N0)? data_i[181] : 1'b0;
  assign data_o[52] = (N1)? data_i[52] : 
                      (N0)? data_i[180] : 1'b0;
  assign data_o[51] = (N1)? data_i[51] : 
                      (N0)? data_i[179] : 1'b0;
  assign data_o[50] = (N1)? data_i[50] : 
                      (N0)? data_i[178] : 1'b0;
  assign data_o[49] = (N1)? data_i[49] : 
                      (N0)? data_i[177] : 1'b0;
  assign data_o[48] = (N1)? data_i[48] : 
                      (N0)? data_i[176] : 1'b0;
  assign data_o[47] = (N1)? data_i[47] : 
                      (N0)? data_i[175] : 1'b0;
  assign data_o[46] = (N1)? data_i[46] : 
                      (N0)? data_i[174] : 1'b0;
  assign data_o[45] = (N1)? data_i[45] : 
                      (N0)? data_i[173] : 1'b0;
  assign data_o[44] = (N1)? data_i[44] : 
                      (N0)? data_i[172] : 1'b0;
  assign data_o[43] = (N1)? data_i[43] : 
                      (N0)? data_i[171] : 1'b0;
  assign data_o[42] = (N1)? data_i[42] : 
                      (N0)? data_i[170] : 1'b0;
  assign data_o[41] = (N1)? data_i[41] : 
                      (N0)? data_i[169] : 1'b0;
  assign data_o[40] = (N1)? data_i[40] : 
                      (N0)? data_i[168] : 1'b0;
  assign data_o[39] = (N1)? data_i[39] : 
                      (N0)? data_i[167] : 1'b0;
  assign data_o[38] = (N1)? data_i[38] : 
                      (N0)? data_i[166] : 1'b0;
  assign data_o[37] = (N1)? data_i[37] : 
                      (N0)? data_i[165] : 1'b0;
  assign data_o[36] = (N1)? data_i[36] : 
                      (N0)? data_i[164] : 1'b0;
  assign data_o[35] = (N1)? data_i[35] : 
                      (N0)? data_i[163] : 1'b0;
  assign data_o[34] = (N1)? data_i[34] : 
                      (N0)? data_i[162] : 1'b0;
  assign data_o[33] = (N1)? data_i[33] : 
                      (N0)? data_i[161] : 1'b0;
  assign data_o[32] = (N1)? data_i[32] : 
                      (N0)? data_i[160] : 1'b0;
  assign data_o[31] = (N1)? data_i[31] : 
                      (N0)? data_i[159] : 1'b0;
  assign data_o[30] = (N1)? data_i[30] : 
                      (N0)? data_i[158] : 1'b0;
  assign data_o[29] = (N1)? data_i[29] : 
                      (N0)? data_i[157] : 1'b0;
  assign data_o[28] = (N1)? data_i[28] : 
                      (N0)? data_i[156] : 1'b0;
  assign data_o[27] = (N1)? data_i[27] : 
                      (N0)? data_i[155] : 1'b0;
  assign data_o[26] = (N1)? data_i[26] : 
                      (N0)? data_i[154] : 1'b0;
  assign data_o[25] = (N1)? data_i[25] : 
                      (N0)? data_i[153] : 1'b0;
  assign data_o[24] = (N1)? data_i[24] : 
                      (N0)? data_i[152] : 1'b0;
  assign data_o[23] = (N1)? data_i[23] : 
                      (N0)? data_i[151] : 1'b0;
  assign data_o[22] = (N1)? data_i[22] : 
                      (N0)? data_i[150] : 1'b0;
  assign data_o[21] = (N1)? data_i[21] : 
                      (N0)? data_i[149] : 1'b0;
  assign data_o[20] = (N1)? data_i[20] : 
                      (N0)? data_i[148] : 1'b0;
  assign data_o[19] = (N1)? data_i[19] : 
                      (N0)? data_i[147] : 1'b0;
  assign data_o[18] = (N1)? data_i[18] : 
                      (N0)? data_i[146] : 1'b0;
  assign data_o[17] = (N1)? data_i[17] : 
                      (N0)? data_i[145] : 1'b0;
  assign data_o[16] = (N1)? data_i[16] : 
                      (N0)? data_i[144] : 1'b0;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[143] : 1'b0;
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[142] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[141] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[140] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[139] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[138] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[137] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[136] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[135] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[134] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[133] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[132] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[131] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[130] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[129] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[128] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_rotate_right_00000080
(
  data_i,
  rot_i,
  o
);

  input [127:0] data_i;
  input [6:0] rot_i;
  output [127:0] o;
  wire [127:0] o;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,
  sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,
  sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,sv2v_dc_21,sv2v_dc_22,
  sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,sv2v_dc_27,sv2v_dc_28,sv2v_dc_29,
  sv2v_dc_30,sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,sv2v_dc_34,sv2v_dc_35,sv2v_dc_36,sv2v_dc_37,
  sv2v_dc_38,sv2v_dc_39,sv2v_dc_40,sv2v_dc_41,sv2v_dc_42,sv2v_dc_43,sv2v_dc_44,
  sv2v_dc_45,sv2v_dc_46,sv2v_dc_47,sv2v_dc_48,sv2v_dc_49,sv2v_dc_50,sv2v_dc_51,
  sv2v_dc_52,sv2v_dc_53,sv2v_dc_54,sv2v_dc_55,sv2v_dc_56,sv2v_dc_57,sv2v_dc_58,sv2v_dc_59,
  sv2v_dc_60,sv2v_dc_61,sv2v_dc_62,sv2v_dc_63,sv2v_dc_64,sv2v_dc_65,sv2v_dc_66,
  sv2v_dc_67,sv2v_dc_68,sv2v_dc_69,sv2v_dc_70,sv2v_dc_71,sv2v_dc_72,sv2v_dc_73,
  sv2v_dc_74,sv2v_dc_75,sv2v_dc_76,sv2v_dc_77,sv2v_dc_78,sv2v_dc_79,sv2v_dc_80,
  sv2v_dc_81,sv2v_dc_82,sv2v_dc_83,sv2v_dc_84,sv2v_dc_85,sv2v_dc_86,sv2v_dc_87,sv2v_dc_88,
  sv2v_dc_89,sv2v_dc_90,sv2v_dc_91,sv2v_dc_92,sv2v_dc_93,sv2v_dc_94,sv2v_dc_95,
  sv2v_dc_96,sv2v_dc_97,sv2v_dc_98,sv2v_dc_99,sv2v_dc_100,sv2v_dc_101,sv2v_dc_102,
  sv2v_dc_103,sv2v_dc_104,sv2v_dc_105,sv2v_dc_106,sv2v_dc_107,sv2v_dc_108,sv2v_dc_109,
  sv2v_dc_110,sv2v_dc_111,sv2v_dc_112,sv2v_dc_113,sv2v_dc_114,sv2v_dc_115,
  sv2v_dc_116,sv2v_dc_117,sv2v_dc_118,sv2v_dc_119,sv2v_dc_120,sv2v_dc_121,sv2v_dc_122,
  sv2v_dc_123,sv2v_dc_124,sv2v_dc_125,sv2v_dc_126,sv2v_dc_127;
  assign { sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36, sv2v_dc_37, sv2v_dc_38, sv2v_dc_39, sv2v_dc_40, sv2v_dc_41, sv2v_dc_42, sv2v_dc_43, sv2v_dc_44, sv2v_dc_45, sv2v_dc_46, sv2v_dc_47, sv2v_dc_48, sv2v_dc_49, sv2v_dc_50, sv2v_dc_51, sv2v_dc_52, sv2v_dc_53, sv2v_dc_54, sv2v_dc_55, sv2v_dc_56, sv2v_dc_57, sv2v_dc_58, sv2v_dc_59, sv2v_dc_60, sv2v_dc_61, sv2v_dc_62, sv2v_dc_63, sv2v_dc_64, sv2v_dc_65, sv2v_dc_66, sv2v_dc_67, sv2v_dc_68, sv2v_dc_69, sv2v_dc_70, sv2v_dc_71, sv2v_dc_72, sv2v_dc_73, sv2v_dc_74, sv2v_dc_75, sv2v_dc_76, sv2v_dc_77, sv2v_dc_78, sv2v_dc_79, sv2v_dc_80, sv2v_dc_81, sv2v_dc_82, sv2v_dc_83, sv2v_dc_84, sv2v_dc_85, sv2v_dc_86, sv2v_dc_87, sv2v_dc_88, sv2v_dc_89, sv2v_dc_90, sv2v_dc_91, sv2v_dc_92, sv2v_dc_93, sv2v_dc_94, sv2v_dc_95, sv2v_dc_96, sv2v_dc_97, sv2v_dc_98, sv2v_dc_99, sv2v_dc_100, sv2v_dc_101, sv2v_dc_102, sv2v_dc_103, sv2v_dc_104, sv2v_dc_105, sv2v_dc_106, sv2v_dc_107, sv2v_dc_108, sv2v_dc_109, sv2v_dc_110, sv2v_dc_111, sv2v_dc_112, sv2v_dc_113, sv2v_dc_114, sv2v_dc_115, sv2v_dc_116, sv2v_dc_117, sv2v_dc_118, sv2v_dc_119, sv2v_dc_120, sv2v_dc_121, sv2v_dc_122, sv2v_dc_123, sv2v_dc_124, sv2v_dc_125, sv2v_dc_126, sv2v_dc_127, o } = { data_i[126:0], data_i } >> rot_i;

endmodule



module bsg_mux_00000080_00000008
(
  data_i,
  sel_i,
  data_o
);

  input [1023:0] data_i;
  input [2:0] sel_i;
  output [127:0] data_o;
  wire [127:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;
  assign data_o[127] = (N7)? data_i[127] : 
                       (N9)? data_i[255] : 
                       (N11)? data_i[383] : 
                       (N13)? data_i[511] : 
                       (N8)? data_i[639] : 
                       (N10)? data_i[767] : 
                       (N12)? data_i[895] : 
                       (N14)? data_i[1023] : 1'b0;
  assign data_o[126] = (N7)? data_i[126] : 
                       (N9)? data_i[254] : 
                       (N11)? data_i[382] : 
                       (N13)? data_i[510] : 
                       (N8)? data_i[638] : 
                       (N10)? data_i[766] : 
                       (N12)? data_i[894] : 
                       (N14)? data_i[1022] : 1'b0;
  assign data_o[125] = (N7)? data_i[125] : 
                       (N9)? data_i[253] : 
                       (N11)? data_i[381] : 
                       (N13)? data_i[509] : 
                       (N8)? data_i[637] : 
                       (N10)? data_i[765] : 
                       (N12)? data_i[893] : 
                       (N14)? data_i[1021] : 1'b0;
  assign data_o[124] = (N7)? data_i[124] : 
                       (N9)? data_i[252] : 
                       (N11)? data_i[380] : 
                       (N13)? data_i[508] : 
                       (N8)? data_i[636] : 
                       (N10)? data_i[764] : 
                       (N12)? data_i[892] : 
                       (N14)? data_i[1020] : 1'b0;
  assign data_o[123] = (N7)? data_i[123] : 
                       (N9)? data_i[251] : 
                       (N11)? data_i[379] : 
                       (N13)? data_i[507] : 
                       (N8)? data_i[635] : 
                       (N10)? data_i[763] : 
                       (N12)? data_i[891] : 
                       (N14)? data_i[1019] : 1'b0;
  assign data_o[122] = (N7)? data_i[122] : 
                       (N9)? data_i[250] : 
                       (N11)? data_i[378] : 
                       (N13)? data_i[506] : 
                       (N8)? data_i[634] : 
                       (N10)? data_i[762] : 
                       (N12)? data_i[890] : 
                       (N14)? data_i[1018] : 1'b0;
  assign data_o[121] = (N7)? data_i[121] : 
                       (N9)? data_i[249] : 
                       (N11)? data_i[377] : 
                       (N13)? data_i[505] : 
                       (N8)? data_i[633] : 
                       (N10)? data_i[761] : 
                       (N12)? data_i[889] : 
                       (N14)? data_i[1017] : 1'b0;
  assign data_o[120] = (N7)? data_i[120] : 
                       (N9)? data_i[248] : 
                       (N11)? data_i[376] : 
                       (N13)? data_i[504] : 
                       (N8)? data_i[632] : 
                       (N10)? data_i[760] : 
                       (N12)? data_i[888] : 
                       (N14)? data_i[1016] : 1'b0;
  assign data_o[119] = (N7)? data_i[119] : 
                       (N9)? data_i[247] : 
                       (N11)? data_i[375] : 
                       (N13)? data_i[503] : 
                       (N8)? data_i[631] : 
                       (N10)? data_i[759] : 
                       (N12)? data_i[887] : 
                       (N14)? data_i[1015] : 1'b0;
  assign data_o[118] = (N7)? data_i[118] : 
                       (N9)? data_i[246] : 
                       (N11)? data_i[374] : 
                       (N13)? data_i[502] : 
                       (N8)? data_i[630] : 
                       (N10)? data_i[758] : 
                       (N12)? data_i[886] : 
                       (N14)? data_i[1014] : 1'b0;
  assign data_o[117] = (N7)? data_i[117] : 
                       (N9)? data_i[245] : 
                       (N11)? data_i[373] : 
                       (N13)? data_i[501] : 
                       (N8)? data_i[629] : 
                       (N10)? data_i[757] : 
                       (N12)? data_i[885] : 
                       (N14)? data_i[1013] : 1'b0;
  assign data_o[116] = (N7)? data_i[116] : 
                       (N9)? data_i[244] : 
                       (N11)? data_i[372] : 
                       (N13)? data_i[500] : 
                       (N8)? data_i[628] : 
                       (N10)? data_i[756] : 
                       (N12)? data_i[884] : 
                       (N14)? data_i[1012] : 1'b0;
  assign data_o[115] = (N7)? data_i[115] : 
                       (N9)? data_i[243] : 
                       (N11)? data_i[371] : 
                       (N13)? data_i[499] : 
                       (N8)? data_i[627] : 
                       (N10)? data_i[755] : 
                       (N12)? data_i[883] : 
                       (N14)? data_i[1011] : 1'b0;
  assign data_o[114] = (N7)? data_i[114] : 
                       (N9)? data_i[242] : 
                       (N11)? data_i[370] : 
                       (N13)? data_i[498] : 
                       (N8)? data_i[626] : 
                       (N10)? data_i[754] : 
                       (N12)? data_i[882] : 
                       (N14)? data_i[1010] : 1'b0;
  assign data_o[113] = (N7)? data_i[113] : 
                       (N9)? data_i[241] : 
                       (N11)? data_i[369] : 
                       (N13)? data_i[497] : 
                       (N8)? data_i[625] : 
                       (N10)? data_i[753] : 
                       (N12)? data_i[881] : 
                       (N14)? data_i[1009] : 1'b0;
  assign data_o[112] = (N7)? data_i[112] : 
                       (N9)? data_i[240] : 
                       (N11)? data_i[368] : 
                       (N13)? data_i[496] : 
                       (N8)? data_i[624] : 
                       (N10)? data_i[752] : 
                       (N12)? data_i[880] : 
                       (N14)? data_i[1008] : 1'b0;
  assign data_o[111] = (N7)? data_i[111] : 
                       (N9)? data_i[239] : 
                       (N11)? data_i[367] : 
                       (N13)? data_i[495] : 
                       (N8)? data_i[623] : 
                       (N10)? data_i[751] : 
                       (N12)? data_i[879] : 
                       (N14)? data_i[1007] : 1'b0;
  assign data_o[110] = (N7)? data_i[110] : 
                       (N9)? data_i[238] : 
                       (N11)? data_i[366] : 
                       (N13)? data_i[494] : 
                       (N8)? data_i[622] : 
                       (N10)? data_i[750] : 
                       (N12)? data_i[878] : 
                       (N14)? data_i[1006] : 1'b0;
  assign data_o[109] = (N7)? data_i[109] : 
                       (N9)? data_i[237] : 
                       (N11)? data_i[365] : 
                       (N13)? data_i[493] : 
                       (N8)? data_i[621] : 
                       (N10)? data_i[749] : 
                       (N12)? data_i[877] : 
                       (N14)? data_i[1005] : 1'b0;
  assign data_o[108] = (N7)? data_i[108] : 
                       (N9)? data_i[236] : 
                       (N11)? data_i[364] : 
                       (N13)? data_i[492] : 
                       (N8)? data_i[620] : 
                       (N10)? data_i[748] : 
                       (N12)? data_i[876] : 
                       (N14)? data_i[1004] : 1'b0;
  assign data_o[107] = (N7)? data_i[107] : 
                       (N9)? data_i[235] : 
                       (N11)? data_i[363] : 
                       (N13)? data_i[491] : 
                       (N8)? data_i[619] : 
                       (N10)? data_i[747] : 
                       (N12)? data_i[875] : 
                       (N14)? data_i[1003] : 1'b0;
  assign data_o[106] = (N7)? data_i[106] : 
                       (N9)? data_i[234] : 
                       (N11)? data_i[362] : 
                       (N13)? data_i[490] : 
                       (N8)? data_i[618] : 
                       (N10)? data_i[746] : 
                       (N12)? data_i[874] : 
                       (N14)? data_i[1002] : 1'b0;
  assign data_o[105] = (N7)? data_i[105] : 
                       (N9)? data_i[233] : 
                       (N11)? data_i[361] : 
                       (N13)? data_i[489] : 
                       (N8)? data_i[617] : 
                       (N10)? data_i[745] : 
                       (N12)? data_i[873] : 
                       (N14)? data_i[1001] : 1'b0;
  assign data_o[104] = (N7)? data_i[104] : 
                       (N9)? data_i[232] : 
                       (N11)? data_i[360] : 
                       (N13)? data_i[488] : 
                       (N8)? data_i[616] : 
                       (N10)? data_i[744] : 
                       (N12)? data_i[872] : 
                       (N14)? data_i[1000] : 1'b0;
  assign data_o[103] = (N7)? data_i[103] : 
                       (N9)? data_i[231] : 
                       (N11)? data_i[359] : 
                       (N13)? data_i[487] : 
                       (N8)? data_i[615] : 
                       (N10)? data_i[743] : 
                       (N12)? data_i[871] : 
                       (N14)? data_i[999] : 1'b0;
  assign data_o[102] = (N7)? data_i[102] : 
                       (N9)? data_i[230] : 
                       (N11)? data_i[358] : 
                       (N13)? data_i[486] : 
                       (N8)? data_i[614] : 
                       (N10)? data_i[742] : 
                       (N12)? data_i[870] : 
                       (N14)? data_i[998] : 1'b0;
  assign data_o[101] = (N7)? data_i[101] : 
                       (N9)? data_i[229] : 
                       (N11)? data_i[357] : 
                       (N13)? data_i[485] : 
                       (N8)? data_i[613] : 
                       (N10)? data_i[741] : 
                       (N12)? data_i[869] : 
                       (N14)? data_i[997] : 1'b0;
  assign data_o[100] = (N7)? data_i[100] : 
                       (N9)? data_i[228] : 
                       (N11)? data_i[356] : 
                       (N13)? data_i[484] : 
                       (N8)? data_i[612] : 
                       (N10)? data_i[740] : 
                       (N12)? data_i[868] : 
                       (N14)? data_i[996] : 1'b0;
  assign data_o[99] = (N7)? data_i[99] : 
                      (N9)? data_i[227] : 
                      (N11)? data_i[355] : 
                      (N13)? data_i[483] : 
                      (N8)? data_i[611] : 
                      (N10)? data_i[739] : 
                      (N12)? data_i[867] : 
                      (N14)? data_i[995] : 1'b0;
  assign data_o[98] = (N7)? data_i[98] : 
                      (N9)? data_i[226] : 
                      (N11)? data_i[354] : 
                      (N13)? data_i[482] : 
                      (N8)? data_i[610] : 
                      (N10)? data_i[738] : 
                      (N12)? data_i[866] : 
                      (N14)? data_i[994] : 1'b0;
  assign data_o[97] = (N7)? data_i[97] : 
                      (N9)? data_i[225] : 
                      (N11)? data_i[353] : 
                      (N13)? data_i[481] : 
                      (N8)? data_i[609] : 
                      (N10)? data_i[737] : 
                      (N12)? data_i[865] : 
                      (N14)? data_i[993] : 1'b0;
  assign data_o[96] = (N7)? data_i[96] : 
                      (N9)? data_i[224] : 
                      (N11)? data_i[352] : 
                      (N13)? data_i[480] : 
                      (N8)? data_i[608] : 
                      (N10)? data_i[736] : 
                      (N12)? data_i[864] : 
                      (N14)? data_i[992] : 1'b0;
  assign data_o[95] = (N7)? data_i[95] : 
                      (N9)? data_i[223] : 
                      (N11)? data_i[351] : 
                      (N13)? data_i[479] : 
                      (N8)? data_i[607] : 
                      (N10)? data_i[735] : 
                      (N12)? data_i[863] : 
                      (N14)? data_i[991] : 1'b0;
  assign data_o[94] = (N7)? data_i[94] : 
                      (N9)? data_i[222] : 
                      (N11)? data_i[350] : 
                      (N13)? data_i[478] : 
                      (N8)? data_i[606] : 
                      (N10)? data_i[734] : 
                      (N12)? data_i[862] : 
                      (N14)? data_i[990] : 1'b0;
  assign data_o[93] = (N7)? data_i[93] : 
                      (N9)? data_i[221] : 
                      (N11)? data_i[349] : 
                      (N13)? data_i[477] : 
                      (N8)? data_i[605] : 
                      (N10)? data_i[733] : 
                      (N12)? data_i[861] : 
                      (N14)? data_i[989] : 1'b0;
  assign data_o[92] = (N7)? data_i[92] : 
                      (N9)? data_i[220] : 
                      (N11)? data_i[348] : 
                      (N13)? data_i[476] : 
                      (N8)? data_i[604] : 
                      (N10)? data_i[732] : 
                      (N12)? data_i[860] : 
                      (N14)? data_i[988] : 1'b0;
  assign data_o[91] = (N7)? data_i[91] : 
                      (N9)? data_i[219] : 
                      (N11)? data_i[347] : 
                      (N13)? data_i[475] : 
                      (N8)? data_i[603] : 
                      (N10)? data_i[731] : 
                      (N12)? data_i[859] : 
                      (N14)? data_i[987] : 1'b0;
  assign data_o[90] = (N7)? data_i[90] : 
                      (N9)? data_i[218] : 
                      (N11)? data_i[346] : 
                      (N13)? data_i[474] : 
                      (N8)? data_i[602] : 
                      (N10)? data_i[730] : 
                      (N12)? data_i[858] : 
                      (N14)? data_i[986] : 1'b0;
  assign data_o[89] = (N7)? data_i[89] : 
                      (N9)? data_i[217] : 
                      (N11)? data_i[345] : 
                      (N13)? data_i[473] : 
                      (N8)? data_i[601] : 
                      (N10)? data_i[729] : 
                      (N12)? data_i[857] : 
                      (N14)? data_i[985] : 1'b0;
  assign data_o[88] = (N7)? data_i[88] : 
                      (N9)? data_i[216] : 
                      (N11)? data_i[344] : 
                      (N13)? data_i[472] : 
                      (N8)? data_i[600] : 
                      (N10)? data_i[728] : 
                      (N12)? data_i[856] : 
                      (N14)? data_i[984] : 1'b0;
  assign data_o[87] = (N7)? data_i[87] : 
                      (N9)? data_i[215] : 
                      (N11)? data_i[343] : 
                      (N13)? data_i[471] : 
                      (N8)? data_i[599] : 
                      (N10)? data_i[727] : 
                      (N12)? data_i[855] : 
                      (N14)? data_i[983] : 1'b0;
  assign data_o[86] = (N7)? data_i[86] : 
                      (N9)? data_i[214] : 
                      (N11)? data_i[342] : 
                      (N13)? data_i[470] : 
                      (N8)? data_i[598] : 
                      (N10)? data_i[726] : 
                      (N12)? data_i[854] : 
                      (N14)? data_i[982] : 1'b0;
  assign data_o[85] = (N7)? data_i[85] : 
                      (N9)? data_i[213] : 
                      (N11)? data_i[341] : 
                      (N13)? data_i[469] : 
                      (N8)? data_i[597] : 
                      (N10)? data_i[725] : 
                      (N12)? data_i[853] : 
                      (N14)? data_i[981] : 1'b0;
  assign data_o[84] = (N7)? data_i[84] : 
                      (N9)? data_i[212] : 
                      (N11)? data_i[340] : 
                      (N13)? data_i[468] : 
                      (N8)? data_i[596] : 
                      (N10)? data_i[724] : 
                      (N12)? data_i[852] : 
                      (N14)? data_i[980] : 1'b0;
  assign data_o[83] = (N7)? data_i[83] : 
                      (N9)? data_i[211] : 
                      (N11)? data_i[339] : 
                      (N13)? data_i[467] : 
                      (N8)? data_i[595] : 
                      (N10)? data_i[723] : 
                      (N12)? data_i[851] : 
                      (N14)? data_i[979] : 1'b0;
  assign data_o[82] = (N7)? data_i[82] : 
                      (N9)? data_i[210] : 
                      (N11)? data_i[338] : 
                      (N13)? data_i[466] : 
                      (N8)? data_i[594] : 
                      (N10)? data_i[722] : 
                      (N12)? data_i[850] : 
                      (N14)? data_i[978] : 1'b0;
  assign data_o[81] = (N7)? data_i[81] : 
                      (N9)? data_i[209] : 
                      (N11)? data_i[337] : 
                      (N13)? data_i[465] : 
                      (N8)? data_i[593] : 
                      (N10)? data_i[721] : 
                      (N12)? data_i[849] : 
                      (N14)? data_i[977] : 1'b0;
  assign data_o[80] = (N7)? data_i[80] : 
                      (N9)? data_i[208] : 
                      (N11)? data_i[336] : 
                      (N13)? data_i[464] : 
                      (N8)? data_i[592] : 
                      (N10)? data_i[720] : 
                      (N12)? data_i[848] : 
                      (N14)? data_i[976] : 1'b0;
  assign data_o[79] = (N7)? data_i[79] : 
                      (N9)? data_i[207] : 
                      (N11)? data_i[335] : 
                      (N13)? data_i[463] : 
                      (N8)? data_i[591] : 
                      (N10)? data_i[719] : 
                      (N12)? data_i[847] : 
                      (N14)? data_i[975] : 1'b0;
  assign data_o[78] = (N7)? data_i[78] : 
                      (N9)? data_i[206] : 
                      (N11)? data_i[334] : 
                      (N13)? data_i[462] : 
                      (N8)? data_i[590] : 
                      (N10)? data_i[718] : 
                      (N12)? data_i[846] : 
                      (N14)? data_i[974] : 1'b0;
  assign data_o[77] = (N7)? data_i[77] : 
                      (N9)? data_i[205] : 
                      (N11)? data_i[333] : 
                      (N13)? data_i[461] : 
                      (N8)? data_i[589] : 
                      (N10)? data_i[717] : 
                      (N12)? data_i[845] : 
                      (N14)? data_i[973] : 1'b0;
  assign data_o[76] = (N7)? data_i[76] : 
                      (N9)? data_i[204] : 
                      (N11)? data_i[332] : 
                      (N13)? data_i[460] : 
                      (N8)? data_i[588] : 
                      (N10)? data_i[716] : 
                      (N12)? data_i[844] : 
                      (N14)? data_i[972] : 1'b0;
  assign data_o[75] = (N7)? data_i[75] : 
                      (N9)? data_i[203] : 
                      (N11)? data_i[331] : 
                      (N13)? data_i[459] : 
                      (N8)? data_i[587] : 
                      (N10)? data_i[715] : 
                      (N12)? data_i[843] : 
                      (N14)? data_i[971] : 1'b0;
  assign data_o[74] = (N7)? data_i[74] : 
                      (N9)? data_i[202] : 
                      (N11)? data_i[330] : 
                      (N13)? data_i[458] : 
                      (N8)? data_i[586] : 
                      (N10)? data_i[714] : 
                      (N12)? data_i[842] : 
                      (N14)? data_i[970] : 1'b0;
  assign data_o[73] = (N7)? data_i[73] : 
                      (N9)? data_i[201] : 
                      (N11)? data_i[329] : 
                      (N13)? data_i[457] : 
                      (N8)? data_i[585] : 
                      (N10)? data_i[713] : 
                      (N12)? data_i[841] : 
                      (N14)? data_i[969] : 1'b0;
  assign data_o[72] = (N7)? data_i[72] : 
                      (N9)? data_i[200] : 
                      (N11)? data_i[328] : 
                      (N13)? data_i[456] : 
                      (N8)? data_i[584] : 
                      (N10)? data_i[712] : 
                      (N12)? data_i[840] : 
                      (N14)? data_i[968] : 1'b0;
  assign data_o[71] = (N7)? data_i[71] : 
                      (N9)? data_i[199] : 
                      (N11)? data_i[327] : 
                      (N13)? data_i[455] : 
                      (N8)? data_i[583] : 
                      (N10)? data_i[711] : 
                      (N12)? data_i[839] : 
                      (N14)? data_i[967] : 1'b0;
  assign data_o[70] = (N7)? data_i[70] : 
                      (N9)? data_i[198] : 
                      (N11)? data_i[326] : 
                      (N13)? data_i[454] : 
                      (N8)? data_i[582] : 
                      (N10)? data_i[710] : 
                      (N12)? data_i[838] : 
                      (N14)? data_i[966] : 1'b0;
  assign data_o[69] = (N7)? data_i[69] : 
                      (N9)? data_i[197] : 
                      (N11)? data_i[325] : 
                      (N13)? data_i[453] : 
                      (N8)? data_i[581] : 
                      (N10)? data_i[709] : 
                      (N12)? data_i[837] : 
                      (N14)? data_i[965] : 1'b0;
  assign data_o[68] = (N7)? data_i[68] : 
                      (N9)? data_i[196] : 
                      (N11)? data_i[324] : 
                      (N13)? data_i[452] : 
                      (N8)? data_i[580] : 
                      (N10)? data_i[708] : 
                      (N12)? data_i[836] : 
                      (N14)? data_i[964] : 1'b0;
  assign data_o[67] = (N7)? data_i[67] : 
                      (N9)? data_i[195] : 
                      (N11)? data_i[323] : 
                      (N13)? data_i[451] : 
                      (N8)? data_i[579] : 
                      (N10)? data_i[707] : 
                      (N12)? data_i[835] : 
                      (N14)? data_i[963] : 1'b0;
  assign data_o[66] = (N7)? data_i[66] : 
                      (N9)? data_i[194] : 
                      (N11)? data_i[322] : 
                      (N13)? data_i[450] : 
                      (N8)? data_i[578] : 
                      (N10)? data_i[706] : 
                      (N12)? data_i[834] : 
                      (N14)? data_i[962] : 1'b0;
  assign data_o[65] = (N7)? data_i[65] : 
                      (N9)? data_i[193] : 
                      (N11)? data_i[321] : 
                      (N13)? data_i[449] : 
                      (N8)? data_i[577] : 
                      (N10)? data_i[705] : 
                      (N12)? data_i[833] : 
                      (N14)? data_i[961] : 1'b0;
  assign data_o[64] = (N7)? data_i[64] : 
                      (N9)? data_i[192] : 
                      (N11)? data_i[320] : 
                      (N13)? data_i[448] : 
                      (N8)? data_i[576] : 
                      (N10)? data_i[704] : 
                      (N12)? data_i[832] : 
                      (N14)? data_i[960] : 1'b0;
  assign data_o[63] = (N7)? data_i[63] : 
                      (N9)? data_i[191] : 
                      (N11)? data_i[319] : 
                      (N13)? data_i[447] : 
                      (N8)? data_i[575] : 
                      (N10)? data_i[703] : 
                      (N12)? data_i[831] : 
                      (N14)? data_i[959] : 1'b0;
  assign data_o[62] = (N7)? data_i[62] : 
                      (N9)? data_i[190] : 
                      (N11)? data_i[318] : 
                      (N13)? data_i[446] : 
                      (N8)? data_i[574] : 
                      (N10)? data_i[702] : 
                      (N12)? data_i[830] : 
                      (N14)? data_i[958] : 1'b0;
  assign data_o[61] = (N7)? data_i[61] : 
                      (N9)? data_i[189] : 
                      (N11)? data_i[317] : 
                      (N13)? data_i[445] : 
                      (N8)? data_i[573] : 
                      (N10)? data_i[701] : 
                      (N12)? data_i[829] : 
                      (N14)? data_i[957] : 1'b0;
  assign data_o[60] = (N7)? data_i[60] : 
                      (N9)? data_i[188] : 
                      (N11)? data_i[316] : 
                      (N13)? data_i[444] : 
                      (N8)? data_i[572] : 
                      (N10)? data_i[700] : 
                      (N12)? data_i[828] : 
                      (N14)? data_i[956] : 1'b0;
  assign data_o[59] = (N7)? data_i[59] : 
                      (N9)? data_i[187] : 
                      (N11)? data_i[315] : 
                      (N13)? data_i[443] : 
                      (N8)? data_i[571] : 
                      (N10)? data_i[699] : 
                      (N12)? data_i[827] : 
                      (N14)? data_i[955] : 1'b0;
  assign data_o[58] = (N7)? data_i[58] : 
                      (N9)? data_i[186] : 
                      (N11)? data_i[314] : 
                      (N13)? data_i[442] : 
                      (N8)? data_i[570] : 
                      (N10)? data_i[698] : 
                      (N12)? data_i[826] : 
                      (N14)? data_i[954] : 1'b0;
  assign data_o[57] = (N7)? data_i[57] : 
                      (N9)? data_i[185] : 
                      (N11)? data_i[313] : 
                      (N13)? data_i[441] : 
                      (N8)? data_i[569] : 
                      (N10)? data_i[697] : 
                      (N12)? data_i[825] : 
                      (N14)? data_i[953] : 1'b0;
  assign data_o[56] = (N7)? data_i[56] : 
                      (N9)? data_i[184] : 
                      (N11)? data_i[312] : 
                      (N13)? data_i[440] : 
                      (N8)? data_i[568] : 
                      (N10)? data_i[696] : 
                      (N12)? data_i[824] : 
                      (N14)? data_i[952] : 1'b0;
  assign data_o[55] = (N7)? data_i[55] : 
                      (N9)? data_i[183] : 
                      (N11)? data_i[311] : 
                      (N13)? data_i[439] : 
                      (N8)? data_i[567] : 
                      (N10)? data_i[695] : 
                      (N12)? data_i[823] : 
                      (N14)? data_i[951] : 1'b0;
  assign data_o[54] = (N7)? data_i[54] : 
                      (N9)? data_i[182] : 
                      (N11)? data_i[310] : 
                      (N13)? data_i[438] : 
                      (N8)? data_i[566] : 
                      (N10)? data_i[694] : 
                      (N12)? data_i[822] : 
                      (N14)? data_i[950] : 1'b0;
  assign data_o[53] = (N7)? data_i[53] : 
                      (N9)? data_i[181] : 
                      (N11)? data_i[309] : 
                      (N13)? data_i[437] : 
                      (N8)? data_i[565] : 
                      (N10)? data_i[693] : 
                      (N12)? data_i[821] : 
                      (N14)? data_i[949] : 1'b0;
  assign data_o[52] = (N7)? data_i[52] : 
                      (N9)? data_i[180] : 
                      (N11)? data_i[308] : 
                      (N13)? data_i[436] : 
                      (N8)? data_i[564] : 
                      (N10)? data_i[692] : 
                      (N12)? data_i[820] : 
                      (N14)? data_i[948] : 1'b0;
  assign data_o[51] = (N7)? data_i[51] : 
                      (N9)? data_i[179] : 
                      (N11)? data_i[307] : 
                      (N13)? data_i[435] : 
                      (N8)? data_i[563] : 
                      (N10)? data_i[691] : 
                      (N12)? data_i[819] : 
                      (N14)? data_i[947] : 1'b0;
  assign data_o[50] = (N7)? data_i[50] : 
                      (N9)? data_i[178] : 
                      (N11)? data_i[306] : 
                      (N13)? data_i[434] : 
                      (N8)? data_i[562] : 
                      (N10)? data_i[690] : 
                      (N12)? data_i[818] : 
                      (N14)? data_i[946] : 1'b0;
  assign data_o[49] = (N7)? data_i[49] : 
                      (N9)? data_i[177] : 
                      (N11)? data_i[305] : 
                      (N13)? data_i[433] : 
                      (N8)? data_i[561] : 
                      (N10)? data_i[689] : 
                      (N12)? data_i[817] : 
                      (N14)? data_i[945] : 1'b0;
  assign data_o[48] = (N7)? data_i[48] : 
                      (N9)? data_i[176] : 
                      (N11)? data_i[304] : 
                      (N13)? data_i[432] : 
                      (N8)? data_i[560] : 
                      (N10)? data_i[688] : 
                      (N12)? data_i[816] : 
                      (N14)? data_i[944] : 1'b0;
  assign data_o[47] = (N7)? data_i[47] : 
                      (N9)? data_i[175] : 
                      (N11)? data_i[303] : 
                      (N13)? data_i[431] : 
                      (N8)? data_i[559] : 
                      (N10)? data_i[687] : 
                      (N12)? data_i[815] : 
                      (N14)? data_i[943] : 1'b0;
  assign data_o[46] = (N7)? data_i[46] : 
                      (N9)? data_i[174] : 
                      (N11)? data_i[302] : 
                      (N13)? data_i[430] : 
                      (N8)? data_i[558] : 
                      (N10)? data_i[686] : 
                      (N12)? data_i[814] : 
                      (N14)? data_i[942] : 1'b0;
  assign data_o[45] = (N7)? data_i[45] : 
                      (N9)? data_i[173] : 
                      (N11)? data_i[301] : 
                      (N13)? data_i[429] : 
                      (N8)? data_i[557] : 
                      (N10)? data_i[685] : 
                      (N12)? data_i[813] : 
                      (N14)? data_i[941] : 1'b0;
  assign data_o[44] = (N7)? data_i[44] : 
                      (N9)? data_i[172] : 
                      (N11)? data_i[300] : 
                      (N13)? data_i[428] : 
                      (N8)? data_i[556] : 
                      (N10)? data_i[684] : 
                      (N12)? data_i[812] : 
                      (N14)? data_i[940] : 1'b0;
  assign data_o[43] = (N7)? data_i[43] : 
                      (N9)? data_i[171] : 
                      (N11)? data_i[299] : 
                      (N13)? data_i[427] : 
                      (N8)? data_i[555] : 
                      (N10)? data_i[683] : 
                      (N12)? data_i[811] : 
                      (N14)? data_i[939] : 1'b0;
  assign data_o[42] = (N7)? data_i[42] : 
                      (N9)? data_i[170] : 
                      (N11)? data_i[298] : 
                      (N13)? data_i[426] : 
                      (N8)? data_i[554] : 
                      (N10)? data_i[682] : 
                      (N12)? data_i[810] : 
                      (N14)? data_i[938] : 1'b0;
  assign data_o[41] = (N7)? data_i[41] : 
                      (N9)? data_i[169] : 
                      (N11)? data_i[297] : 
                      (N13)? data_i[425] : 
                      (N8)? data_i[553] : 
                      (N10)? data_i[681] : 
                      (N12)? data_i[809] : 
                      (N14)? data_i[937] : 1'b0;
  assign data_o[40] = (N7)? data_i[40] : 
                      (N9)? data_i[168] : 
                      (N11)? data_i[296] : 
                      (N13)? data_i[424] : 
                      (N8)? data_i[552] : 
                      (N10)? data_i[680] : 
                      (N12)? data_i[808] : 
                      (N14)? data_i[936] : 1'b0;
  assign data_o[39] = (N7)? data_i[39] : 
                      (N9)? data_i[167] : 
                      (N11)? data_i[295] : 
                      (N13)? data_i[423] : 
                      (N8)? data_i[551] : 
                      (N10)? data_i[679] : 
                      (N12)? data_i[807] : 
                      (N14)? data_i[935] : 1'b0;
  assign data_o[38] = (N7)? data_i[38] : 
                      (N9)? data_i[166] : 
                      (N11)? data_i[294] : 
                      (N13)? data_i[422] : 
                      (N8)? data_i[550] : 
                      (N10)? data_i[678] : 
                      (N12)? data_i[806] : 
                      (N14)? data_i[934] : 1'b0;
  assign data_o[37] = (N7)? data_i[37] : 
                      (N9)? data_i[165] : 
                      (N11)? data_i[293] : 
                      (N13)? data_i[421] : 
                      (N8)? data_i[549] : 
                      (N10)? data_i[677] : 
                      (N12)? data_i[805] : 
                      (N14)? data_i[933] : 1'b0;
  assign data_o[36] = (N7)? data_i[36] : 
                      (N9)? data_i[164] : 
                      (N11)? data_i[292] : 
                      (N13)? data_i[420] : 
                      (N8)? data_i[548] : 
                      (N10)? data_i[676] : 
                      (N12)? data_i[804] : 
                      (N14)? data_i[932] : 1'b0;
  assign data_o[35] = (N7)? data_i[35] : 
                      (N9)? data_i[163] : 
                      (N11)? data_i[291] : 
                      (N13)? data_i[419] : 
                      (N8)? data_i[547] : 
                      (N10)? data_i[675] : 
                      (N12)? data_i[803] : 
                      (N14)? data_i[931] : 1'b0;
  assign data_o[34] = (N7)? data_i[34] : 
                      (N9)? data_i[162] : 
                      (N11)? data_i[290] : 
                      (N13)? data_i[418] : 
                      (N8)? data_i[546] : 
                      (N10)? data_i[674] : 
                      (N12)? data_i[802] : 
                      (N14)? data_i[930] : 1'b0;
  assign data_o[33] = (N7)? data_i[33] : 
                      (N9)? data_i[161] : 
                      (N11)? data_i[289] : 
                      (N13)? data_i[417] : 
                      (N8)? data_i[545] : 
                      (N10)? data_i[673] : 
                      (N12)? data_i[801] : 
                      (N14)? data_i[929] : 1'b0;
  assign data_o[32] = (N7)? data_i[32] : 
                      (N9)? data_i[160] : 
                      (N11)? data_i[288] : 
                      (N13)? data_i[416] : 
                      (N8)? data_i[544] : 
                      (N10)? data_i[672] : 
                      (N12)? data_i[800] : 
                      (N14)? data_i[928] : 1'b0;
  assign data_o[31] = (N7)? data_i[31] : 
                      (N9)? data_i[159] : 
                      (N11)? data_i[287] : 
                      (N13)? data_i[415] : 
                      (N8)? data_i[543] : 
                      (N10)? data_i[671] : 
                      (N12)? data_i[799] : 
                      (N14)? data_i[927] : 1'b0;
  assign data_o[30] = (N7)? data_i[30] : 
                      (N9)? data_i[158] : 
                      (N11)? data_i[286] : 
                      (N13)? data_i[414] : 
                      (N8)? data_i[542] : 
                      (N10)? data_i[670] : 
                      (N12)? data_i[798] : 
                      (N14)? data_i[926] : 1'b0;
  assign data_o[29] = (N7)? data_i[29] : 
                      (N9)? data_i[157] : 
                      (N11)? data_i[285] : 
                      (N13)? data_i[413] : 
                      (N8)? data_i[541] : 
                      (N10)? data_i[669] : 
                      (N12)? data_i[797] : 
                      (N14)? data_i[925] : 1'b0;
  assign data_o[28] = (N7)? data_i[28] : 
                      (N9)? data_i[156] : 
                      (N11)? data_i[284] : 
                      (N13)? data_i[412] : 
                      (N8)? data_i[540] : 
                      (N10)? data_i[668] : 
                      (N12)? data_i[796] : 
                      (N14)? data_i[924] : 1'b0;
  assign data_o[27] = (N7)? data_i[27] : 
                      (N9)? data_i[155] : 
                      (N11)? data_i[283] : 
                      (N13)? data_i[411] : 
                      (N8)? data_i[539] : 
                      (N10)? data_i[667] : 
                      (N12)? data_i[795] : 
                      (N14)? data_i[923] : 1'b0;
  assign data_o[26] = (N7)? data_i[26] : 
                      (N9)? data_i[154] : 
                      (N11)? data_i[282] : 
                      (N13)? data_i[410] : 
                      (N8)? data_i[538] : 
                      (N10)? data_i[666] : 
                      (N12)? data_i[794] : 
                      (N14)? data_i[922] : 1'b0;
  assign data_o[25] = (N7)? data_i[25] : 
                      (N9)? data_i[153] : 
                      (N11)? data_i[281] : 
                      (N13)? data_i[409] : 
                      (N8)? data_i[537] : 
                      (N10)? data_i[665] : 
                      (N12)? data_i[793] : 
                      (N14)? data_i[921] : 1'b0;
  assign data_o[24] = (N7)? data_i[24] : 
                      (N9)? data_i[152] : 
                      (N11)? data_i[280] : 
                      (N13)? data_i[408] : 
                      (N8)? data_i[536] : 
                      (N10)? data_i[664] : 
                      (N12)? data_i[792] : 
                      (N14)? data_i[920] : 1'b0;
  assign data_o[23] = (N7)? data_i[23] : 
                      (N9)? data_i[151] : 
                      (N11)? data_i[279] : 
                      (N13)? data_i[407] : 
                      (N8)? data_i[535] : 
                      (N10)? data_i[663] : 
                      (N12)? data_i[791] : 
                      (N14)? data_i[919] : 1'b0;
  assign data_o[22] = (N7)? data_i[22] : 
                      (N9)? data_i[150] : 
                      (N11)? data_i[278] : 
                      (N13)? data_i[406] : 
                      (N8)? data_i[534] : 
                      (N10)? data_i[662] : 
                      (N12)? data_i[790] : 
                      (N14)? data_i[918] : 1'b0;
  assign data_o[21] = (N7)? data_i[21] : 
                      (N9)? data_i[149] : 
                      (N11)? data_i[277] : 
                      (N13)? data_i[405] : 
                      (N8)? data_i[533] : 
                      (N10)? data_i[661] : 
                      (N12)? data_i[789] : 
                      (N14)? data_i[917] : 1'b0;
  assign data_o[20] = (N7)? data_i[20] : 
                      (N9)? data_i[148] : 
                      (N11)? data_i[276] : 
                      (N13)? data_i[404] : 
                      (N8)? data_i[532] : 
                      (N10)? data_i[660] : 
                      (N12)? data_i[788] : 
                      (N14)? data_i[916] : 1'b0;
  assign data_o[19] = (N7)? data_i[19] : 
                      (N9)? data_i[147] : 
                      (N11)? data_i[275] : 
                      (N13)? data_i[403] : 
                      (N8)? data_i[531] : 
                      (N10)? data_i[659] : 
                      (N12)? data_i[787] : 
                      (N14)? data_i[915] : 1'b0;
  assign data_o[18] = (N7)? data_i[18] : 
                      (N9)? data_i[146] : 
                      (N11)? data_i[274] : 
                      (N13)? data_i[402] : 
                      (N8)? data_i[530] : 
                      (N10)? data_i[658] : 
                      (N12)? data_i[786] : 
                      (N14)? data_i[914] : 1'b0;
  assign data_o[17] = (N7)? data_i[17] : 
                      (N9)? data_i[145] : 
                      (N11)? data_i[273] : 
                      (N13)? data_i[401] : 
                      (N8)? data_i[529] : 
                      (N10)? data_i[657] : 
                      (N12)? data_i[785] : 
                      (N14)? data_i[913] : 1'b0;
  assign data_o[16] = (N7)? data_i[16] : 
                      (N9)? data_i[144] : 
                      (N11)? data_i[272] : 
                      (N13)? data_i[400] : 
                      (N8)? data_i[528] : 
                      (N10)? data_i[656] : 
                      (N12)? data_i[784] : 
                      (N14)? data_i[912] : 1'b0;
  assign data_o[15] = (N7)? data_i[15] : 
                      (N9)? data_i[143] : 
                      (N11)? data_i[271] : 
                      (N13)? data_i[399] : 
                      (N8)? data_i[527] : 
                      (N10)? data_i[655] : 
                      (N12)? data_i[783] : 
                      (N14)? data_i[911] : 1'b0;
  assign data_o[14] = (N7)? data_i[14] : 
                      (N9)? data_i[142] : 
                      (N11)? data_i[270] : 
                      (N13)? data_i[398] : 
                      (N8)? data_i[526] : 
                      (N10)? data_i[654] : 
                      (N12)? data_i[782] : 
                      (N14)? data_i[910] : 1'b0;
  assign data_o[13] = (N7)? data_i[13] : 
                      (N9)? data_i[141] : 
                      (N11)? data_i[269] : 
                      (N13)? data_i[397] : 
                      (N8)? data_i[525] : 
                      (N10)? data_i[653] : 
                      (N12)? data_i[781] : 
                      (N14)? data_i[909] : 1'b0;
  assign data_o[12] = (N7)? data_i[12] : 
                      (N9)? data_i[140] : 
                      (N11)? data_i[268] : 
                      (N13)? data_i[396] : 
                      (N8)? data_i[524] : 
                      (N10)? data_i[652] : 
                      (N12)? data_i[780] : 
                      (N14)? data_i[908] : 1'b0;
  assign data_o[11] = (N7)? data_i[11] : 
                      (N9)? data_i[139] : 
                      (N11)? data_i[267] : 
                      (N13)? data_i[395] : 
                      (N8)? data_i[523] : 
                      (N10)? data_i[651] : 
                      (N12)? data_i[779] : 
                      (N14)? data_i[907] : 1'b0;
  assign data_o[10] = (N7)? data_i[10] : 
                      (N9)? data_i[138] : 
                      (N11)? data_i[266] : 
                      (N13)? data_i[394] : 
                      (N8)? data_i[522] : 
                      (N10)? data_i[650] : 
                      (N12)? data_i[778] : 
                      (N14)? data_i[906] : 1'b0;
  assign data_o[9] = (N7)? data_i[9] : 
                     (N9)? data_i[137] : 
                     (N11)? data_i[265] : 
                     (N13)? data_i[393] : 
                     (N8)? data_i[521] : 
                     (N10)? data_i[649] : 
                     (N12)? data_i[777] : 
                     (N14)? data_i[905] : 1'b0;
  assign data_o[8] = (N7)? data_i[8] : 
                     (N9)? data_i[136] : 
                     (N11)? data_i[264] : 
                     (N13)? data_i[392] : 
                     (N8)? data_i[520] : 
                     (N10)? data_i[648] : 
                     (N12)? data_i[776] : 
                     (N14)? data_i[904] : 1'b0;
  assign data_o[7] = (N7)? data_i[7] : 
                     (N9)? data_i[135] : 
                     (N11)? data_i[263] : 
                     (N13)? data_i[391] : 
                     (N8)? data_i[519] : 
                     (N10)? data_i[647] : 
                     (N12)? data_i[775] : 
                     (N14)? data_i[903] : 1'b0;
  assign data_o[6] = (N7)? data_i[6] : 
                     (N9)? data_i[134] : 
                     (N11)? data_i[262] : 
                     (N13)? data_i[390] : 
                     (N8)? data_i[518] : 
                     (N10)? data_i[646] : 
                     (N12)? data_i[774] : 
                     (N14)? data_i[902] : 1'b0;
  assign data_o[5] = (N7)? data_i[5] : 
                     (N9)? data_i[133] : 
                     (N11)? data_i[261] : 
                     (N13)? data_i[389] : 
                     (N8)? data_i[517] : 
                     (N10)? data_i[645] : 
                     (N12)? data_i[773] : 
                     (N14)? data_i[901] : 1'b0;
  assign data_o[4] = (N7)? data_i[4] : 
                     (N9)? data_i[132] : 
                     (N11)? data_i[260] : 
                     (N13)? data_i[388] : 
                     (N8)? data_i[516] : 
                     (N10)? data_i[644] : 
                     (N12)? data_i[772] : 
                     (N14)? data_i[900] : 1'b0;
  assign data_o[3] = (N7)? data_i[3] : 
                     (N9)? data_i[131] : 
                     (N11)? data_i[259] : 
                     (N13)? data_i[387] : 
                     (N8)? data_i[515] : 
                     (N10)? data_i[643] : 
                     (N12)? data_i[771] : 
                     (N14)? data_i[899] : 1'b0;
  assign data_o[2] = (N7)? data_i[2] : 
                     (N9)? data_i[130] : 
                     (N11)? data_i[258] : 
                     (N13)? data_i[386] : 
                     (N8)? data_i[514] : 
                     (N10)? data_i[642] : 
                     (N12)? data_i[770] : 
                     (N14)? data_i[898] : 1'b0;
  assign data_o[1] = (N7)? data_i[1] : 
                     (N9)? data_i[129] : 
                     (N11)? data_i[257] : 
                     (N13)? data_i[385] : 
                     (N8)? data_i[513] : 
                     (N10)? data_i[641] : 
                     (N12)? data_i[769] : 
                     (N14)? data_i[897] : 1'b0;
  assign data_o[0] = (N7)? data_i[0] : 
                     (N9)? data_i[128] : 
                     (N11)? data_i[256] : 
                     (N13)? data_i[384] : 
                     (N8)? data_i[512] : 
                     (N10)? data_i[640] : 
                     (N12)? data_i[768] : 
                     (N14)? data_i[896] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];
  assign N6 = ~sel_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & sel_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & sel_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & sel_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & sel_i[2];

endmodule



module bsg_bus_pack_00000080
(
  data_i,
  sel_i,
  size_i,
  data_o
);

  input [127:0] data_i;
  input [3:0] sel_i;
  input [2:0] size_i;
  output [127:0] data_o;
  wire [127:0] data_o,data_rot_lo;
  wire data_repl_lo_7__127_,data_repl_lo_7__126_,data_repl_lo_7__125_,
  data_repl_lo_7__124_,data_repl_lo_7__123_,data_repl_lo_7__122_,data_repl_lo_7__121_,
  data_repl_lo_7__120_,data_repl_lo_7__119_,data_repl_lo_7__118_,data_repl_lo_7__117_,
  data_repl_lo_7__116_,data_repl_lo_7__115_,data_repl_lo_7__114_,data_repl_lo_7__113_,
  data_repl_lo_7__112_,data_repl_lo_7__111_,data_repl_lo_7__110_,data_repl_lo_7__109_,
  data_repl_lo_7__108_,data_repl_lo_7__107_,data_repl_lo_7__106_,
  data_repl_lo_7__105_,data_repl_lo_7__104_,data_repl_lo_7__103_,data_repl_lo_7__102_,
  data_repl_lo_7__101_,data_repl_lo_7__100_,data_repl_lo_7__99_,data_repl_lo_7__98_,
  data_repl_lo_7__97_,data_repl_lo_7__96_,data_repl_lo_7__95_,data_repl_lo_7__94_,
  data_repl_lo_7__93_,data_repl_lo_7__92_,data_repl_lo_7__91_,data_repl_lo_7__90_,
  data_repl_lo_7__89_,data_repl_lo_7__88_,data_repl_lo_7__87_,data_repl_lo_7__86_,
  data_repl_lo_7__85_,data_repl_lo_7__84_,data_repl_lo_7__83_,data_repl_lo_7__82_,
  data_repl_lo_7__81_,data_repl_lo_7__80_,data_repl_lo_7__79_,data_repl_lo_7__78_,
  data_repl_lo_7__77_,data_repl_lo_7__76_,data_repl_lo_7__75_,data_repl_lo_7__74_,
  data_repl_lo_7__73_,data_repl_lo_7__72_,data_repl_lo_7__71_,data_repl_lo_7__70_,
  data_repl_lo_7__69_,data_repl_lo_7__68_,data_repl_lo_7__67_,data_repl_lo_7__66_,
  data_repl_lo_7__65_,data_repl_lo_7__64_,data_repl_lo_7__63_,data_repl_lo_7__62_,
  data_repl_lo_7__61_,data_repl_lo_7__60_,data_repl_lo_7__59_,data_repl_lo_7__58_,
  data_repl_lo_7__57_,data_repl_lo_7__56_,data_repl_lo_7__55_,data_repl_lo_7__54_,
  data_repl_lo_7__53_,data_repl_lo_7__52_,data_repl_lo_7__51_,data_repl_lo_7__50_,
  data_repl_lo_7__49_,data_repl_lo_7__48_,data_repl_lo_7__47_,data_repl_lo_7__46_,
  data_repl_lo_7__45_,data_repl_lo_7__44_,data_repl_lo_7__43_,data_repl_lo_7__42_,
  data_repl_lo_7__41_,data_repl_lo_7__40_,data_repl_lo_7__39_,data_repl_lo_7__38_,
  data_repl_lo_7__37_,data_repl_lo_7__36_,data_repl_lo_7__35_,data_repl_lo_7__34_,
  data_repl_lo_7__33_,data_repl_lo_7__32_,data_repl_lo_7__31_,data_repl_lo_7__30_,
  data_repl_lo_7__29_,data_repl_lo_7__28_,data_repl_lo_7__27_,data_repl_lo_7__26_,
  data_repl_lo_7__25_,data_repl_lo_7__24_,data_repl_lo_7__23_,data_repl_lo_7__22_,
  data_repl_lo_7__21_,data_repl_lo_7__20_,data_repl_lo_7__19_,data_repl_lo_7__18_,
  data_repl_lo_7__17_,data_repl_lo_7__16_,data_repl_lo_7__15_,data_repl_lo_7__14_,
  data_repl_lo_7__13_,data_repl_lo_7__12_,data_repl_lo_7__11_,data_repl_lo_7__10_,
  data_repl_lo_7__9_,data_repl_lo_7__8_,data_repl_lo_7__7_,data_repl_lo_7__6_,
  data_repl_lo_7__5_,data_repl_lo_7__4_,data_repl_lo_7__3_,data_repl_lo_7__2_,data_repl_lo_7__1_,
  data_repl_lo_7__0_,data_repl_lo_6__127_,data_repl_lo_6__126_,
  data_repl_lo_6__125_,data_repl_lo_6__124_,data_repl_lo_6__123_,data_repl_lo_6__122_,
  data_repl_lo_6__121_,data_repl_lo_6__120_,data_repl_lo_6__119_,data_repl_lo_6__118_,
  data_repl_lo_6__117_,data_repl_lo_6__116_,data_repl_lo_6__115_,data_repl_lo_6__114_,
  data_repl_lo_6__113_,data_repl_lo_6__112_,data_repl_lo_6__111_,data_repl_lo_6__110_,
  data_repl_lo_6__109_,data_repl_lo_6__108_,data_repl_lo_6__107_,data_repl_lo_6__106_,
  data_repl_lo_6__105_,data_repl_lo_6__104_,data_repl_lo_6__103_,
  data_repl_lo_6__102_,data_repl_lo_6__101_,data_repl_lo_6__100_,data_repl_lo_6__99_,
  data_repl_lo_6__98_,data_repl_lo_6__97_,data_repl_lo_6__96_,data_repl_lo_6__95_,
  data_repl_lo_6__94_,data_repl_lo_6__93_,data_repl_lo_6__92_,data_repl_lo_6__91_,
  data_repl_lo_6__90_,data_repl_lo_6__89_,data_repl_lo_6__88_,data_repl_lo_6__87_,
  data_repl_lo_6__86_,data_repl_lo_6__85_,data_repl_lo_6__84_,data_repl_lo_6__83_,
  data_repl_lo_6__82_,data_repl_lo_6__81_,data_repl_lo_6__80_,data_repl_lo_6__79_,
  data_repl_lo_6__78_,data_repl_lo_6__77_,data_repl_lo_6__76_,data_repl_lo_6__75_,
  data_repl_lo_6__74_,data_repl_lo_6__73_,data_repl_lo_6__72_,data_repl_lo_6__71_,
  data_repl_lo_6__70_,data_repl_lo_6__69_,data_repl_lo_6__68_,data_repl_lo_6__67_,
  data_repl_lo_6__66_,data_repl_lo_6__65_,data_repl_lo_6__64_,data_repl_lo_6__63_,
  data_repl_lo_6__62_,data_repl_lo_6__61_,data_repl_lo_6__60_,data_repl_lo_6__59_,
  data_repl_lo_6__58_,data_repl_lo_6__57_,data_repl_lo_6__56_,data_repl_lo_6__55_,
  data_repl_lo_6__54_,data_repl_lo_6__53_,data_repl_lo_6__52_,data_repl_lo_6__51_,
  data_repl_lo_6__50_,data_repl_lo_6__49_,data_repl_lo_6__48_,data_repl_lo_6__47_,
  data_repl_lo_6__46_,data_repl_lo_6__45_,data_repl_lo_6__44_,data_repl_lo_6__43_,
  data_repl_lo_6__42_,data_repl_lo_6__41_,data_repl_lo_6__40_,data_repl_lo_6__39_,
  data_repl_lo_6__38_,data_repl_lo_6__37_,data_repl_lo_6__36_,data_repl_lo_6__35_,
  data_repl_lo_6__34_,data_repl_lo_6__33_,data_repl_lo_6__32_,data_repl_lo_6__31_,
  data_repl_lo_6__30_,data_repl_lo_6__29_,data_repl_lo_6__28_,data_repl_lo_6__27_,
  data_repl_lo_6__26_,data_repl_lo_6__25_,data_repl_lo_6__24_,data_repl_lo_6__23_,
  data_repl_lo_6__22_,data_repl_lo_6__21_,data_repl_lo_6__20_,data_repl_lo_6__19_,
  data_repl_lo_6__18_,data_repl_lo_6__17_,data_repl_lo_6__16_,data_repl_lo_6__15_,
  data_repl_lo_6__14_,data_repl_lo_6__13_,data_repl_lo_6__12_,data_repl_lo_6__11_,
  data_repl_lo_6__10_,data_repl_lo_6__9_,data_repl_lo_6__8_,data_repl_lo_6__7_,
  data_repl_lo_6__6_,data_repl_lo_6__5_,data_repl_lo_6__4_,data_repl_lo_6__3_,data_repl_lo_6__2_,
  data_repl_lo_6__1_,data_repl_lo_6__0_,data_repl_lo_5__127_,data_repl_lo_5__126_,
  data_repl_lo_5__125_,data_repl_lo_5__124_,data_repl_lo_5__123_,
  data_repl_lo_5__122_,data_repl_lo_5__121_,data_repl_lo_5__120_,data_repl_lo_5__119_,
  data_repl_lo_5__118_,data_repl_lo_5__117_,data_repl_lo_5__116_,data_repl_lo_5__115_,
  data_repl_lo_5__114_,data_repl_lo_5__113_,data_repl_lo_5__112_,data_repl_lo_5__111_,
  data_repl_lo_5__110_,data_repl_lo_5__109_,data_repl_lo_5__108_,data_repl_lo_5__107_,
  data_repl_lo_5__106_,data_repl_lo_5__105_,data_repl_lo_5__104_,
  data_repl_lo_5__103_,data_repl_lo_5__102_,data_repl_lo_5__101_,data_repl_lo_5__100_,
  data_repl_lo_5__99_,data_repl_lo_5__98_,data_repl_lo_5__97_,data_repl_lo_5__96_,
  data_repl_lo_5__95_,data_repl_lo_5__94_,data_repl_lo_5__93_,data_repl_lo_5__92_,
  data_repl_lo_5__91_,data_repl_lo_5__90_,data_repl_lo_5__89_,data_repl_lo_5__88_,
  data_repl_lo_5__87_,data_repl_lo_5__86_,data_repl_lo_5__85_,data_repl_lo_5__84_,
  data_repl_lo_5__83_,data_repl_lo_5__82_,data_repl_lo_5__81_,data_repl_lo_5__80_,
  data_repl_lo_5__79_,data_repl_lo_5__78_,data_repl_lo_5__77_,data_repl_lo_5__76_,
  data_repl_lo_5__75_,data_repl_lo_5__74_,data_repl_lo_5__73_,data_repl_lo_5__72_,
  data_repl_lo_5__71_,data_repl_lo_5__70_,data_repl_lo_5__69_,data_repl_lo_5__68_,
  data_repl_lo_5__67_,data_repl_lo_5__66_,data_repl_lo_5__65_,data_repl_lo_5__64_,
  data_repl_lo_5__63_,data_repl_lo_5__62_,data_repl_lo_5__61_,data_repl_lo_5__60_,
  data_repl_lo_5__59_,data_repl_lo_5__58_,data_repl_lo_5__57_,data_repl_lo_5__56_,
  data_repl_lo_5__55_,data_repl_lo_5__54_,data_repl_lo_5__53_,data_repl_lo_5__52_,
  data_repl_lo_5__51_,data_repl_lo_5__50_,data_repl_lo_5__49_,data_repl_lo_5__48_,
  data_repl_lo_5__47_,data_repl_lo_5__46_,data_repl_lo_5__45_,data_repl_lo_5__44_,
  data_repl_lo_5__43_,data_repl_lo_5__42_,data_repl_lo_5__41_,data_repl_lo_5__40_,
  data_repl_lo_5__39_,data_repl_lo_5__38_,data_repl_lo_5__37_,data_repl_lo_5__36_,
  data_repl_lo_5__35_,data_repl_lo_5__34_,data_repl_lo_5__33_,data_repl_lo_5__32_,
  data_repl_lo_5__31_,data_repl_lo_5__30_,data_repl_lo_5__29_,data_repl_lo_5__28_,
  data_repl_lo_5__27_,data_repl_lo_5__26_,data_repl_lo_5__25_,data_repl_lo_5__24_,
  data_repl_lo_5__23_,data_repl_lo_5__22_,data_repl_lo_5__21_,data_repl_lo_5__20_,
  data_repl_lo_5__19_,data_repl_lo_5__18_,data_repl_lo_5__17_,data_repl_lo_5__16_,
  data_repl_lo_5__15_,data_repl_lo_5__14_,data_repl_lo_5__13_,data_repl_lo_5__12_,
  data_repl_lo_5__11_,data_repl_lo_5__10_,data_repl_lo_5__9_,data_repl_lo_5__8_,
  data_repl_lo_5__7_,data_repl_lo_5__6_,data_repl_lo_5__5_,data_repl_lo_5__4_,data_repl_lo_5__3_,
  data_repl_lo_5__2_,data_repl_lo_5__1_,data_repl_lo_5__0_;

  bsg_rotate_right_00000080
  rot
  (
    .data_i(data_i),
    .rot_i({ sel_i, 1'b0, 1'b0, 1'b0 }),
    .o(data_rot_lo)
  );


  bsg_mux_00000080_00000008
  repl_mux
  (
    .data_i({ data_repl_lo_7__127_, data_repl_lo_7__126_, data_repl_lo_7__125_, data_repl_lo_7__124_, data_repl_lo_7__123_, data_repl_lo_7__122_, data_repl_lo_7__121_, data_repl_lo_7__120_, data_repl_lo_7__119_, data_repl_lo_7__118_, data_repl_lo_7__117_, data_repl_lo_7__116_, data_repl_lo_7__115_, data_repl_lo_7__114_, data_repl_lo_7__113_, data_repl_lo_7__112_, data_repl_lo_7__111_, data_repl_lo_7__110_, data_repl_lo_7__109_, data_repl_lo_7__108_, data_repl_lo_7__107_, data_repl_lo_7__106_, data_repl_lo_7__105_, data_repl_lo_7__104_, data_repl_lo_7__103_, data_repl_lo_7__102_, data_repl_lo_7__101_, data_repl_lo_7__100_, data_repl_lo_7__99_, data_repl_lo_7__98_, data_repl_lo_7__97_, data_repl_lo_7__96_, data_repl_lo_7__95_, data_repl_lo_7__94_, data_repl_lo_7__93_, data_repl_lo_7__92_, data_repl_lo_7__91_, data_repl_lo_7__90_, data_repl_lo_7__89_, data_repl_lo_7__88_, data_repl_lo_7__87_, data_repl_lo_7__86_, data_repl_lo_7__85_, data_repl_lo_7__84_, data_repl_lo_7__83_, data_repl_lo_7__82_, data_repl_lo_7__81_, data_repl_lo_7__80_, data_repl_lo_7__79_, data_repl_lo_7__78_, data_repl_lo_7__77_, data_repl_lo_7__76_, data_repl_lo_7__75_, data_repl_lo_7__74_, data_repl_lo_7__73_, data_repl_lo_7__72_, data_repl_lo_7__71_, data_repl_lo_7__70_, data_repl_lo_7__69_, data_repl_lo_7__68_, data_repl_lo_7__67_, data_repl_lo_7__66_, data_repl_lo_7__65_, data_repl_lo_7__64_, data_repl_lo_7__63_, data_repl_lo_7__62_, data_repl_lo_7__61_, data_repl_lo_7__60_, data_repl_lo_7__59_, data_repl_lo_7__58_, data_repl_lo_7__57_, data_repl_lo_7__56_, data_repl_lo_7__55_, data_repl_lo_7__54_, data_repl_lo_7__53_, data_repl_lo_7__52_, data_repl_lo_7__51_, data_repl_lo_7__50_, data_repl_lo_7__49_, data_repl_lo_7__48_, data_repl_lo_7__47_, data_repl_lo_7__46_, data_repl_lo_7__45_, data_repl_lo_7__44_, data_repl_lo_7__43_, data_repl_lo_7__42_, data_repl_lo_7__41_, data_repl_lo_7__40_, data_repl_lo_7__39_, data_repl_lo_7__38_, data_repl_lo_7__37_, data_repl_lo_7__36_, data_repl_lo_7__35_, data_repl_lo_7__34_, data_repl_lo_7__33_, data_repl_lo_7__32_, data_repl_lo_7__31_, data_repl_lo_7__30_, data_repl_lo_7__29_, data_repl_lo_7__28_, data_repl_lo_7__27_, data_repl_lo_7__26_, data_repl_lo_7__25_, data_repl_lo_7__24_, data_repl_lo_7__23_, data_repl_lo_7__22_, data_repl_lo_7__21_, data_repl_lo_7__20_, data_repl_lo_7__19_, data_repl_lo_7__18_, data_repl_lo_7__17_, data_repl_lo_7__16_, data_repl_lo_7__15_, data_repl_lo_7__14_, data_repl_lo_7__13_, data_repl_lo_7__12_, data_repl_lo_7__11_, data_repl_lo_7__10_, data_repl_lo_7__9_, data_repl_lo_7__8_, data_repl_lo_7__7_, data_repl_lo_7__6_, data_repl_lo_7__5_, data_repl_lo_7__4_, data_repl_lo_7__3_, data_repl_lo_7__2_, data_repl_lo_7__1_, data_repl_lo_7__0_, data_repl_lo_6__127_, data_repl_lo_6__126_, data_repl_lo_6__125_, data_repl_lo_6__124_, data_repl_lo_6__123_, data_repl_lo_6__122_, data_repl_lo_6__121_, data_repl_lo_6__120_, data_repl_lo_6__119_, data_repl_lo_6__118_, data_repl_lo_6__117_, data_repl_lo_6__116_, data_repl_lo_6__115_, data_repl_lo_6__114_, data_repl_lo_6__113_, data_repl_lo_6__112_, data_repl_lo_6__111_, data_repl_lo_6__110_, data_repl_lo_6__109_, data_repl_lo_6__108_, data_repl_lo_6__107_, data_repl_lo_6__106_, data_repl_lo_6__105_, data_repl_lo_6__104_, data_repl_lo_6__103_, data_repl_lo_6__102_, data_repl_lo_6__101_, data_repl_lo_6__100_, data_repl_lo_6__99_, data_repl_lo_6__98_, data_repl_lo_6__97_, data_repl_lo_6__96_, data_repl_lo_6__95_, data_repl_lo_6__94_, data_repl_lo_6__93_, data_repl_lo_6__92_, data_repl_lo_6__91_, data_repl_lo_6__90_, data_repl_lo_6__89_, data_repl_lo_6__88_, data_repl_lo_6__87_, data_repl_lo_6__86_, data_repl_lo_6__85_, data_repl_lo_6__84_, data_repl_lo_6__83_, data_repl_lo_6__82_, data_repl_lo_6__81_, data_repl_lo_6__80_, data_repl_lo_6__79_, data_repl_lo_6__78_, data_repl_lo_6__77_, data_repl_lo_6__76_, data_repl_lo_6__75_, data_repl_lo_6__74_, data_repl_lo_6__73_, data_repl_lo_6__72_, data_repl_lo_6__71_, data_repl_lo_6__70_, data_repl_lo_6__69_, data_repl_lo_6__68_, data_repl_lo_6__67_, data_repl_lo_6__66_, data_repl_lo_6__65_, data_repl_lo_6__64_, data_repl_lo_6__63_, data_repl_lo_6__62_, data_repl_lo_6__61_, data_repl_lo_6__60_, data_repl_lo_6__59_, data_repl_lo_6__58_, data_repl_lo_6__57_, data_repl_lo_6__56_, data_repl_lo_6__55_, data_repl_lo_6__54_, data_repl_lo_6__53_, data_repl_lo_6__52_, data_repl_lo_6__51_, data_repl_lo_6__50_, data_repl_lo_6__49_, data_repl_lo_6__48_, data_repl_lo_6__47_, data_repl_lo_6__46_, data_repl_lo_6__45_, data_repl_lo_6__44_, data_repl_lo_6__43_, data_repl_lo_6__42_, data_repl_lo_6__41_, data_repl_lo_6__40_, data_repl_lo_6__39_, data_repl_lo_6__38_, data_repl_lo_6__37_, data_repl_lo_6__36_, data_repl_lo_6__35_, data_repl_lo_6__34_, data_repl_lo_6__33_, data_repl_lo_6__32_, data_repl_lo_6__31_, data_repl_lo_6__30_, data_repl_lo_6__29_, data_repl_lo_6__28_, data_repl_lo_6__27_, data_repl_lo_6__26_, data_repl_lo_6__25_, data_repl_lo_6__24_, data_repl_lo_6__23_, data_repl_lo_6__22_, data_repl_lo_6__21_, data_repl_lo_6__20_, data_repl_lo_6__19_, data_repl_lo_6__18_, data_repl_lo_6__17_, data_repl_lo_6__16_, data_repl_lo_6__15_, data_repl_lo_6__14_, data_repl_lo_6__13_, data_repl_lo_6__12_, data_repl_lo_6__11_, data_repl_lo_6__10_, data_repl_lo_6__9_, data_repl_lo_6__8_, data_repl_lo_6__7_, data_repl_lo_6__6_, data_repl_lo_6__5_, data_repl_lo_6__4_, data_repl_lo_6__3_, data_repl_lo_6__2_, data_repl_lo_6__1_, data_repl_lo_6__0_, data_repl_lo_5__127_, data_repl_lo_5__126_, data_repl_lo_5__125_, data_repl_lo_5__124_, data_repl_lo_5__123_, data_repl_lo_5__122_, data_repl_lo_5__121_, data_repl_lo_5__120_, data_repl_lo_5__119_, data_repl_lo_5__118_, data_repl_lo_5__117_, data_repl_lo_5__116_, data_repl_lo_5__115_, data_repl_lo_5__114_, data_repl_lo_5__113_, data_repl_lo_5__112_, data_repl_lo_5__111_, data_repl_lo_5__110_, data_repl_lo_5__109_, data_repl_lo_5__108_, data_repl_lo_5__107_, data_repl_lo_5__106_, data_repl_lo_5__105_, data_repl_lo_5__104_, data_repl_lo_5__103_, data_repl_lo_5__102_, data_repl_lo_5__101_, data_repl_lo_5__100_, data_repl_lo_5__99_, data_repl_lo_5__98_, data_repl_lo_5__97_, data_repl_lo_5__96_, data_repl_lo_5__95_, data_repl_lo_5__94_, data_repl_lo_5__93_, data_repl_lo_5__92_, data_repl_lo_5__91_, data_repl_lo_5__90_, data_repl_lo_5__89_, data_repl_lo_5__88_, data_repl_lo_5__87_, data_repl_lo_5__86_, data_repl_lo_5__85_, data_repl_lo_5__84_, data_repl_lo_5__83_, data_repl_lo_5__82_, data_repl_lo_5__81_, data_repl_lo_5__80_, data_repl_lo_5__79_, data_repl_lo_5__78_, data_repl_lo_5__77_, data_repl_lo_5__76_, data_repl_lo_5__75_, data_repl_lo_5__74_, data_repl_lo_5__73_, data_repl_lo_5__72_, data_repl_lo_5__71_, data_repl_lo_5__70_, data_repl_lo_5__69_, data_repl_lo_5__68_, data_repl_lo_5__67_, data_repl_lo_5__66_, data_repl_lo_5__65_, data_repl_lo_5__64_, data_repl_lo_5__63_, data_repl_lo_5__62_, data_repl_lo_5__61_, data_repl_lo_5__60_, data_repl_lo_5__59_, data_repl_lo_5__58_, data_repl_lo_5__57_, data_repl_lo_5__56_, data_repl_lo_5__55_, data_repl_lo_5__54_, data_repl_lo_5__53_, data_repl_lo_5__52_, data_repl_lo_5__51_, data_repl_lo_5__50_, data_repl_lo_5__49_, data_repl_lo_5__48_, data_repl_lo_5__47_, data_repl_lo_5__46_, data_repl_lo_5__45_, data_repl_lo_5__44_, data_repl_lo_5__43_, data_repl_lo_5__42_, data_repl_lo_5__41_, data_repl_lo_5__40_, data_repl_lo_5__39_, data_repl_lo_5__38_, data_repl_lo_5__37_, data_repl_lo_5__36_, data_repl_lo_5__35_, data_repl_lo_5__34_, data_repl_lo_5__33_, data_repl_lo_5__32_, data_repl_lo_5__31_, data_repl_lo_5__30_, data_repl_lo_5__29_, data_repl_lo_5__28_, data_repl_lo_5__27_, data_repl_lo_5__26_, data_repl_lo_5__25_, data_repl_lo_5__24_, data_repl_lo_5__23_, data_repl_lo_5__22_, data_repl_lo_5__21_, data_repl_lo_5__20_, data_repl_lo_5__19_, data_repl_lo_5__18_, data_repl_lo_5__17_, data_repl_lo_5__16_, data_repl_lo_5__15_, data_repl_lo_5__14_, data_repl_lo_5__13_, data_repl_lo_5__12_, data_repl_lo_5__11_, data_repl_lo_5__10_, data_repl_lo_5__9_, data_repl_lo_5__8_, data_repl_lo_5__7_, data_repl_lo_5__6_, data_repl_lo_5__5_, data_repl_lo_5__4_, data_repl_lo_5__3_, data_repl_lo_5__2_, data_repl_lo_5__1_, data_repl_lo_5__0_, data_rot_lo, data_rot_lo[63:0], data_rot_lo[63:0], data_rot_lo[31:0], data_rot_lo[31:0], data_rot_lo[31:0], data_rot_lo[31:0], data_rot_lo[15:0], data_rot_lo[15:0], data_rot_lo[15:0], data_rot_lo[15:0], data_rot_lo[15:0], data_rot_lo[15:0], data_rot_lo[15:0], data_rot_lo[15:0], data_rot_lo[7:0], data_rot_lo[7:0], data_rot_lo[7:0], data_rot_lo[7:0], data_rot_lo[7:0], data_rot_lo[7:0], data_rot_lo[7:0], data_rot_lo[7:0], data_rot_lo[7:0], data_rot_lo[7:0], data_rot_lo[7:0], data_rot_lo[7:0], data_rot_lo[7:0], data_rot_lo[7:0], data_rot_lo[7:0], data_rot_lo[7:0] }),
    .sel_i(size_i),
    .data_o(data_o)
  );


endmodule



module bp_me_cache_controller_00
(
  clk_i,
  reset_i,
  mem_fwd_header_i,
  mem_fwd_data_i,
  mem_fwd_v_i,
  mem_fwd_ready_and_o,
  mem_rev_header_o,
  mem_rev_data_o,
  mem_rev_v_o,
  mem_rev_ready_and_i,
  cache_pkt_o,
  cache_pkt_v_o,
  cache_pkt_yumi_i,
  cache_data_i,
  cache_data_v_i,
  cache_data_yumi_o
);

  input [64:0] mem_fwd_header_i;
  input [127:0] mem_fwd_data_i;
  output [64:0] mem_rev_header_o;
  output [127:0] mem_rev_data_o;
  output [365:0] cache_pkt_o;
  output [1:0] cache_pkt_v_o;
  input [1:0] cache_pkt_yumi_i;
  input [255:0] cache_data_i;
  input [1:0] cache_data_v_i;
  output [1:0] cache_data_yumi_o;
  input clk_i;
  input reset_i;
  input mem_fwd_v_i;
  input mem_rev_ready_and_i;
  output mem_fwd_ready_and_o;
  output mem_rev_v_o;
  wire [64:0] mem_rev_header_o,fsm_fwd_header_li;
  wire [127:0] mem_rev_data_o,fsm_fwd_data_li,fsm_rev_data_lo,fwd_pkt_data_lo,cache_data_li;
  wire [365:0] cache_pkt_o;
  wire [1:0] cache_pkt_v_o,cache_data_yumi_o,op_data_lo,op_v_lo,
  \cache_pkt_sel_3_.non_max_size.decoded_slice_index ;
  wire mem_fwd_ready_and_o,mem_rev_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,
  N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,
  N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,cache_pkt_o_1__182_,cache_pkt_o_1__181_,
  cache_pkt_o_1__180_,cache_pkt_o_1__179_,cache_pkt_o_1__178_,cache_pkt_o_1__177_,
  cache_pkt_o_1__176_,cache_pkt_o_1__175_,cache_pkt_o_1__174_,cache_pkt_o_1__173_,
  cache_pkt_o_1__172_,cache_pkt_o_1__171_,cache_pkt_o_1__170_,cache_pkt_o_1__169_,
  cache_pkt_o_1__168_,cache_pkt_o_1__167_,cache_pkt_o_1__166_,cache_pkt_o_1__165_,
  cache_pkt_o_1__164_,cache_pkt_o_1__163_,cache_pkt_o_1__162_,cache_pkt_o_1__161_,
  cache_pkt_o_1__160_,cache_pkt_o_1__159_,cache_pkt_o_1__158_,cache_pkt_o_1__157_,
  cache_pkt_o_1__156_,cache_pkt_o_1__155_,cache_pkt_o_1__154_,cache_pkt_o_1__153_,
  cache_pkt_o_1__152_,cache_pkt_o_1__151_,cache_pkt_o_1__150_,cache_pkt_o_1__149_,
  cache_pkt_o_1__148_,cache_pkt_o_1__147_,cache_pkt_o_1__146_,cache_pkt_o_1__145_,
  cache_pkt_o_1__144_,cache_pkt_o_1__143_,cache_pkt_o_1__142_,cache_pkt_o_1__141_,
  cache_pkt_o_1__140_,cache_pkt_o_1__139_,cache_pkt_o_1__138_,cache_pkt_o_1__137_,
  cache_pkt_o_1__136_,cache_pkt_o_1__135_,cache_pkt_o_1__134_,cache_pkt_o_1__133_,
  cache_pkt_o_1__132_,cache_pkt_o_1__131_,cache_pkt_o_1__130_,cache_pkt_o_1__129_,
  cache_pkt_o_1__128_,cache_pkt_o_1__127_,cache_pkt_o_1__126_,cache_pkt_o_1__125_,
  cache_pkt_o_1__124_,cache_pkt_o_1__123_,cache_pkt_o_1__122_,cache_pkt_o_1__121_,
  cache_pkt_o_1__120_,cache_pkt_o_1__119_,cache_pkt_o_1__118_,cache_pkt_o_1__117_,
  cache_pkt_o_1__116_,cache_pkt_o_1__115_,cache_pkt_o_1__114_,cache_pkt_o_1__113_,
  cache_pkt_o_1__112_,cache_pkt_o_1__111_,cache_pkt_o_1__110_,cache_pkt_o_1__109_,
  cache_pkt_o_1__108_,cache_pkt_o_1__107_,cache_pkt_o_1__106_,cache_pkt_o_1__105_,
  cache_pkt_o_1__104_,cache_pkt_o_1__103_,cache_pkt_o_1__102_,cache_pkt_o_1__101_,
  cache_pkt_o_1__100_,cache_pkt_o_1__99_,cache_pkt_o_1__98_,cache_pkt_o_1__97_,cache_pkt_o_1__96_,
  cache_pkt_o_1__95_,cache_pkt_o_1__94_,cache_pkt_o_1__93_,cache_pkt_o_1__92_,
  cache_pkt_o_1__91_,cache_pkt_o_1__90_,cache_pkt_o_1__89_,cache_pkt_o_1__88_,
  cache_pkt_o_1__87_,cache_pkt_o_1__86_,cache_pkt_o_1__85_,cache_pkt_o_1__84_,
  cache_pkt_o_1__83_,cache_pkt_o_1__82_,cache_pkt_o_1__81_,cache_pkt_o_1__80_,
  cache_pkt_o_1__79_,cache_pkt_o_1__78_,cache_pkt_o_1__77_,cache_pkt_o_1__76_,cache_pkt_o_1__75_,
  cache_pkt_o_1__74_,cache_pkt_o_1__73_,cache_pkt_o_1__72_,cache_pkt_o_1__71_,
  cache_pkt_o_1__70_,cache_pkt_o_1__69_,cache_pkt_o_1__68_,cache_pkt_o_1__67_,
  cache_pkt_o_1__66_,cache_pkt_o_1__65_,cache_pkt_o_1__64_,cache_pkt_o_1__63_,
  cache_pkt_o_1__62_,cache_pkt_o_1__61_,cache_pkt_o_1__60_,cache_pkt_o_1__59_,cache_pkt_o_1__58_,
  cache_pkt_o_1__57_,cache_pkt_o_1__56_,cache_pkt_o_1__55_,cache_pkt_o_1__54_,
  cache_pkt_o_1__53_,cache_pkt_o_1__52_,cache_pkt_o_1__51_,cache_pkt_o_1__50_,
  cache_pkt_o_1__49_,cache_pkt_o_1__48_,cache_pkt_o_1__47_,cache_pkt_o_1__46_,
  cache_pkt_o_1__45_,cache_pkt_o_1__44_,cache_pkt_o_1__43_,cache_pkt_o_1__42_,
  cache_pkt_o_1__41_,cache_pkt_o_1__40_,cache_pkt_o_1__39_,cache_pkt_o_1__38_,cache_pkt_o_1__37_,
  cache_pkt_o_1__36_,cache_pkt_o_1__35_,cache_pkt_o_1__34_,cache_pkt_o_1__33_,
  cache_pkt_o_1__32_,cache_pkt_o_1__31_,cache_pkt_o_1__30_,cache_pkt_o_1__29_,
  cache_pkt_o_1__28_,cache_pkt_o_1__27_,cache_pkt_o_1__26_,cache_pkt_o_1__25_,
  cache_pkt_o_1__24_,cache_pkt_o_1__23_,cache_pkt_o_1__22_,cache_pkt_o_1__21_,
  cache_pkt_o_1__20_,cache_pkt_o_1__19_,cache_pkt_o_1__18_,cache_pkt_o_1__17_,cache_pkt_o_1__16_,
  cache_pkt_o_1__15_,cache_pkt_o_1__14_,cache_pkt_o_1__13_,cache_pkt_o_1__12_,
  cache_pkt_o_1__11_,cache_pkt_o_1__10_,cache_pkt_o_1__9_,cache_pkt_o_1__8_,
  cache_pkt_o_1__7_,cache_pkt_o_1__6_,cache_pkt_o_1__5_,cache_pkt_o_1__4_,cache_pkt_o_1__3_,
  cache_pkt_o_1__2_,cache_pkt_o_1__1_,cache_pkt_o_1__0_,fsm_fwd_v_li,
  fsm_fwd_yumi_lo,fsm_fwd_new_li,fsm_fwd_critical_li,fsm_fwd_last_li,fsm_rev_v_lo,
  fsm_rev_ready_then_li,fsm_rev_new_lo,fsm_rev_critical_lo,fsm_rev_last_lo,N60,N61,is_uc_op,
  set_clear,set_up,cache_pkt_mask_mux_li_3__15_,cache_pkt_mask_mux_li_3__14_,
  cache_pkt_mask_mux_li_3__13_,cache_pkt_mask_mux_li_3__12_,cache_pkt_mask_mux_li_3__11_,
  cache_pkt_mask_mux_li_3__10_,cache_pkt_mask_mux_li_3__9_,
  cache_pkt_mask_mux_li_3__8_,cache_pkt_mask_mux_li_3__7_,cache_pkt_mask_mux_li_3__6_,
  cache_pkt_mask_mux_li_3__5_,cache_pkt_mask_mux_li_3__4_,cache_pkt_mask_mux_li_3__3_,
  cache_pkt_mask_mux_li_3__2_,cache_pkt_mask_mux_li_3__1_,cache_pkt_mask_mux_li_3__0_,
  cache_pkt_mask_mux_li_2__15_,cache_pkt_mask_mux_li_2__14_,cache_pkt_mask_mux_li_2__13_,
  cache_pkt_mask_mux_li_2__12_,cache_pkt_mask_mux_li_2__11_,cache_pkt_mask_mux_li_2__10_,
  cache_pkt_mask_mux_li_2__9_,cache_pkt_mask_mux_li_2__8_,
  cache_pkt_mask_mux_li_2__7_,cache_pkt_mask_mux_li_2__6_,cache_pkt_mask_mux_li_2__5_,
  cache_pkt_mask_mux_li_2__4_,cache_pkt_mask_mux_li_2__3_,cache_pkt_mask_mux_li_2__2_,
  cache_pkt_mask_mux_li_2__1_,cache_pkt_mask_mux_li_2__0_,cache_pkt_mask_mux_li_1__15_,
  cache_pkt_mask_mux_li_1__14_,cache_pkt_mask_mux_li_1__13_,cache_pkt_mask_mux_li_1__12_,
  cache_pkt_mask_mux_li_1__11_,cache_pkt_mask_mux_li_1__10_,
  cache_pkt_mask_mux_li_1__9_,cache_pkt_mask_mux_li_1__8_,cache_pkt_mask_mux_li_1__7_,
  cache_pkt_mask_mux_li_1__6_,cache_pkt_mask_mux_li_1__5_,cache_pkt_mask_mux_li_1__4_,
  cache_pkt_mask_mux_li_1__3_,cache_pkt_mask_mux_li_1__2_,cache_pkt_mask_mux_li_1__1_,
  cache_pkt_mask_mux_li_1__0_,cache_pkt_mask_mux_li_0__15_,cache_pkt_mask_mux_li_0__14_,
  cache_pkt_mask_mux_li_0__13_,cache_pkt_mask_mux_li_0__12_,cache_pkt_mask_mux_li_0__11_,
  cache_pkt_mask_mux_li_0__10_,cache_pkt_mask_mux_li_0__9_,
  cache_pkt_mask_mux_li_0__8_,cache_pkt_mask_mux_li_0__7_,cache_pkt_mask_mux_li_0__6_,
  cache_pkt_mask_mux_li_0__5_,cache_pkt_mask_mux_li_0__4_,cache_pkt_mask_mux_li_0__3_,
  cache_pkt_mask_mux_li_0__2_,cache_pkt_mask_mux_li_0__1_,cache_pkt_mask_mux_li_0__0_,N62,N63,N64,
  N65,N66,N67,N68,N69,N70,N71,fwd_pkt_dram_lo,cache_pkt_v_lo,N72,N73,
  cache_pkt_yumi_li,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,
  N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,
  N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,
  N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,
  N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,
  N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,
  N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,
  N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,
  N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,
  N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,
  N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,
  N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
  N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,
  N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,
  N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,
  N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,
  N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,
  N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,
  N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,
  N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,
  N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,
  N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,
  N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,
  N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,
  N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,
  sv2v_dc_1;
  wire [2:0] state_r,cache_pkt_sel_li,fsm_rev_size_li,state_n;
  wire [39:0] fsm_fwd_addr_li,fsm_rev_addr_lo;
  wire [65:0] fsm_rev_metadata_lo;
  wire [10:0] set_cnt;
  wire [15:0] \cache_pkt_sel_0_.non_max_size.decoded_slice_index ,cache_pkt_mask_lo;
  wire [7:0] \cache_pkt_sel_1_.non_max_size.decoded_slice_index ;
  wire [3:0] \cache_pkt_sel_2_.non_max_size.decoded_slice_index ;
  wire [32:0] fwd_pkt_daddr_lo;
  wire [0:0] fwd_pkt_bank_lo,cache_fwd_bank_lo;
  reg state_r_2_sv2v_reg,state_r_1_sv2v_reg,state_r_0_sv2v_reg;
  assign state_r[2] = state_r_2_sv2v_reg;
  assign state_r[1] = state_r_1_sv2v_reg;
  assign state_r[0] = state_r_0_sv2v_reg;
  assign cache_pkt_o[182] = cache_pkt_o_1__182_;
  assign cache_pkt_o[365] = cache_pkt_o_1__182_;
  assign cache_pkt_o[181] = cache_pkt_o_1__181_;
  assign cache_pkt_o[364] = cache_pkt_o_1__181_;
  assign cache_pkt_o[180] = cache_pkt_o_1__180_;
  assign cache_pkt_o[363] = cache_pkt_o_1__180_;
  assign cache_pkt_o[179] = cache_pkt_o_1__179_;
  assign cache_pkt_o[362] = cache_pkt_o_1__179_;
  assign cache_pkt_o[178] = cache_pkt_o_1__178_;
  assign cache_pkt_o[361] = cache_pkt_o_1__178_;
  assign cache_pkt_o[177] = cache_pkt_o_1__177_;
  assign cache_pkt_o[360] = cache_pkt_o_1__177_;
  assign cache_pkt_o[176] = cache_pkt_o_1__176_;
  assign cache_pkt_o[359] = cache_pkt_o_1__176_;
  assign cache_pkt_o[175] = cache_pkt_o_1__175_;
  assign cache_pkt_o[358] = cache_pkt_o_1__175_;
  assign cache_pkt_o[174] = cache_pkt_o_1__174_;
  assign cache_pkt_o[357] = cache_pkt_o_1__174_;
  assign cache_pkt_o[173] = cache_pkt_o_1__173_;
  assign cache_pkt_o[356] = cache_pkt_o_1__173_;
  assign cache_pkt_o[172] = cache_pkt_o_1__172_;
  assign cache_pkt_o[355] = cache_pkt_o_1__172_;
  assign cache_pkt_o[171] = cache_pkt_o_1__171_;
  assign cache_pkt_o[354] = cache_pkt_o_1__171_;
  assign cache_pkt_o[170] = cache_pkt_o_1__170_;
  assign cache_pkt_o[353] = cache_pkt_o_1__170_;
  assign cache_pkt_o[169] = cache_pkt_o_1__169_;
  assign cache_pkt_o[352] = cache_pkt_o_1__169_;
  assign cache_pkt_o[168] = cache_pkt_o_1__168_;
  assign cache_pkt_o[351] = cache_pkt_o_1__168_;
  assign cache_pkt_o[167] = cache_pkt_o_1__167_;
  assign cache_pkt_o[350] = cache_pkt_o_1__167_;
  assign cache_pkt_o[166] = cache_pkt_o_1__166_;
  assign cache_pkt_o[349] = cache_pkt_o_1__166_;
  assign cache_pkt_o[165] = cache_pkt_o_1__165_;
  assign cache_pkt_o[348] = cache_pkt_o_1__165_;
  assign cache_pkt_o[164] = cache_pkt_o_1__164_;
  assign cache_pkt_o[347] = cache_pkt_o_1__164_;
  assign cache_pkt_o[163] = cache_pkt_o_1__163_;
  assign cache_pkt_o[346] = cache_pkt_o_1__163_;
  assign cache_pkt_o[162] = cache_pkt_o_1__162_;
  assign cache_pkt_o[345] = cache_pkt_o_1__162_;
  assign cache_pkt_o[161] = cache_pkt_o_1__161_;
  assign cache_pkt_o[344] = cache_pkt_o_1__161_;
  assign cache_pkt_o[160] = cache_pkt_o_1__160_;
  assign cache_pkt_o[343] = cache_pkt_o_1__160_;
  assign cache_pkt_o[159] = cache_pkt_o_1__159_;
  assign cache_pkt_o[342] = cache_pkt_o_1__159_;
  assign cache_pkt_o[158] = cache_pkt_o_1__158_;
  assign cache_pkt_o[341] = cache_pkt_o_1__158_;
  assign cache_pkt_o[157] = cache_pkt_o_1__157_;
  assign cache_pkt_o[340] = cache_pkt_o_1__157_;
  assign cache_pkt_o[156] = cache_pkt_o_1__156_;
  assign cache_pkt_o[339] = cache_pkt_o_1__156_;
  assign cache_pkt_o[155] = cache_pkt_o_1__155_;
  assign cache_pkt_o[338] = cache_pkt_o_1__155_;
  assign cache_pkt_o[154] = cache_pkt_o_1__154_;
  assign cache_pkt_o[337] = cache_pkt_o_1__154_;
  assign cache_pkt_o[153] = cache_pkt_o_1__153_;
  assign cache_pkt_o[336] = cache_pkt_o_1__153_;
  assign cache_pkt_o[152] = cache_pkt_o_1__152_;
  assign cache_pkt_o[335] = cache_pkt_o_1__152_;
  assign cache_pkt_o[151] = cache_pkt_o_1__151_;
  assign cache_pkt_o[334] = cache_pkt_o_1__151_;
  assign cache_pkt_o[150] = cache_pkt_o_1__150_;
  assign cache_pkt_o[333] = cache_pkt_o_1__150_;
  assign cache_pkt_o[149] = cache_pkt_o_1__149_;
  assign cache_pkt_o[332] = cache_pkt_o_1__149_;
  assign cache_pkt_o[148] = cache_pkt_o_1__148_;
  assign cache_pkt_o[331] = cache_pkt_o_1__148_;
  assign cache_pkt_o[147] = cache_pkt_o_1__147_;
  assign cache_pkt_o[330] = cache_pkt_o_1__147_;
  assign cache_pkt_o[146] = cache_pkt_o_1__146_;
  assign cache_pkt_o[329] = cache_pkt_o_1__146_;
  assign cache_pkt_o[145] = cache_pkt_o_1__145_;
  assign cache_pkt_o[328] = cache_pkt_o_1__145_;
  assign cache_pkt_o[144] = cache_pkt_o_1__144_;
  assign cache_pkt_o[327] = cache_pkt_o_1__144_;
  assign cache_pkt_o[143] = cache_pkt_o_1__143_;
  assign cache_pkt_o[326] = cache_pkt_o_1__143_;
  assign cache_pkt_o[142] = cache_pkt_o_1__142_;
  assign cache_pkt_o[325] = cache_pkt_o_1__142_;
  assign cache_pkt_o[141] = cache_pkt_o_1__141_;
  assign cache_pkt_o[324] = cache_pkt_o_1__141_;
  assign cache_pkt_o[140] = cache_pkt_o_1__140_;
  assign cache_pkt_o[323] = cache_pkt_o_1__140_;
  assign cache_pkt_o[139] = cache_pkt_o_1__139_;
  assign cache_pkt_o[322] = cache_pkt_o_1__139_;
  assign cache_pkt_o[138] = cache_pkt_o_1__138_;
  assign cache_pkt_o[321] = cache_pkt_o_1__138_;
  assign cache_pkt_o[137] = cache_pkt_o_1__137_;
  assign cache_pkt_o[320] = cache_pkt_o_1__137_;
  assign cache_pkt_o[136] = cache_pkt_o_1__136_;
  assign cache_pkt_o[319] = cache_pkt_o_1__136_;
  assign cache_pkt_o[135] = cache_pkt_o_1__135_;
  assign cache_pkt_o[318] = cache_pkt_o_1__135_;
  assign cache_pkt_o[134] = cache_pkt_o_1__134_;
  assign cache_pkt_o[317] = cache_pkt_o_1__134_;
  assign cache_pkt_o[133] = cache_pkt_o_1__133_;
  assign cache_pkt_o[316] = cache_pkt_o_1__133_;
  assign cache_pkt_o[132] = cache_pkt_o_1__132_;
  assign cache_pkt_o[315] = cache_pkt_o_1__132_;
  assign cache_pkt_o[131] = cache_pkt_o_1__131_;
  assign cache_pkt_o[314] = cache_pkt_o_1__131_;
  assign cache_pkt_o[130] = cache_pkt_o_1__130_;
  assign cache_pkt_o[313] = cache_pkt_o_1__130_;
  assign cache_pkt_o[129] = cache_pkt_o_1__129_;
  assign cache_pkt_o[312] = cache_pkt_o_1__129_;
  assign cache_pkt_o[128] = cache_pkt_o_1__128_;
  assign cache_pkt_o[311] = cache_pkt_o_1__128_;
  assign cache_pkt_o[127] = cache_pkt_o_1__127_;
  assign cache_pkt_o[310] = cache_pkt_o_1__127_;
  assign cache_pkt_o[126] = cache_pkt_o_1__126_;
  assign cache_pkt_o[309] = cache_pkt_o_1__126_;
  assign cache_pkt_o[125] = cache_pkt_o_1__125_;
  assign cache_pkt_o[308] = cache_pkt_o_1__125_;
  assign cache_pkt_o[124] = cache_pkt_o_1__124_;
  assign cache_pkt_o[307] = cache_pkt_o_1__124_;
  assign cache_pkt_o[123] = cache_pkt_o_1__123_;
  assign cache_pkt_o[306] = cache_pkt_o_1__123_;
  assign cache_pkt_o[122] = cache_pkt_o_1__122_;
  assign cache_pkt_o[305] = cache_pkt_o_1__122_;
  assign cache_pkt_o[121] = cache_pkt_o_1__121_;
  assign cache_pkt_o[304] = cache_pkt_o_1__121_;
  assign cache_pkt_o[120] = cache_pkt_o_1__120_;
  assign cache_pkt_o[303] = cache_pkt_o_1__120_;
  assign cache_pkt_o[119] = cache_pkt_o_1__119_;
  assign cache_pkt_o[302] = cache_pkt_o_1__119_;
  assign cache_pkt_o[118] = cache_pkt_o_1__118_;
  assign cache_pkt_o[301] = cache_pkt_o_1__118_;
  assign cache_pkt_o[117] = cache_pkt_o_1__117_;
  assign cache_pkt_o[300] = cache_pkt_o_1__117_;
  assign cache_pkt_o[116] = cache_pkt_o_1__116_;
  assign cache_pkt_o[299] = cache_pkt_o_1__116_;
  assign cache_pkt_o[115] = cache_pkt_o_1__115_;
  assign cache_pkt_o[298] = cache_pkt_o_1__115_;
  assign cache_pkt_o[114] = cache_pkt_o_1__114_;
  assign cache_pkt_o[297] = cache_pkt_o_1__114_;
  assign cache_pkt_o[113] = cache_pkt_o_1__113_;
  assign cache_pkt_o[296] = cache_pkt_o_1__113_;
  assign cache_pkt_o[112] = cache_pkt_o_1__112_;
  assign cache_pkt_o[295] = cache_pkt_o_1__112_;
  assign cache_pkt_o[111] = cache_pkt_o_1__111_;
  assign cache_pkt_o[294] = cache_pkt_o_1__111_;
  assign cache_pkt_o[110] = cache_pkt_o_1__110_;
  assign cache_pkt_o[293] = cache_pkt_o_1__110_;
  assign cache_pkt_o[109] = cache_pkt_o_1__109_;
  assign cache_pkt_o[292] = cache_pkt_o_1__109_;
  assign cache_pkt_o[108] = cache_pkt_o_1__108_;
  assign cache_pkt_o[291] = cache_pkt_o_1__108_;
  assign cache_pkt_o[107] = cache_pkt_o_1__107_;
  assign cache_pkt_o[290] = cache_pkt_o_1__107_;
  assign cache_pkt_o[106] = cache_pkt_o_1__106_;
  assign cache_pkt_o[289] = cache_pkt_o_1__106_;
  assign cache_pkt_o[105] = cache_pkt_o_1__105_;
  assign cache_pkt_o[288] = cache_pkt_o_1__105_;
  assign cache_pkt_o[104] = cache_pkt_o_1__104_;
  assign cache_pkt_o[287] = cache_pkt_o_1__104_;
  assign cache_pkt_o[103] = cache_pkt_o_1__103_;
  assign cache_pkt_o[286] = cache_pkt_o_1__103_;
  assign cache_pkt_o[102] = cache_pkt_o_1__102_;
  assign cache_pkt_o[285] = cache_pkt_o_1__102_;
  assign cache_pkt_o[101] = cache_pkt_o_1__101_;
  assign cache_pkt_o[284] = cache_pkt_o_1__101_;
  assign cache_pkt_o[100] = cache_pkt_o_1__100_;
  assign cache_pkt_o[283] = cache_pkt_o_1__100_;
  assign cache_pkt_o[99] = cache_pkt_o_1__99_;
  assign cache_pkt_o[282] = cache_pkt_o_1__99_;
  assign cache_pkt_o[98] = cache_pkt_o_1__98_;
  assign cache_pkt_o[281] = cache_pkt_o_1__98_;
  assign cache_pkt_o[97] = cache_pkt_o_1__97_;
  assign cache_pkt_o[280] = cache_pkt_o_1__97_;
  assign cache_pkt_o[96] = cache_pkt_o_1__96_;
  assign cache_pkt_o[279] = cache_pkt_o_1__96_;
  assign cache_pkt_o[95] = cache_pkt_o_1__95_;
  assign cache_pkt_o[278] = cache_pkt_o_1__95_;
  assign cache_pkt_o[94] = cache_pkt_o_1__94_;
  assign cache_pkt_o[277] = cache_pkt_o_1__94_;
  assign cache_pkt_o[93] = cache_pkt_o_1__93_;
  assign cache_pkt_o[276] = cache_pkt_o_1__93_;
  assign cache_pkt_o[92] = cache_pkt_o_1__92_;
  assign cache_pkt_o[275] = cache_pkt_o_1__92_;
  assign cache_pkt_o[91] = cache_pkt_o_1__91_;
  assign cache_pkt_o[274] = cache_pkt_o_1__91_;
  assign cache_pkt_o[90] = cache_pkt_o_1__90_;
  assign cache_pkt_o[273] = cache_pkt_o_1__90_;
  assign cache_pkt_o[89] = cache_pkt_o_1__89_;
  assign cache_pkt_o[272] = cache_pkt_o_1__89_;
  assign cache_pkt_o[88] = cache_pkt_o_1__88_;
  assign cache_pkt_o[271] = cache_pkt_o_1__88_;
  assign cache_pkt_o[87] = cache_pkt_o_1__87_;
  assign cache_pkt_o[270] = cache_pkt_o_1__87_;
  assign cache_pkt_o[86] = cache_pkt_o_1__86_;
  assign cache_pkt_o[269] = cache_pkt_o_1__86_;
  assign cache_pkt_o[85] = cache_pkt_o_1__85_;
  assign cache_pkt_o[268] = cache_pkt_o_1__85_;
  assign cache_pkt_o[84] = cache_pkt_o_1__84_;
  assign cache_pkt_o[267] = cache_pkt_o_1__84_;
  assign cache_pkt_o[83] = cache_pkt_o_1__83_;
  assign cache_pkt_o[266] = cache_pkt_o_1__83_;
  assign cache_pkt_o[82] = cache_pkt_o_1__82_;
  assign cache_pkt_o[265] = cache_pkt_o_1__82_;
  assign cache_pkt_o[81] = cache_pkt_o_1__81_;
  assign cache_pkt_o[264] = cache_pkt_o_1__81_;
  assign cache_pkt_o[80] = cache_pkt_o_1__80_;
  assign cache_pkt_o[263] = cache_pkt_o_1__80_;
  assign cache_pkt_o[79] = cache_pkt_o_1__79_;
  assign cache_pkt_o[262] = cache_pkt_o_1__79_;
  assign cache_pkt_o[78] = cache_pkt_o_1__78_;
  assign cache_pkt_o[261] = cache_pkt_o_1__78_;
  assign cache_pkt_o[77] = cache_pkt_o_1__77_;
  assign cache_pkt_o[260] = cache_pkt_o_1__77_;
  assign cache_pkt_o[76] = cache_pkt_o_1__76_;
  assign cache_pkt_o[259] = cache_pkt_o_1__76_;
  assign cache_pkt_o[75] = cache_pkt_o_1__75_;
  assign cache_pkt_o[258] = cache_pkt_o_1__75_;
  assign cache_pkt_o[74] = cache_pkt_o_1__74_;
  assign cache_pkt_o[257] = cache_pkt_o_1__74_;
  assign cache_pkt_o[73] = cache_pkt_o_1__73_;
  assign cache_pkt_o[256] = cache_pkt_o_1__73_;
  assign cache_pkt_o[72] = cache_pkt_o_1__72_;
  assign cache_pkt_o[255] = cache_pkt_o_1__72_;
  assign cache_pkt_o[71] = cache_pkt_o_1__71_;
  assign cache_pkt_o[254] = cache_pkt_o_1__71_;
  assign cache_pkt_o[70] = cache_pkt_o_1__70_;
  assign cache_pkt_o[253] = cache_pkt_o_1__70_;
  assign cache_pkt_o[69] = cache_pkt_o_1__69_;
  assign cache_pkt_o[252] = cache_pkt_o_1__69_;
  assign cache_pkt_o[68] = cache_pkt_o_1__68_;
  assign cache_pkt_o[251] = cache_pkt_o_1__68_;
  assign cache_pkt_o[67] = cache_pkt_o_1__67_;
  assign cache_pkt_o[250] = cache_pkt_o_1__67_;
  assign cache_pkt_o[66] = cache_pkt_o_1__66_;
  assign cache_pkt_o[249] = cache_pkt_o_1__66_;
  assign cache_pkt_o[65] = cache_pkt_o_1__65_;
  assign cache_pkt_o[248] = cache_pkt_o_1__65_;
  assign cache_pkt_o[64] = cache_pkt_o_1__64_;
  assign cache_pkt_o[247] = cache_pkt_o_1__64_;
  assign cache_pkt_o[63] = cache_pkt_o_1__63_;
  assign cache_pkt_o[246] = cache_pkt_o_1__63_;
  assign cache_pkt_o[62] = cache_pkt_o_1__62_;
  assign cache_pkt_o[245] = cache_pkt_o_1__62_;
  assign cache_pkt_o[61] = cache_pkt_o_1__61_;
  assign cache_pkt_o[244] = cache_pkt_o_1__61_;
  assign cache_pkt_o[60] = cache_pkt_o_1__60_;
  assign cache_pkt_o[243] = cache_pkt_o_1__60_;
  assign cache_pkt_o[59] = cache_pkt_o_1__59_;
  assign cache_pkt_o[242] = cache_pkt_o_1__59_;
  assign cache_pkt_o[58] = cache_pkt_o_1__58_;
  assign cache_pkt_o[241] = cache_pkt_o_1__58_;
  assign cache_pkt_o[57] = cache_pkt_o_1__57_;
  assign cache_pkt_o[240] = cache_pkt_o_1__57_;
  assign cache_pkt_o[56] = cache_pkt_o_1__56_;
  assign cache_pkt_o[239] = cache_pkt_o_1__56_;
  assign cache_pkt_o[55] = cache_pkt_o_1__55_;
  assign cache_pkt_o[238] = cache_pkt_o_1__55_;
  assign cache_pkt_o[54] = cache_pkt_o_1__54_;
  assign cache_pkt_o[237] = cache_pkt_o_1__54_;
  assign cache_pkt_o[53] = cache_pkt_o_1__53_;
  assign cache_pkt_o[236] = cache_pkt_o_1__53_;
  assign cache_pkt_o[52] = cache_pkt_o_1__52_;
  assign cache_pkt_o[235] = cache_pkt_o_1__52_;
  assign cache_pkt_o[51] = cache_pkt_o_1__51_;
  assign cache_pkt_o[234] = cache_pkt_o_1__51_;
  assign cache_pkt_o[50] = cache_pkt_o_1__50_;
  assign cache_pkt_o[233] = cache_pkt_o_1__50_;
  assign cache_pkt_o[49] = cache_pkt_o_1__49_;
  assign cache_pkt_o[232] = cache_pkt_o_1__49_;
  assign cache_pkt_o[48] = cache_pkt_o_1__48_;
  assign cache_pkt_o[231] = cache_pkt_o_1__48_;
  assign cache_pkt_o[47] = cache_pkt_o_1__47_;
  assign cache_pkt_o[230] = cache_pkt_o_1__47_;
  assign cache_pkt_o[46] = cache_pkt_o_1__46_;
  assign cache_pkt_o[229] = cache_pkt_o_1__46_;
  assign cache_pkt_o[45] = cache_pkt_o_1__45_;
  assign cache_pkt_o[228] = cache_pkt_o_1__45_;
  assign cache_pkt_o[44] = cache_pkt_o_1__44_;
  assign cache_pkt_o[227] = cache_pkt_o_1__44_;
  assign cache_pkt_o[43] = cache_pkt_o_1__43_;
  assign cache_pkt_o[226] = cache_pkt_o_1__43_;
  assign cache_pkt_o[42] = cache_pkt_o_1__42_;
  assign cache_pkt_o[225] = cache_pkt_o_1__42_;
  assign cache_pkt_o[41] = cache_pkt_o_1__41_;
  assign cache_pkt_o[224] = cache_pkt_o_1__41_;
  assign cache_pkt_o[40] = cache_pkt_o_1__40_;
  assign cache_pkt_o[223] = cache_pkt_o_1__40_;
  assign cache_pkt_o[39] = cache_pkt_o_1__39_;
  assign cache_pkt_o[222] = cache_pkt_o_1__39_;
  assign cache_pkt_o[38] = cache_pkt_o_1__38_;
  assign cache_pkt_o[221] = cache_pkt_o_1__38_;
  assign cache_pkt_o[37] = cache_pkt_o_1__37_;
  assign cache_pkt_o[220] = cache_pkt_o_1__37_;
  assign cache_pkt_o[36] = cache_pkt_o_1__36_;
  assign cache_pkt_o[219] = cache_pkt_o_1__36_;
  assign cache_pkt_o[35] = cache_pkt_o_1__35_;
  assign cache_pkt_o[218] = cache_pkt_o_1__35_;
  assign cache_pkt_o[34] = cache_pkt_o_1__34_;
  assign cache_pkt_o[217] = cache_pkt_o_1__34_;
  assign cache_pkt_o[33] = cache_pkt_o_1__33_;
  assign cache_pkt_o[216] = cache_pkt_o_1__33_;
  assign cache_pkt_o[32] = cache_pkt_o_1__32_;
  assign cache_pkt_o[215] = cache_pkt_o_1__32_;
  assign cache_pkt_o[31] = cache_pkt_o_1__31_;
  assign cache_pkt_o[214] = cache_pkt_o_1__31_;
  assign cache_pkt_o[30] = cache_pkt_o_1__30_;
  assign cache_pkt_o[213] = cache_pkt_o_1__30_;
  assign cache_pkt_o[29] = cache_pkt_o_1__29_;
  assign cache_pkt_o[212] = cache_pkt_o_1__29_;
  assign cache_pkt_o[28] = cache_pkt_o_1__28_;
  assign cache_pkt_o[211] = cache_pkt_o_1__28_;
  assign cache_pkt_o[27] = cache_pkt_o_1__27_;
  assign cache_pkt_o[210] = cache_pkt_o_1__27_;
  assign cache_pkt_o[26] = cache_pkt_o_1__26_;
  assign cache_pkt_o[209] = cache_pkt_o_1__26_;
  assign cache_pkt_o[25] = cache_pkt_o_1__25_;
  assign cache_pkt_o[208] = cache_pkt_o_1__25_;
  assign cache_pkt_o[24] = cache_pkt_o_1__24_;
  assign cache_pkt_o[207] = cache_pkt_o_1__24_;
  assign cache_pkt_o[23] = cache_pkt_o_1__23_;
  assign cache_pkt_o[206] = cache_pkt_o_1__23_;
  assign cache_pkt_o[22] = cache_pkt_o_1__22_;
  assign cache_pkt_o[205] = cache_pkt_o_1__22_;
  assign cache_pkt_o[21] = cache_pkt_o_1__21_;
  assign cache_pkt_o[204] = cache_pkt_o_1__21_;
  assign cache_pkt_o[20] = cache_pkt_o_1__20_;
  assign cache_pkt_o[203] = cache_pkt_o_1__20_;
  assign cache_pkt_o[19] = cache_pkt_o_1__19_;
  assign cache_pkt_o[202] = cache_pkt_o_1__19_;
  assign cache_pkt_o[18] = cache_pkt_o_1__18_;
  assign cache_pkt_o[201] = cache_pkt_o_1__18_;
  assign cache_pkt_o[17] = cache_pkt_o_1__17_;
  assign cache_pkt_o[200] = cache_pkt_o_1__17_;
  assign cache_pkt_o[16] = cache_pkt_o_1__16_;
  assign cache_pkt_o[199] = cache_pkt_o_1__16_;
  assign cache_pkt_o[15] = cache_pkt_o_1__15_;
  assign cache_pkt_o[198] = cache_pkt_o_1__15_;
  assign cache_pkt_o[14] = cache_pkt_o_1__14_;
  assign cache_pkt_o[197] = cache_pkt_o_1__14_;
  assign cache_pkt_o[13] = cache_pkt_o_1__13_;
  assign cache_pkt_o[196] = cache_pkt_o_1__13_;
  assign cache_pkt_o[12] = cache_pkt_o_1__12_;
  assign cache_pkt_o[195] = cache_pkt_o_1__12_;
  assign cache_pkt_o[11] = cache_pkt_o_1__11_;
  assign cache_pkt_o[194] = cache_pkt_o_1__11_;
  assign cache_pkt_o[10] = cache_pkt_o_1__10_;
  assign cache_pkt_o[193] = cache_pkt_o_1__10_;
  assign cache_pkt_o[9] = cache_pkt_o_1__9_;
  assign cache_pkt_o[192] = cache_pkt_o_1__9_;
  assign cache_pkt_o[8] = cache_pkt_o_1__8_;
  assign cache_pkt_o[191] = cache_pkt_o_1__8_;
  assign cache_pkt_o[7] = cache_pkt_o_1__7_;
  assign cache_pkt_o[190] = cache_pkt_o_1__7_;
  assign cache_pkt_o[6] = cache_pkt_o_1__6_;
  assign cache_pkt_o[189] = cache_pkt_o_1__6_;
  assign cache_pkt_o[5] = cache_pkt_o_1__5_;
  assign cache_pkt_o[188] = cache_pkt_o_1__5_;
  assign cache_pkt_o[4] = cache_pkt_o_1__4_;
  assign cache_pkt_o[187] = cache_pkt_o_1__4_;
  assign cache_pkt_o[3] = cache_pkt_o_1__3_;
  assign cache_pkt_o[186] = cache_pkt_o_1__3_;
  assign cache_pkt_o[2] = cache_pkt_o_1__2_;
  assign cache_pkt_o[185] = cache_pkt_o_1__2_;
  assign cache_pkt_o[1] = cache_pkt_o_1__1_;
  assign cache_pkt_o[184] = cache_pkt_o_1__1_;
  assign cache_pkt_o[0] = cache_pkt_o_1__0_;
  assign cache_pkt_o[183] = cache_pkt_o_1__0_;

  bsg_fifo_1r1w_small_width_p1_els_p3_ready_THEN_valid_p1
  \tag_0_.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(cache_pkt_yumi_i[0]),
    .data_i(N446),
    .v_o(op_v_lo[0]),
    .data_o(op_data_lo[0]),
    .yumi_i(cache_data_yumi_o[0])
  );


  bsg_fifo_1r1w_small_width_p1_els_p3_ready_THEN_valid_p1
  \tag_1_.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(cache_pkt_yumi_i[1]),
    .data_i(N446),
    .v_o(op_v_lo[1]),
    .data_o(op_data_lo[1]),
    .yumi_i(cache_data_yumi_o[1])
  );


  bp_me_stream_pump_00_00000080_0000000e_6_7_00000080_0000000e_5_7_00000042_00000006
  stream_pump
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .in_msg_header_i(mem_fwd_header_i),
    .in_msg_data_i(mem_fwd_data_i),
    .in_msg_v_i(mem_fwd_v_i),
    .in_msg_ready_and_o(mem_fwd_ready_and_o),
    .in_fsm_header_o(fsm_fwd_header_li),
    .in_fsm_data_o(fsm_fwd_data_li),
    .in_fsm_v_o(fsm_fwd_v_li),
    .in_fsm_yumi_i(fsm_fwd_yumi_lo),
    .in_fsm_metadata_i({ fwd_pkt_bank_lo[0:0], fsm_fwd_header_li }),
    .in_fsm_addr_o(fsm_fwd_addr_li),
    .in_fsm_new_o(fsm_fwd_new_li),
    .in_fsm_critical_o(fsm_fwd_critical_li),
    .in_fsm_last_o(fsm_fwd_last_li),
    .out_msg_header_o(mem_rev_header_o),
    .out_msg_data_o(mem_rev_data_o),
    .out_msg_v_o(mem_rev_v_o),
    .out_msg_ready_and_i(mem_rev_ready_and_i),
    .out_fsm_header_i(fsm_rev_metadata_lo[64:0]),
    .out_fsm_data_i(fsm_rev_data_lo),
    .out_fsm_v_i(fsm_rev_v_lo),
    .out_fsm_ready_then_o(fsm_rev_ready_then_li),
    .out_fsm_metadata_o(fsm_rev_metadata_lo),
    .out_fsm_addr_o(fsm_rev_addr_lo),
    .out_fsm_new_o(fsm_rev_new_lo),
    .out_fsm_last_o(fsm_rev_last_lo),
    .out_fsm_critical_o(fsm_rev_critical_lo)
  );

  assign N60 = fsm_fwd_addr_li >= { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign N61 = fsm_fwd_addr_li < { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };

  bsg_counter_clear_up_000007ff_0
  set_counter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(set_clear),
    .up_i(set_up),
    .count_o(set_cnt)
  );

  assign \cache_pkt_sel_0_.non_max_size.decoded_slice_index  = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fsm_fwd_addr_li[3:0];

  bsg_expand_bitmask_00000010_1
  \cache_pkt_sel_0_.non_max_size.mask_expand 
  (
    .i(\cache_pkt_sel_0_.non_max_size.decoded_slice_index ),
    .o({ cache_pkt_mask_mux_li_0__15_, cache_pkt_mask_mux_li_0__14_, cache_pkt_mask_mux_li_0__13_, cache_pkt_mask_mux_li_0__12_, cache_pkt_mask_mux_li_0__11_, cache_pkt_mask_mux_li_0__10_, cache_pkt_mask_mux_li_0__9_, cache_pkt_mask_mux_li_0__8_, cache_pkt_mask_mux_li_0__7_, cache_pkt_mask_mux_li_0__6_, cache_pkt_mask_mux_li_0__5_, cache_pkt_mask_mux_li_0__4_, cache_pkt_mask_mux_li_0__3_, cache_pkt_mask_mux_li_0__2_, cache_pkt_mask_mux_li_0__1_, cache_pkt_mask_mux_li_0__0_ })
  );

  assign \cache_pkt_sel_1_.non_max_size.decoded_slice_index  = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fsm_fwd_addr_li[3:1];

  bsg_expand_bitmask_00000008_2
  \cache_pkt_sel_1_.non_max_size.mask_expand 
  (
    .i(\cache_pkt_sel_1_.non_max_size.decoded_slice_index ),
    .o({ cache_pkt_mask_mux_li_1__15_, cache_pkt_mask_mux_li_1__14_, cache_pkt_mask_mux_li_1__13_, cache_pkt_mask_mux_li_1__12_, cache_pkt_mask_mux_li_1__11_, cache_pkt_mask_mux_li_1__10_, cache_pkt_mask_mux_li_1__9_, cache_pkt_mask_mux_li_1__8_, cache_pkt_mask_mux_li_1__7_, cache_pkt_mask_mux_li_1__6_, cache_pkt_mask_mux_li_1__5_, cache_pkt_mask_mux_li_1__4_, cache_pkt_mask_mux_li_1__3_, cache_pkt_mask_mux_li_1__2_, cache_pkt_mask_mux_li_1__1_, cache_pkt_mask_mux_li_1__0_ })
  );

  assign \cache_pkt_sel_2_.non_max_size.decoded_slice_index  = { 1'b0, 1'b0, 1'b0, 1'b1 } << fsm_fwd_addr_li[3:2];

  bsg_expand_bitmask_00000004_4
  \cache_pkt_sel_2_.non_max_size.mask_expand 
  (
    .i(\cache_pkt_sel_2_.non_max_size.decoded_slice_index ),
    .o({ cache_pkt_mask_mux_li_2__15_, cache_pkt_mask_mux_li_2__14_, cache_pkt_mask_mux_li_2__13_, cache_pkt_mask_mux_li_2__12_, cache_pkt_mask_mux_li_2__11_, cache_pkt_mask_mux_li_2__10_, cache_pkt_mask_mux_li_2__9_, cache_pkt_mask_mux_li_2__8_, cache_pkt_mask_mux_li_2__7_, cache_pkt_mask_mux_li_2__6_, cache_pkt_mask_mux_li_2__5_, cache_pkt_mask_mux_li_2__4_, cache_pkt_mask_mux_li_2__3_, cache_pkt_mask_mux_li_2__2_, cache_pkt_mask_mux_li_2__1_, cache_pkt_mask_mux_li_2__0_ })
  );

  assign \cache_pkt_sel_3_.non_max_size.decoded_slice_index  = { 1'b0, 1'b1 } << fsm_fwd_addr_li[3];

  bsg_expand_bitmask_00000002_8
  \cache_pkt_sel_3_.non_max_size.mask_expand 
  (
    .i(\cache_pkt_sel_3_.non_max_size.decoded_slice_index ),
    .o({ cache_pkt_mask_mux_li_3__15_, cache_pkt_mask_mux_li_3__14_, cache_pkt_mask_mux_li_3__13_, cache_pkt_mask_mux_li_3__12_, cache_pkt_mask_mux_li_3__11_, cache_pkt_mask_mux_li_3__10_, cache_pkt_mask_mux_li_3__9_, cache_pkt_mask_mux_li_3__8_, cache_pkt_mask_mux_li_3__7_, cache_pkt_mask_mux_li_3__6_, cache_pkt_mask_mux_li_3__5_, cache_pkt_mask_mux_li_3__4_, cache_pkt_mask_mux_li_3__3_, cache_pkt_mask_mux_li_3__2_, cache_pkt_mask_mux_li_3__1_, cache_pkt_mask_mux_li_3__0_ })
  );

  assign N70 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N69, N68, N67, N66, N65, N64, N63, N62 } > { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 };

  bsg_mux_00000010_00000005
  cache_pkt_mask_mux
  (
    .data_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, cache_pkt_mask_mux_li_3__15_, cache_pkt_mask_mux_li_3__14_, cache_pkt_mask_mux_li_3__13_, cache_pkt_mask_mux_li_3__12_, cache_pkt_mask_mux_li_3__11_, cache_pkt_mask_mux_li_3__10_, cache_pkt_mask_mux_li_3__9_, cache_pkt_mask_mux_li_3__8_, cache_pkt_mask_mux_li_3__7_, cache_pkt_mask_mux_li_3__6_, cache_pkt_mask_mux_li_3__5_, cache_pkt_mask_mux_li_3__4_, cache_pkt_mask_mux_li_3__3_, cache_pkt_mask_mux_li_3__2_, cache_pkt_mask_mux_li_3__1_, cache_pkt_mask_mux_li_3__0_, cache_pkt_mask_mux_li_2__15_, cache_pkt_mask_mux_li_2__14_, cache_pkt_mask_mux_li_2__13_, cache_pkt_mask_mux_li_2__12_, cache_pkt_mask_mux_li_2__11_, cache_pkt_mask_mux_li_2__10_, cache_pkt_mask_mux_li_2__9_, cache_pkt_mask_mux_li_2__8_, cache_pkt_mask_mux_li_2__7_, cache_pkt_mask_mux_li_2__6_, cache_pkt_mask_mux_li_2__5_, cache_pkt_mask_mux_li_2__4_, cache_pkt_mask_mux_li_2__3_, cache_pkt_mask_mux_li_2__2_, cache_pkt_mask_mux_li_2__1_, cache_pkt_mask_mux_li_2__0_, cache_pkt_mask_mux_li_1__15_, cache_pkt_mask_mux_li_1__14_, cache_pkt_mask_mux_li_1__13_, cache_pkt_mask_mux_li_1__12_, cache_pkt_mask_mux_li_1__11_, cache_pkt_mask_mux_li_1__10_, cache_pkt_mask_mux_li_1__9_, cache_pkt_mask_mux_li_1__8_, cache_pkt_mask_mux_li_1__7_, cache_pkt_mask_mux_li_1__6_, cache_pkt_mask_mux_li_1__5_, cache_pkt_mask_mux_li_1__4_, cache_pkt_mask_mux_li_1__3_, cache_pkt_mask_mux_li_1__2_, cache_pkt_mask_mux_li_1__1_, cache_pkt_mask_mux_li_1__0_, cache_pkt_mask_mux_li_0__15_, cache_pkt_mask_mux_li_0__14_, cache_pkt_mask_mux_li_0__13_, cache_pkt_mask_mux_li_0__12_, cache_pkt_mask_mux_li_0__11_, cache_pkt_mask_mux_li_0__10_, cache_pkt_mask_mux_li_0__9_, cache_pkt_mask_mux_li_0__8_, cache_pkt_mask_mux_li_0__7_, cache_pkt_mask_mux_li_0__6_, cache_pkt_mask_mux_li_0__5_, cache_pkt_mask_mux_li_0__4_, cache_pkt_mask_mux_li_0__3_, cache_pkt_mask_mux_li_0__2_, cache_pkt_mask_mux_li_0__1_, cache_pkt_mask_mux_li_0__0_ }),
    .sel_i(cache_pkt_sel_li),
    .data_o(cache_pkt_mask_lo)
  );


  bp_me_dram_hash_encode_00
  bank_select
  (
    .paddr_i(fsm_fwd_addr_li),
    .data_i(fsm_fwd_data_li),
    .dram_o(fwd_pkt_dram_lo),
    .daddr_o(fwd_pkt_daddr_lo),
    .slice_o(sv2v_dc_1),
    .bank_o(fwd_pkt_bank_lo[0]),
    .data_o(fwd_pkt_data_lo)
  );


  bsg_decode_with_v_00000002
  decode
  (
    .i(cache_fwd_bank_lo[0]),
    .v_i(cache_pkt_v_lo),
    .o(cache_pkt_v_o)
  );

  assign N73 = (N72)? cache_pkt_yumi_i[0] : 
               (N0)? cache_pkt_yumi_i[1] : 1'b0;
  assign N0 = cache_fwd_bank_lo[0];
  assign N82 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N81, N80, N79, N78, N77, N76, N75, N74 } > { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 };

  bsg_mux_00000080_00000002
  resp_bank_sel
  (
    .data_i(cache_data_i),
    .sel_i(fsm_rev_metadata_lo[65]),
    .data_o(cache_data_li)
  );


  bsg_bus_pack_00000080
  mem_rev_data_bus_pack
  (
    .data_i(cache_data_li),
    .sel_i({ 1'b0, 1'b0, 1'b0, 1'b0 }),
    .size_i(fsm_rev_size_li),
    .data_o(fsm_rev_data_lo)
  );

  assign N85 = N84 & N442;
  assign N86 = N85 & N443;
  assign N87 = state_r[2] | state_r[1];
  assign N88 = N87 | N443;
  assign N90 = state_r[2] | N442;
  assign N91 = N90 | state_r[0];
  assign N93 = state_r[2] | N442;
  assign N94 = N93 | N443;
  assign N96 = N84 | state_r[1];
  assign N97 = N96 | state_r[0];
  assign N99 = state_r[2] & state_r[0];
  assign N100 = state_r[2] & state_r[1];
  assign N109 = N108 | fsm_fwd_addr_li[4];
  assign N110 = fsm_fwd_addr_li[3] | fsm_fwd_addr_li[2];
  assign N111 = fsm_fwd_addr_li[1] | fsm_fwd_addr_li[0];
  assign N112 = N109 | N110;
  assign N113 = N112 | N111;
  assign N117 = N115 | fsm_fwd_addr_li[4];
  assign N118 = N116 | fsm_fwd_addr_li[2];
  assign N119 = fsm_fwd_addr_li[1] | fsm_fwd_addr_li[0];
  assign N120 = N117 | N118;
  assign N121 = N120 | N119;
  assign N125 = N123 | N124;
  assign N126 = fsm_fwd_addr_li[3] | fsm_fwd_addr_li[2];
  assign N127 = fsm_fwd_addr_li[1] | fsm_fwd_addr_li[0];
  assign N128 = N125 | N126;
  assign N129 = N128 | N127;
  assign N134 = N131 | N132;
  assign N135 = N133 | fsm_fwd_addr_li[2];
  assign N136 = fsm_fwd_addr_li[1] | fsm_fwd_addr_li[0];
  assign N137 = N134 | N135;
  assign N138 = N137 | N136;
  assign N160 = N140 & N141;
  assign N161 = N142 & N143;
  assign N162 = N144 & N145;
  assign N163 = N146 & N147;
  assign N164 = N148 & N149;
  assign N165 = N150 & N151;
  assign N166 = N152 & N153;
  assign N167 = N154 & N155;
  assign N168 = N156 & N157;
  assign N169 = N158 & N159;
  assign N170 = N160 & N161;
  assign N171 = N162 & N163;
  assign N172 = N164 & N165;
  assign N173 = N166 & N167;
  assign N174 = N168 & N169;
  assign N175 = N170 & N171;
  assign N176 = N172 & N173;
  assign N177 = N175 & N176;
  assign N178 = N177 & N174;
  assign N180 = fsm_fwd_addr_li[19] | fsm_fwd_addr_li[18];
  assign N181 = fsm_fwd_addr_li[17] | fsm_fwd_addr_li[16];
  assign N182 = fsm_fwd_addr_li[15] | fsm_fwd_addr_li[14];
  assign N183 = fsm_fwd_addr_li[13] | fsm_fwd_addr_li[12];
  assign N184 = fsm_fwd_addr_li[11] | fsm_fwd_addr_li[10];
  assign N185 = fsm_fwd_addr_li[9] | fsm_fwd_addr_li[8];
  assign N186 = fsm_fwd_addr_li[7] | fsm_fwd_addr_li[6];
  assign N187 = fsm_fwd_addr_li[5] | fsm_fwd_addr_li[4];
  assign N188 = N179 | fsm_fwd_addr_li[2];
  assign N189 = fsm_fwd_addr_li[1] | fsm_fwd_addr_li[0];
  assign N190 = N180 | N181;
  assign N191 = N182 | N183;
  assign N192 = N184 | N185;
  assign N193 = N186 | N187;
  assign N194 = N188 | N189;
  assign N195 = N190 | N191;
  assign N196 = N192 | N193;
  assign N197 = N195 | N196;
  assign N198 = N197 | N194;
  assign N201 = fsm_fwd_addr_li[19] | fsm_fwd_addr_li[18];
  assign N202 = fsm_fwd_addr_li[17] | fsm_fwd_addr_li[16];
  assign N203 = fsm_fwd_addr_li[15] | fsm_fwd_addr_li[14];
  assign N204 = fsm_fwd_addr_li[13] | fsm_fwd_addr_li[12];
  assign N205 = fsm_fwd_addr_li[11] | fsm_fwd_addr_li[10];
  assign N206 = fsm_fwd_addr_li[9] | fsm_fwd_addr_li[8];
  assign N207 = fsm_fwd_addr_li[7] | fsm_fwd_addr_li[6];
  assign N208 = fsm_fwd_addr_li[5] | N200;
  assign N209 = fsm_fwd_addr_li[3] | fsm_fwd_addr_li[2];
  assign N210 = fsm_fwd_addr_li[1] | fsm_fwd_addr_li[0];
  assign N211 = N201 | N202;
  assign N212 = N203 | N204;
  assign N213 = N205 | N206;
  assign N214 = N207 | N208;
  assign N215 = N209 | N210;
  assign N216 = N211 | N212;
  assign N217 = N213 | N214;
  assign N218 = N216 | N217;
  assign N219 = N218 | N215;
  assign N223 = fsm_fwd_addr_li[19] | fsm_fwd_addr_li[18];
  assign N224 = fsm_fwd_addr_li[17] | fsm_fwd_addr_li[16];
  assign N225 = fsm_fwd_addr_li[15] | fsm_fwd_addr_li[14];
  assign N226 = fsm_fwd_addr_li[13] | fsm_fwd_addr_li[12];
  assign N227 = fsm_fwd_addr_li[11] | fsm_fwd_addr_li[10];
  assign N228 = fsm_fwd_addr_li[9] | fsm_fwd_addr_li[8];
  assign N229 = fsm_fwd_addr_li[7] | fsm_fwd_addr_li[6];
  assign N230 = fsm_fwd_addr_li[5] | N221;
  assign N231 = N222 | fsm_fwd_addr_li[2];
  assign N232 = fsm_fwd_addr_li[1] | fsm_fwd_addr_li[0];
  assign N233 = N223 | N224;
  assign N234 = N225 | N226;
  assign N235 = N227 | N228;
  assign N236 = N229 | N230;
  assign N237 = N231 | N232;
  assign N238 = N233 | N234;
  assign N239 = N235 | N236;
  assign N240 = N238 | N239;
  assign N241 = N240 | N237;
  assign N260 = N258 & N259;
  assign N264 = N262 & N263;
  assign N266 = fsm_fwd_header_li[1] | N265;
  assign N268 = N267 | fsm_fwd_header_li[0];
  assign N270 = fsm_fwd_header_li[1] & fsm_fwd_header_li[0];
  assign N274 = N272 & N273;
  assign N276 = fsm_fwd_header_li[49] | N275;
  assign N279 = N278 | fsm_fwd_header_li[48];
  assign N281 = fsm_fwd_header_li[49] & fsm_fwd_header_li[48];
  assign N291 = N289 & N290;
  assign N293 = fsm_fwd_header_li[49] | N292;
  assign N296 = N295 | fsm_fwd_header_li[48];
  assign N297 = fsm_fwd_header_li[49] & fsm_fwd_header_li[48];
  assign N303 = N299 & N300;
  assign N304 = N301 & N302;
  assign N305 = N303 & N304;
  assign N308 = fsm_fwd_header_li[7] | fsm_fwd_header_li[6];
  assign N309 = N306 | N307;
  assign N310 = N308 | N309;
  assign N313 = fsm_fwd_header_li[7] | N312;
  assign N314 = fsm_fwd_header_li[5] | fsm_fwd_header_li[4];
  assign N315 = N313 | N314;
  assign N319 = fsm_fwd_header_li[7] | N317;
  assign N320 = fsm_fwd_header_li[5] | N318;
  assign N321 = N319 | N320;
  assign N325 = fsm_fwd_header_li[7] | N323;
  assign N326 = N324 | fsm_fwd_header_li[4];
  assign N327 = N325 | N326;
  assign N332 = fsm_fwd_header_li[7] | N329;
  assign N333 = N330 | N331;
  assign N334 = N332 | N333;
  assign N337 = N336 | fsm_fwd_header_li[6];
  assign N338 = fsm_fwd_header_li[5] | fsm_fwd_header_li[4];
  assign N339 = N337 | N338;
  assign N343 = N341 | fsm_fwd_header_li[6];
  assign N344 = fsm_fwd_header_li[5] | N342;
  assign N345 = N343 | N344;
  assign N349 = N347 | fsm_fwd_header_li[6];
  assign N350 = N348 | fsm_fwd_header_li[4];
  assign N351 = N349 | N350;
  assign N356 = N353 | fsm_fwd_header_li[6];
  assign N357 = N354 | N355;
  assign N358 = N356 | N357;
  assign N361 = fsm_fwd_header_li[7] | fsm_fwd_header_li[6];
  assign N362 = fsm_fwd_header_li[5] | N360;
  assign N363 = N361 | N362;
  assign N365 = fsm_fwd_header_li[7] | fsm_fwd_header_li[6];
  assign N366 = N364 | fsm_fwd_header_li[4];
  assign N367 = N365 | N366;
  assign N368 = fsm_fwd_header_li[7] & fsm_fwd_header_li[6];
  assign N442 = ~state_r[1];
  assign N443 = ~state_r[0];
  assign N444 = N442 | state_r[2];
  assign N445 = N443 | N444;
  assign N446 = ~N445;
  assign N447 = ~fsm_rev_metadata_lo[65];
  assign N448 = set_cnt[9] & set_cnt[10];
  assign N449 = set_cnt[8] & N448;
  assign N450 = set_cnt[7] & N449;
  assign N451 = set_cnt[6] & N450;
  assign N452 = set_cnt[5] & N451;
  assign N453 = set_cnt[4] & N452;
  assign N454 = set_cnt[3] & N453;
  assign N455 = set_cnt[2] & N454;
  assign N456 = set_cnt[1] & N455;
  assign N457 = set_cnt[0] & N456;
  assign N458 = ~fsm_fwd_header_li[49];
  assign N459 = N458 | fsm_fwd_header_li[50];
  assign N460 = fsm_fwd_header_li[48] | N459;
  assign N461 = state_r[1] | state_r[2];
  assign N462 = N443 | N461;
  assign N463 = ~N462;
  assign { N69, N68, N67, N66, N65, N64, N63, N62 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fsm_fwd_header_li[50:48];
  assign { N81, N80, N79, N78, N77, N76, N75, N74 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fsm_rev_metadata_lo[50:48];
  assign cache_pkt_sel_li = (N1)? { 1'b1, 1'b0, 1'b0 } : 
                            (N71)? fsm_fwd_header_li[50:48] : 1'b0;
  assign N1 = N70;
  assign cache_fwd_bank_lo[0] = (N2)? set_cnt[10] : 
                                (N3)? fwd_pkt_bank_lo[0] : 1'b0;
  assign N2 = N463;
  assign N3 = N462;
  assign fsm_rev_size_li = (N4)? { 1'b1, 1'b0, 1'b0 } : 
                           (N83)? fsm_rev_metadata_lo[50:48] : 1'b0;
  assign N4 = N82;
  assign N106 = ~N105;
  assign N251 = ~fwd_pkt_data_lo[0];
  assign { N257, N256, N253, N252 } = (N5)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                                      (N6)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                                      (N7)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                      (N8)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                      (N9)? { 1'b1, 1'b1, 1'b0, 1'b0 } : 
                                      (N10)? { 1'b1, 1'b1, 1'b0, 1'b1 } : 
                                      (N11)? { 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                      (N12)? { 1'b1, 1'b1, fwd_pkt_data_lo[0:0], fwd_pkt_data_lo[0:0] } : 
                                      (N250)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N5 = N114;
  assign N6 = N122;
  assign N7 = N130;
  assign N8 = N139;
  assign N9 = N178;
  assign N10 = N199;
  assign N11 = N220;
  assign N12 = N242;
  assign N255 = (N12)? N251 : 
                (N254)? 1'b0 : 1'b0;
  assign { N283, N282 } = (N13)? { 1'b0, 1'b0 } : 
                          (N14)? { 1'b0, 1'b1 } : 
                          (N15)? { 1'b1, 1'b0 } : 
                          (N16)? { 1'b1, 1'b1 } : 1'b0;
  assign N13 = N274;
  assign N14 = N277;
  assign N15 = N280;
  assign N16 = N281;
  assign { N285, N284 } = (N17)? { N283, N282 } : 
                          (N18)? { 1'b0, 1'b0 } : 1'b0;
  assign N17 = N271;
  assign N18 = N286;
  assign { N375, N374, N373, N372, N371, N370 } = (N19)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, N460 } : 
                                                  (N20)? { 1'b1, N460, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                  (N21)? { 1'b1, N460, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                                  (N22)? { 1'b1, N460, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                                  (N23)? { 1'b1, N460, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                  (N24)? { 1'b1, N460, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                                  (N25)? { 1'b1, N460, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                                  (N26)? { 1'b1, N460, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                                  (N27)? { 1'b1, N460, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                  (N28)? { 1'b1, N460, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                                  (N29)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N19 = N305;
  assign N20 = N311;
  assign N21 = N316;
  assign N22 = N322;
  assign N23 = N328;
  assign N24 = N335;
  assign N25 = N340;
  assign N26 = N346;
  assign N27 = N352;
  assign N28 = N359;
  assign N29 = N369;
  assign { N381, N376 } = (N30)? { 1'b1, 1'b0 } : 
                          (N31)? { 1'b1, 1'b1 } : 
                          (N32)? { N373, N370 } : 1'b0;
  assign N30 = N291;
  assign N31 = N294;
  assign N32 = N298;
  assign { N383, N382, N380, N379 } = (N32)? { N375, N374, N372, N371 } : 
                                      (N378)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N389, N388, N387, N386, N385, N384 } = (N33)? { N383, N382, N381, N380, N379, N376 } : 
                                                  (N34)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1 } : 1'b0;
  assign N33 = N287;
  assign N34 = N288;
  assign { N393, N392, N391, N390 } = (N35)? { N286, N286, N285, N284 } : 
                                      (N36)? { N387, N386, N385, N384 } : 
                                      (N37)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N35 = N264;
  assign N36 = N269;
  assign N37 = N270;
  assign { N397, N396 } = (N36)? { N389, N388 } : 
                          (N395)? { 1'b0, 1'b0 } : 1'b0;
  assign { N403, N402, N401, N400, N399, N398 } = (N38)? { N397, N396, N393, N392, N391, N390 } : 
                                                  (N261)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N38 = N260;
  assign { N409, N408, N407, N406, N405, N404 } = (N39)? { 1'b0, N257, N256, N255, N253, N252 } : 
                                                  (N40)? { N403, N402, N401, N400, N399, N398 } : 1'b0;
  assign N39 = N107;
  assign N40 = fwd_pkt_dram_lo;
  assign { N416, N415, N414 } = (N41)? { 1'b1, 1'b0, 1'b0 } : 
                                (N413)? state_r : 1'b0;
  assign N41 = N412;
  assign N417 = (N42)? N411 : 
                (N43)? cache_pkt_yumi_li : 1'b0;
  assign N42 = is_uc_op;
  assign N43 = N410;
  assign { N420, N419, N418 } = (N42)? { N416, N415, N414 } : 
                                (N43)? state_r : 1'b0;
  assign { N424, N423, N422 } = (N44)? { 1'b0, 1'b1, 1'b0 } : 
                                (N45)? state_r : 1'b0;
  assign N44 = cache_pkt_yumi_li;
  assign N45 = N421;
  assign state_n = (N46)? { 1'b0, 1'b0, 1'b1 } : 
                   (N47)? { 1'b0, N103, N104 } : 
                   (N48)? { 1'b0, 1'b1, N106 } : 
                   (N49)? { N420, N419, N418 } : 
                   (N50)? { N424, N423, N422 } : 1'b0;
  assign N46 = N86;
  assign N47 = N89;
  assign N48 = N92;
  assign N49 = N95;
  assign N50 = N98;
  assign cache_pkt_v_lo = (N46)? 1'b0 : 
                          (N47)? 1'b1 : 
                          (N48)? 1'b0 : 
                          (N49)? fsm_fwd_v_li : 
                          (N50)? fsm_fwd_v_li : 
                          (N51)? 1'b0 : 1'b0;
  assign N51 = N101;
  assign { cache_pkt_o_1__181_, cache_pkt_o_1__180_, cache_pkt_o_1__177_, cache_pkt_o_1__176_, cache_pkt_o_1__175_, cache_pkt_o_1__174_, cache_pkt_o_1__173_, cache_pkt_o_1__172_, cache_pkt_o_1__171_, cache_pkt_o_1__170_, cache_pkt_o_1__169_, cache_pkt_o_1__168_, cache_pkt_o_1__167_, cache_pkt_o_1__166_, cache_pkt_o_1__165_, cache_pkt_o_1__164_, cache_pkt_o_1__163_, cache_pkt_o_1__162_, cache_pkt_o_1__161_, cache_pkt_o_1__160_, cache_pkt_o_1__159_, cache_pkt_o_1__158_, cache_pkt_o_1__157_, cache_pkt_o_1__156_, cache_pkt_o_1__155_, cache_pkt_o_1__154_, cache_pkt_o_1__153_, cache_pkt_o_1__152_, cache_pkt_o_1__151_, cache_pkt_o_1__150_, cache_pkt_o_1__149_, cache_pkt_o_1__148_, cache_pkt_o_1__147_, cache_pkt_o_1__146_, cache_pkt_o_1__145_, cache_pkt_o_1__144_, cache_pkt_o_1__143_, cache_pkt_o_1__142_, cache_pkt_o_1__141_, cache_pkt_o_1__140_, cache_pkt_o_1__139_, cache_pkt_o_1__138_, cache_pkt_o_1__137_, cache_pkt_o_1__136_, cache_pkt_o_1__135_, cache_pkt_o_1__134_, cache_pkt_o_1__133_, cache_pkt_o_1__132_, cache_pkt_o_1__131_, cache_pkt_o_1__130_, cache_pkt_o_1__129_, cache_pkt_o_1__128_, cache_pkt_o_1__127_, cache_pkt_o_1__126_, cache_pkt_o_1__125_, cache_pkt_o_1__124_, cache_pkt_o_1__123_, cache_pkt_o_1__122_, cache_pkt_o_1__121_, cache_pkt_o_1__120_, cache_pkt_o_1__119_, cache_pkt_o_1__118_, cache_pkt_o_1__117_, cache_pkt_o_1__116_, cache_pkt_o_1__115_, cache_pkt_o_1__114_, cache_pkt_o_1__113_, cache_pkt_o_1__112_, cache_pkt_o_1__111_, cache_pkt_o_1__110_, cache_pkt_o_1__109_, cache_pkt_o_1__108_, cache_pkt_o_1__107_, cache_pkt_o_1__106_, cache_pkt_o_1__105_, cache_pkt_o_1__104_, cache_pkt_o_1__103_, cache_pkt_o_1__102_, cache_pkt_o_1__101_, cache_pkt_o_1__100_, cache_pkt_o_1__99_, cache_pkt_o_1__98_, cache_pkt_o_1__97_, cache_pkt_o_1__96_, cache_pkt_o_1__95_, cache_pkt_o_1__94_, cache_pkt_o_1__93_, cache_pkt_o_1__92_, cache_pkt_o_1__91_, cache_pkt_o_1__90_, cache_pkt_o_1__89_, cache_pkt_o_1__88_, cache_pkt_o_1__87_, cache_pkt_o_1__86_, cache_pkt_o_1__85_, cache_pkt_o_1__84_, cache_pkt_o_1__83_, cache_pkt_o_1__82_, cache_pkt_o_1__81_, cache_pkt_o_1__80_, cache_pkt_o_1__79_, cache_pkt_o_1__78_, cache_pkt_o_1__77_, cache_pkt_o_1__76_, cache_pkt_o_1__75_, cache_pkt_o_1__74_, cache_pkt_o_1__73_, cache_pkt_o_1__72_, cache_pkt_o_1__71_, cache_pkt_o_1__70_, cache_pkt_o_1__69_, cache_pkt_o_1__68_, cache_pkt_o_1__67_, cache_pkt_o_1__66_, cache_pkt_o_1__65_, cache_pkt_o_1__64_, cache_pkt_o_1__63_, cache_pkt_o_1__62_, cache_pkt_o_1__61_, cache_pkt_o_1__60_, cache_pkt_o_1__59_, cache_pkt_o_1__58_, cache_pkt_o_1__57_, cache_pkt_o_1__56_, cache_pkt_o_1__55_, cache_pkt_o_1__54_, cache_pkt_o_1__53_, cache_pkt_o_1__52_, cache_pkt_o_1__51_, cache_pkt_o_1__50_, cache_pkt_o_1__49_, cache_pkt_o_1__48_, cache_pkt_o_1__47_, cache_pkt_o_1__46_, cache_pkt_o_1__45_, cache_pkt_o_1__44_, cache_pkt_o_1__43_, cache_pkt_o_1__42_, cache_pkt_o_1__41_, cache_pkt_o_1__40_, cache_pkt_o_1__39_, cache_pkt_o_1__38_, cache_pkt_o_1__37_, cache_pkt_o_1__36_, cache_pkt_o_1__35_, cache_pkt_o_1__34_, cache_pkt_o_1__33_, cache_pkt_o_1__32_, cache_pkt_o_1__31_, cache_pkt_o_1__30_, cache_pkt_o_1__29_, cache_pkt_o_1__28_, cache_pkt_o_1__27_, cache_pkt_o_1__26_, cache_pkt_o_1__25_, cache_pkt_o_1__24_, cache_pkt_o_1__23_, cache_pkt_o_1__22_, cache_pkt_o_1__21_, cache_pkt_o_1__20_, cache_pkt_o_1__19_, cache_pkt_o_1__18_, cache_pkt_o_1__17_, cache_pkt_o_1__16_, cache_pkt_o_1__15_, cache_pkt_o_1__14_, cache_pkt_o_1__13_, cache_pkt_o_1__12_, cache_pkt_o_1__11_, cache_pkt_o_1__10_, cache_pkt_o_1__9_, cache_pkt_o_1__8_, cache_pkt_o_1__7_, cache_pkt_o_1__6_, cache_pkt_o_1__5_, cache_pkt_o_1__4_, cache_pkt_o_1__3_, cache_pkt_o_1__2_, cache_pkt_o_1__1_, cache_pkt_o_1__0_ } = (N46)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N47)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, set_cnt, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N48)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N49)? { N408, N407, N404, fwd_pkt_daddr_lo, fwd_pkt_data_lo, cache_pkt_mask_lo } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N50)? { 1'b1, 1'b1, 1'b1, fwd_pkt_daddr_lo, fwd_pkt_data_lo, cache_pkt_mask_lo } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N51)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { cache_pkt_o_1__182_, cache_pkt_o_1__179_, cache_pkt_o_1__178_ } = (N49)? { N409, N406, N405 } : 
                                                                             (N425)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign set_up = (N46)? 1'b0 : 
                  (N47)? N102 : 
                  (N48)? 1'b0 : 
                  (N49)? 1'b0 : 
                  (N50)? 1'b0 : 
                  (N51)? 1'b0 : 1'b0;
  assign set_clear = (N46)? 1'b0 : 
                     (N47)? N103 : 
                     (N48)? 1'b0 : 
                     (N49)? 1'b0 : 
                     (N50)? 1'b0 : 
                     (N51)? 1'b0 : 1'b0;
  assign { N427, N426 } = (N46)? { 1'b0, 1'b0 } : 
                          (N47)? cache_data_v_i : 
                          (N48)? cache_data_v_i : 
                          (N49)? { 1'b0, 1'b0 } : 
                          (N50)? { 1'b0, 1'b0 } : 
                          (N51)? { 1'b0, 1'b0 } : 1'b0;
  assign fsm_fwd_yumi_lo = (N46)? 1'b0 : 
                           (N47)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N49)? N417 : 
                           (N50)? cache_pkt_yumi_li : 
                           (N51)? 1'b0 : 1'b0;
  assign N433 = (N52)? cache_data_v_i[0] : 
                (N53)? N426 : 1'b0;
  assign N52 = N431;
  assign N53 = N432;
  assign N434 = (N54)? N430 : 
                (N55)? 1'b0 : 1'b0;
  assign N54 = N428;
  assign N55 = N429;
  assign cache_data_yumi_o[0] = (N54)? N430 : 
                                (N55)? N433 : 1'b0;
  assign N440 = (N56)? cache_data_v_i[1] : 
                (N57)? N427 : 1'b0;
  assign N56 = N438;
  assign N57 = N439;
  assign fsm_rev_v_lo = (N58)? N437 : 
                        (N59)? N434 : 1'b0;
  assign N58 = N435;
  assign N59 = N436;
  assign cache_data_yumi_o[1] = (N58)? N437 : 
                                (N59)? N440 : 1'b0;
  assign is_uc_op = N60 & N61;
  assign N71 = ~N70;
  assign N72 = ~cache_fwd_bank_lo[0];
  assign cache_pkt_yumi_li = fsm_fwd_v_li & N73;
  assign N83 = ~N82;
  assign N84 = ~state_r[2];
  assign N89 = ~N88;
  assign N92 = ~N91;
  assign N95 = ~N94;
  assign N98 = ~N97;
  assign N101 = N99 | N100;
  assign N102 = ~N457;
  assign N103 = N457 & N464;
  assign N464 = cache_pkt_yumi_i[1] | cache_pkt_yumi_i[0];
  assign N104 = ~N103;
  assign N105 = cache_data_v_i[1] | N465;
  assign N465 = fsm_rev_ready_then_li | cache_data_v_i[0];
  assign N107 = ~fwd_pkt_dram_lo;
  assign N108 = ~fsm_fwd_addr_li[5];
  assign N114 = ~N113;
  assign N115 = ~fsm_fwd_addr_li[5];
  assign N116 = ~fsm_fwd_addr_li[3];
  assign N122 = ~N121;
  assign N123 = ~fsm_fwd_addr_li[5];
  assign N124 = ~fsm_fwd_addr_li[4];
  assign N130 = ~N129;
  assign N131 = ~fsm_fwd_addr_li[5];
  assign N132 = ~fsm_fwd_addr_li[4];
  assign N133 = ~fsm_fwd_addr_li[3];
  assign N139 = ~N138;
  assign N140 = ~fsm_fwd_addr_li[19];
  assign N141 = ~fsm_fwd_addr_li[18];
  assign N142 = ~fsm_fwd_addr_li[17];
  assign N143 = ~fsm_fwd_addr_li[16];
  assign N144 = ~fsm_fwd_addr_li[15];
  assign N145 = ~fsm_fwd_addr_li[14];
  assign N146 = ~fsm_fwd_addr_li[13];
  assign N147 = ~fsm_fwd_addr_li[12];
  assign N148 = ~fsm_fwd_addr_li[11];
  assign N149 = ~fsm_fwd_addr_li[10];
  assign N150 = ~fsm_fwd_addr_li[9];
  assign N151 = ~fsm_fwd_addr_li[8];
  assign N152 = ~fsm_fwd_addr_li[7];
  assign N153 = ~fsm_fwd_addr_li[6];
  assign N154 = ~fsm_fwd_addr_li[5];
  assign N155 = ~fsm_fwd_addr_li[4];
  assign N156 = ~fsm_fwd_addr_li[3];
  assign N157 = ~fsm_fwd_addr_li[2];
  assign N158 = ~fsm_fwd_addr_li[1];
  assign N159 = ~fsm_fwd_addr_li[0];
  assign N179 = ~fsm_fwd_addr_li[3];
  assign N199 = ~N198;
  assign N200 = ~fsm_fwd_addr_li[4];
  assign N220 = ~N219;
  assign N221 = ~fsm_fwd_addr_li[4];
  assign N222 = ~fsm_fwd_addr_li[3];
  assign N242 = ~N241;
  assign N243 = N122 | N114;
  assign N244 = N130 | N243;
  assign N245 = N139 | N244;
  assign N246 = N178 | N245;
  assign N247 = N199 | N246;
  assign N248 = N220 | N247;
  assign N249 = N242 | N248;
  assign N250 = ~N249;
  assign N254 = N241;
  assign N258 = ~fsm_fwd_header_li[3];
  assign N259 = ~fsm_fwd_header_li[2];
  assign N261 = ~N260;
  assign N262 = ~fsm_fwd_header_li[1];
  assign N263 = ~fsm_fwd_header_li[0];
  assign N265 = ~fsm_fwd_header_li[0];
  assign N267 = ~fsm_fwd_header_li[1];
  assign N269 = N466 | N467;
  assign N466 = ~N266;
  assign N467 = ~N268;
  assign N271 = ~fsm_fwd_header_li[50];
  assign N286 = fsm_fwd_header_li[50];
  assign N272 = ~fsm_fwd_header_li[49];
  assign N273 = ~fsm_fwd_header_li[48];
  assign N275 = ~fsm_fwd_header_li[48];
  assign N277 = ~N276;
  assign N278 = ~fsm_fwd_header_li[49];
  assign N280 = ~N279;
  assign N287 = ~fsm_fwd_header_li[50];
  assign N288 = fsm_fwd_header_li[50];
  assign N289 = ~fsm_fwd_header_li[49];
  assign N290 = ~fsm_fwd_header_li[48];
  assign N292 = ~fsm_fwd_header_li[48];
  assign N294 = ~N293;
  assign N295 = ~fsm_fwd_header_li[49];
  assign N298 = N468 | N297;
  assign N468 = ~N296;
  assign N299 = ~fsm_fwd_header_li[7];
  assign N300 = ~fsm_fwd_header_li[6];
  assign N301 = ~fsm_fwd_header_li[5];
  assign N302 = ~fsm_fwd_header_li[4];
  assign N306 = ~fsm_fwd_header_li[5];
  assign N307 = ~fsm_fwd_header_li[4];
  assign N311 = ~N310;
  assign N312 = ~fsm_fwd_header_li[6];
  assign N316 = ~N315;
  assign N317 = ~fsm_fwd_header_li[6];
  assign N318 = ~fsm_fwd_header_li[4];
  assign N322 = ~N321;
  assign N323 = ~fsm_fwd_header_li[6];
  assign N324 = ~fsm_fwd_header_li[5];
  assign N328 = ~N327;
  assign N329 = ~fsm_fwd_header_li[6];
  assign N330 = ~fsm_fwd_header_li[5];
  assign N331 = ~fsm_fwd_header_li[4];
  assign N335 = ~N334;
  assign N336 = ~fsm_fwd_header_li[7];
  assign N340 = ~N339;
  assign N341 = ~fsm_fwd_header_li[7];
  assign N342 = ~fsm_fwd_header_li[4];
  assign N346 = ~N345;
  assign N347 = ~fsm_fwd_header_li[7];
  assign N348 = ~fsm_fwd_header_li[5];
  assign N352 = ~N351;
  assign N353 = ~fsm_fwd_header_li[7];
  assign N354 = ~fsm_fwd_header_li[5];
  assign N355 = ~fsm_fwd_header_li[4];
  assign N359 = ~N358;
  assign N360 = ~fsm_fwd_header_li[4];
  assign N364 = ~fsm_fwd_header_li[5];
  assign N369 = N469 | N471;
  assign N469 = ~N363;
  assign N471 = N470 | N368;
  assign N470 = ~N367;
  assign N377 = ~N298;
  assign N378 = N377;
  assign N394 = ~N269;
  assign N395 = N394;
  assign N410 = ~is_uc_op;
  assign N411 = cache_pkt_yumi_li & N472;
  assign N472 = ~fsm_fwd_last_li;
  assign N412 = N473 & cache_pkt_yumi_li;
  assign N473 = fsm_fwd_v_li & fsm_fwd_last_li;
  assign N413 = ~N412;
  assign N421 = ~cache_pkt_yumi_li;
  assign N425 = N94;
  assign N428 = N474 & N447;
  assign N474 = op_v_lo[0] & op_data_lo[0];
  assign N429 = ~N428;
  assign N430 = fsm_rev_ready_then_li & cache_data_v_i[0];
  assign N431 = op_v_lo[0] & N475;
  assign N475 = ~op_data_lo[0];
  assign N432 = ~N431;
  assign N435 = N476 & fsm_rev_metadata_lo[65];
  assign N476 = op_v_lo[1] & op_data_lo[1];
  assign N436 = ~N435;
  assign N437 = fsm_rev_ready_then_li & cache_data_v_i[1];
  assign N438 = op_v_lo[1] & N477;
  assign N477 = ~op_data_lo[1];
  assign N439 = ~N438;
  assign N441 = ~N101;

  always @(posedge clk_i) begin
    if(reset_i) begin
      state_r_2_sv2v_reg <= 1'b0;
      state_r_1_sv2v_reg <= 1'b0;
      state_r_0_sv2v_reg <= 1'b0;
    end else if(N441) begin
      state_r_2_sv2v_reg <= state_n[2];
      state_r_1_sv2v_reg <= state_n[1];
      state_r_0_sv2v_reg <= state_n[0];
    end 
  end


endmodule



module bsg_cache_decode
(
  opcode_i,
  decode_o
);

  input [5:0] opcode_i;
  output [20:0] decode_o;
  wire [20:0] decode_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N146,N147,N148,N150,N152,
  N153,N154,N155,N156,N158,N160,N161,N163,N165,N166,N167,N168,N170,N171,N172,N173,
  N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,
  N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,
  N206,N207,N208,N209,N210,N211,N212,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297;
  assign N17 = N80 | N138;
  assign N18 = opcode_i[3] | opcode_i[2];
  assign N19 = opcode_i[1] | opcode_i[0];
  assign N20 = N17 | N18;
  assign N21 = N20 | N19;
  assign N22 = opcode_i[1] | N139;
  assign N23 = N20 | N22;
  assign N24 = N146 | N139;
  assign N25 = N20 | N24;
  assign N26 = opcode_i[3] | N165;
  assign N27 = N17 | N26;
  assign N28 = N27 | N19;
  assign N29 = N146 | opcode_i[0];
  assign N30 = N20 | N29;
  assign N31 = N27 | N22;
  assign N32 = N27 | N29;
  assign N33 = N27 | N24;
  assign N34 = N152 | opcode_i[2];
  assign N35 = N17 | N34;
  assign N36 = N35 | N19;
  assign N37 = opcode_i[5] | opcode_i[4];
  assign N38 = N37 | N18;
  assign N39 = N38 | N24;
  assign N40 = N37 | N34;
  assign N41 = N40 | N24;
  assign N42 = N37 | N26;
  assign N43 = N42 | N24;
  assign N45 = N80 | opcode_i[4];
  assign N46 = N45 | N18;
  assign N47 = N46 | N19;
  assign N48 = N46 | N22;
  assign N49 = N46 | N24;
  assign N50 = N45 | N26;
  assign N51 = N50 | N19;
  assign N52 = N46 | N29;
  assign N53 = N50 | N22;
  assign N54 = N50 | N29;
  assign N55 = N50 | N24;
  assign N56 = N45 | N34;
  assign N57 = N56 | N19;
  assign N58 = N38 | N29;
  assign N59 = N40 | N29;
  assign N60 = N42 | N29;
  assign N62 = N38 | N22;
  assign N63 = N40 | N22;
  assign N64 = N42 | N22;
  assign N66 = N80 & N138;
  assign N67 = N152 & N165;
  assign N68 = N146 & N139;
  assign N69 = N66 & N67;
  assign N70 = N69 & N68;
  assign N71 = N40 | N19;
  assign N72 = N42 | N19;
  assign N74 = opcode_i[5] & opcode_i[3];
  assign N75 = N74 & opcode_i[0];
  assign N76 = N74 & opcode_i[1];
  assign N77 = opcode_i[3] & opcode_i[2];
  assign N78 = N80 & opcode_i[4];
  assign N81 = N138 & N152;
  assign N82 = N165 & N146;
  assign N83 = N81 & N82;
  assign N84 = N83 & N139;
  assign N85 = N138 | opcode_i[3];
  assign N86 = opcode_i[2] | opcode_i[1];
  assign N87 = N85 | N86;
  assign N88 = N87 | opcode_i[0];
  assign N90 = opcode_i[4] | opcode_i[3];
  assign N91 = N90 | N86;
  assign N92 = N91 | N139;
  assign N93 = N87 | N139;
  assign N95 = opcode_i[2] | N146;
  assign N96 = N90 | N95;
  assign N97 = N96 | opcode_i[0];
  assign N98 = N85 | N95;
  assign N99 = N98 | opcode_i[0];
  assign N101 = N96 | N139;
  assign N102 = N98 | N139;
  assign N104 = N165 | opcode_i[1];
  assign N105 = N90 | N104;
  assign N106 = N105 | opcode_i[0];
  assign N107 = N85 | N104;
  assign N108 = N107 | opcode_i[0];
  assign N110 = N105 | N139;
  assign N111 = N107 | N139;
  assign N113 = N165 | N146;
  assign N114 = N90 | N113;
  assign N115 = N114 | opcode_i[0];
  assign N116 = N85 | N113;
  assign N117 = N116 | opcode_i[0];
  assign N119 = N114 | N139;
  assign N120 = N116 | N139;
  assign N122 = opcode_i[4] | N152;
  assign N123 = N122 | N86;
  assign N124 = N123 | opcode_i[0];
  assign N125 = N138 | N152;
  assign N126 = N125 | N86;
  assign N127 = N126 | opcode_i[0];
  assign N129 = opcode_i[3] & opcode_i[0];
  assign N130 = opcode_i[3] & opcode_i[1];
  assign N138 = ~opcode_i[4];
  assign N139 = ~opcode_i[0];
  assign N140 = N138 | opcode_i[5];
  assign N141 = opcode_i[3] | N140;
  assign N142 = opcode_i[2] | N141;
  assign N143 = opcode_i[1] | N142;
  assign N144 = N139 | N143;
  assign decode_o[13] = ~N144;
  assign N146 = ~opcode_i[1];
  assign N147 = N146 | N142;
  assign N148 = opcode_i[0] | N147;
  assign decode_o[12] = ~N148;
  assign N150 = N139 | N147;
  assign decode_o[11] = ~N150;
  assign N152 = ~opcode_i[3];
  assign N153 = N152 | N140;
  assign N154 = opcode_i[2] | N153;
  assign N155 = opcode_i[1] | N154;
  assign N156 = opcode_i[0] | N155;
  assign decode_o[10] = ~N156;
  assign N158 = N139 | N155;
  assign decode_o[9] = ~N158;
  assign N160 = N146 | N154;
  assign N161 = opcode_i[0] | N160;
  assign decode_o[8] = ~N161;
  assign N163 = N139 | N160;
  assign decode_o[7] = ~N163;
  assign N165 = ~opcode_i[2];
  assign N166 = N165 | N153;
  assign N167 = opcode_i[1] | N166;
  assign N168 = opcode_i[0] | N167;
  assign decode_o[6] = ~N168;
  assign N170 = opcode_i[4] | opcode_i[5];
  assign N171 = opcode_i[3] | N170;
  assign N172 = opcode_i[2] | N171;
  assign N173 = opcode_i[1] | N172;
  assign N174 = opcode_i[0] | N173;
  assign N175 = ~N174;
  assign N176 = N139 | N173;
  assign N177 = ~N176;
  assign N178 = N146 | N172;
  assign N179 = opcode_i[0] | N178;
  assign N180 = ~N179;
  assign N181 = N139 | N178;
  assign N182 = ~N181;
  assign N183 = N152 | N170;
  assign N184 = N165 | N183;
  assign N185 = opcode_i[1] | N184;
  assign N186 = opcode_i[0] | N185;
  assign N187 = ~N186;
  assign N188 = N139 | N185;
  assign N189 = ~N188;
  assign N190 = N165 | N171;
  assign N191 = opcode_i[1] | N190;
  assign N192 = opcode_i[0] | N191;
  assign N193 = ~N192;
  assign N194 = N139 | N191;
  assign N195 = ~N194;
  assign N196 = N146 | N190;
  assign N197 = opcode_i[0] | N196;
  assign N198 = ~N197;
  assign N199 = N139 | N196;
  assign N200 = ~N199;
  assign N201 = opcode_i[2] | N183;
  assign N202 = opcode_i[1] | N201;
  assign N203 = opcode_i[0] | N202;
  assign N204 = ~N203;
  assign N205 = N139 | N202;
  assign N206 = ~N205;
  assign N207 = N146 | N201;
  assign N208 = opcode_i[0] | N207;
  assign N209 = ~N208;
  assign N210 = N139 | N207;
  assign N211 = ~N210;
  assign N212 = opcode_i[0] | N143;
  assign decode_o[14] = ~N212;
  assign decode_o[20:19] = (N0)? { 1'b1, 1'b1 } : 
                           (N1)? { 1'b1, 1'b0 } : 
                           (N2)? { 1'b0, 1'b1 } : 
                           (N3)? { 1'b0, 1'b0 } : 
                           (N4)? { 1'b0, 1'b0 } : 1'b0;
  assign N0 = N44;
  assign N1 = N61;
  assign N2 = N65;
  assign N3 = N73;
  assign N4 = N79;
  assign { N135, N134, N133, N132 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N6)? { 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                      (N7)? { 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                      (N8)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                      (N9)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                      (N10)? { 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                      (N11)? { 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                      (N12)? { 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                      (N13)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                      (N14)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N5 = N89;
  assign N6 = N94;
  assign N7 = N100;
  assign N8 = N103;
  assign N9 = N109;
  assign N10 = N112;
  assign N11 = N118;
  assign N12 = N121;
  assign N13 = N128;
  assign N14 = N131;
  assign decode_o[4:0] = (N15)? { N137, N135, N134, N133, N132 } : 
                         (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = opcode_i[5];
  assign N16 = N80;
  assign N44 = N234 | N235;
  assign N234 = N232 | N233;
  assign N232 = N230 | N231;
  assign N230 = N228 | N229;
  assign N228 = N226 | N227;
  assign N226 = N224 | N225;
  assign N224 = N222 | N223;
  assign N222 = N220 | N221;
  assign N220 = N218 | N219;
  assign N218 = N216 | N217;
  assign N216 = N214 | N215;
  assign N214 = ~N21;
  assign N215 = ~N23;
  assign N217 = ~N25;
  assign N219 = ~N28;
  assign N221 = ~N30;
  assign N223 = ~N31;
  assign N225 = ~N32;
  assign N227 = ~N33;
  assign N229 = ~N36;
  assign N231 = ~N39;
  assign N233 = ~N41;
  assign N235 = ~N43;
  assign N61 = N256 | N257;
  assign N256 = N254 | N255;
  assign N254 = N252 | N253;
  assign N252 = N250 | N251;
  assign N250 = N248 | N249;
  assign N248 = N246 | N247;
  assign N246 = N244 | N245;
  assign N244 = N242 | N243;
  assign N242 = N240 | N241;
  assign N240 = N238 | N239;
  assign N238 = N236 | N237;
  assign N236 = ~N47;
  assign N237 = ~N48;
  assign N239 = ~N49;
  assign N241 = ~N51;
  assign N243 = ~N52;
  assign N245 = ~N53;
  assign N247 = ~N54;
  assign N249 = ~N55;
  assign N251 = ~N57;
  assign N253 = ~N58;
  assign N255 = ~N59;
  assign N257 = ~N60;
  assign N65 = N260 | N261;
  assign N260 = N258 | N259;
  assign N258 = ~N62;
  assign N259 = ~N63;
  assign N261 = ~N64;
  assign N73 = N263 | N264;
  assign N263 = N70 | N262;
  assign N262 = ~N71;
  assign N264 = ~N72;
  assign N79 = N75 | N266;
  assign N266 = N76 | N265;
  assign N265 = N77 | N78;
  assign decode_o[17] = N187 | N189;
  assign decode_o[18] = N269 | decode_o[4];
  assign N269 = N268 | N182;
  assign N268 = N267 | N180;
  assign N267 = N175 | N177;
  assign decode_o[16] = N276 | N187;
  assign N276 = N275 | N200;
  assign N275 = N274 | N198;
  assign N274 = N273 | N195;
  assign N273 = N272 | N193;
  assign N272 = N271 | N182;
  assign N271 = N270 | N180;
  assign N270 = N175 | N177;
  assign decode_o[15] = N279 | N189;
  assign N279 = N278 | N211;
  assign N278 = N277 | N209;
  assign N277 = N204 | N206;
  assign decode_o[5] = ~decode_o[14];
  assign N80 = ~opcode_i[5];
  assign N89 = N84 | N280;
  assign N280 = ~N88;
  assign N94 = N281 | N282;
  assign N281 = ~N92;
  assign N282 = ~N93;
  assign N100 = N283 | N284;
  assign N283 = ~N97;
  assign N284 = ~N99;
  assign N103 = N285 | N286;
  assign N285 = ~N101;
  assign N286 = ~N102;
  assign N109 = N287 | N288;
  assign N287 = ~N106;
  assign N288 = ~N108;
  assign N112 = N289 | N290;
  assign N289 = ~N110;
  assign N290 = ~N111;
  assign N118 = N291 | N292;
  assign N291 = ~N115;
  assign N292 = ~N117;
  assign N121 = N293 | N294;
  assign N293 = ~N119;
  assign N294 = ~N120;
  assign N128 = N295 | N296;
  assign N295 = ~N124;
  assign N296 = ~N127;
  assign N131 = N129 | N297;
  assign N297 = N130 | N77;
  assign N136 = ~N131;
  assign N137 = N136;

endmodule



module bsg_mem_1rw_sync_mask_write_bit_000000b0_00000080_1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [175:0] data_i;
  input [6:0] addr_i;
  input [175:0] w_mask_i;
  output [175:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [175:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_mem_1rw_sync_mask_write_byte_00000200_00000400_1
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  addr_i,
  data_i,
  write_mask_i,
  data_o
);

  input [8:0] addr_i;
  input [1023:0] data_i;
  input [127:0] write_mask_i;
  output [1023:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [1023:0] data_o;

  bsg_mem_1rw_sync_mask_write_byte_synth
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .w_i(w_i),
    .addr_i(addr_i),
    .data_i(data_i),
    .write_mask_i(write_mask_i),
    .data_o(data_o)
  );


endmodule



module bsg_mem_1rw_sync_mask_write_bit_00000020_00000080_1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [31:0] data_i;
  input [6:0] addr_i;
  input [31:0] w_mask_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [31:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_scan_00000008_1_1
(
  i,
  o
);

  input [7:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__7_,t_1__6_,
  t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__7_ = i[0] | 1'b0;
  assign t_1__6_ = i[1] | i[0];
  assign t_1__5_ = i[2] | i[1];
  assign t_1__4_ = i[3] | i[2];
  assign t_1__3_ = i[4] | i[3];
  assign t_1__2_ = i[5] | i[4];
  assign t_1__1_ = i[6] | i[5];
  assign t_1__0_ = i[7] | i[6];
  assign t_2__7_ = t_1__7_ | 1'b0;
  assign t_2__6_ = t_1__6_ | 1'b0;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign o[0] = t_2__7_ | 1'b0;
  assign o[1] = t_2__6_ | 1'b0;
  assign o[2] = t_2__5_ | 1'b0;
  assign o[3] = t_2__4_ | 1'b0;
  assign o[4] = t_2__3_ | t_2__7_;
  assign o[5] = t_2__2_ | t_2__6_;
  assign o[6] = t_2__1_ | t_2__5_;
  assign o[7] = t_2__0_ | t_2__4_;

endmodule



module bsg_priority_encode_one_hot_out_00000008_1
(
  i,
  o,
  v_o
);

  input [7:0] i;
  output [7:0] o;
  output v_o;
  wire [7:0] o;
  wire v_o,N0,N1,N2,N3,N4,N5,N6;
  wire [6:1] scan_lo;

  bsg_scan_00000008_1_1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, scan_lo, o[0:0] })
  );

  assign o[7] = v_o & N0;
  assign N0 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N1;
  assign N1 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N2;
  assign N2 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N3;
  assign N3 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N4;
  assign N4 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N5;
  assign N5 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N6;
  assign N6 = ~o[0];

endmodule



module bsg_encode_one_hot_00000008_1
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o,v_2__0_,v_1__6_,v_1__4_,v_1__2_,v_1__0_,addr_2__4_,addr_2__0_;
  assign v_1__0_ = i[1] | i[0];
  assign v_1__2_ = i[3] | i[2];
  assign v_1__4_ = i[5] | i[4];
  assign v_1__6_ = i[7] | i[6];
  assign v_2__0_ = v_1__2_ | v_1__0_;
  assign addr_2__0_ = i[1] | i[3];
  assign addr_o[2] = v_1__6_ | v_1__4_;
  assign addr_2__4_ = i[5] | i[7];
  assign v_o = addr_o[2] | v_2__0_;
  assign addr_o[1] = v_1__2_ | v_1__6_;
  assign addr_o[0] = addr_2__0_ | addr_2__4_;

endmodule



module bsg_priority_encode_00000008_1
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [7:0] enc_lo;

  bsg_priority_encode_one_hot_out_00000008_1
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_00000008_1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o)
  );


endmodule



module bsg_mem_1rw_sync_mask_write_bit_0000000f_00000080_1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [14:0] data_i;
  input [6:0] addr_i;
  input [14:0] w_mask_i;
  output [14:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [14:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_lru_pseudo_tree_decode_00000008
(
  way_id_i,
  data_o,
  mask_o
);

  input [2:0] way_id_i;
  output [6:0] data_o;
  output [6:0] mask_o;
  wire [6:0] data_o,mask_o;
  wire N0,N1,N2;
  assign mask_o[0] = 1'b1;
  assign data_o[0] = 1'b1 & N0;
  assign N0 = ~way_id_i[2];
  assign mask_o[1] = 1'b1 & N0;
  assign data_o[1] = mask_o[1] & N1;
  assign N1 = ~way_id_i[1];
  assign mask_o[2] = 1'b1 & way_id_i[2];
  assign data_o[2] = mask_o[2] & N1;
  assign mask_o[3] = mask_o[1] & N1;
  assign data_o[3] = mask_o[3] & N2;
  assign N2 = ~way_id_i[0];
  assign mask_o[4] = mask_o[1] & way_id_i[1];
  assign data_o[4] = mask_o[4] & N2;
  assign mask_o[5] = mask_o[2] & N1;
  assign data_o[5] = mask_o[5] & N2;
  assign mask_o[6] = mask_o[2] & way_id_i[1];
  assign data_o[6] = mask_o[6] & N2;

endmodule



module bsg_lru_pseudo_tree_backup_00000008
(
  disabled_ways_i,
  modify_mask_o,
  modify_data_o
);

  input [7:0] disabled_ways_i;
  output [6:0] modify_mask_o;
  output [6:0] modify_data_o;
  wire [6:0] modify_mask_o,modify_data_o;
  wire modify_data_o_6_,modify_data_o_5_,modify_data_o_4_,modify_data_o_3_,
  \lru.genblk1_1_.and_reduce_1 ,N0,N1,N2,N3;
  wire [1:1] \lru.genblk1_0_.and_reduce ;
  wire [3:3] \lru.genblk1_1_.and_reduce ;
  assign modify_data_o_6_ = disabled_ways_i[6];
  assign modify_data_o[6] = modify_data_o_6_;
  assign modify_data_o_5_ = disabled_ways_i[4];
  assign modify_data_o[5] = modify_data_o_5_;
  assign modify_data_o_4_ = disabled_ways_i[2];
  assign modify_data_o[4] = modify_data_o_4_;
  assign modify_data_o_3_ = disabled_ways_i[0];
  assign modify_data_o[3] = modify_data_o_3_;
  assign modify_data_o[0] = N1 & modify_data_o_3_;
  assign N1 = N0 & disabled_ways_i[1];
  assign N0 = disabled_ways_i[3] & modify_data_o_4_;
  assign \lru.genblk1_0_.and_reduce [1] = N3 & modify_data_o_5_;
  assign N3 = N2 & disabled_ways_i[5];
  assign N2 = disabled_ways_i[7] & modify_data_o_6_;
  assign modify_mask_o[0] = \lru.genblk1_0_.and_reduce [1] | modify_data_o[0];
  assign modify_data_o[1] = disabled_ways_i[1] & modify_data_o_3_;
  assign \lru.genblk1_1_.and_reduce_1  = disabled_ways_i[3] & modify_data_o_4_;
  assign modify_data_o[2] = disabled_ways_i[5] & modify_data_o_5_;
  assign \lru.genblk1_1_.and_reduce [3] = disabled_ways_i[7] & modify_data_o_6_;
  assign modify_mask_o[1] = \lru.genblk1_1_.and_reduce_1  | modify_data_o[1];
  assign modify_mask_o[2] = \lru.genblk1_1_.and_reduce [3] | modify_data_o[2];
  assign modify_mask_o[3] = disabled_ways_i[1] | modify_data_o_3_;
  assign modify_mask_o[4] = disabled_ways_i[3] | modify_data_o_4_;
  assign modify_mask_o[5] = disabled_ways_i[5] | modify_data_o_5_;
  assign modify_mask_o[6] = disabled_ways_i[7] | modify_data_o_6_;

endmodule



module bsg_mux_segmented_00000007_1
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [6:0] data0_i;
  input [6:0] data1_i;
  input [6:0] sel_i;
  output [6:0] data_o;
  wire [6:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;
  assign data_o[0] = (N0)? data1_i[0] : 
                     (N7)? data0_i[0] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[1] = (N1)? data1_i[1] : 
                     (N8)? data0_i[1] : 1'b0;
  assign N1 = sel_i[1];
  assign data_o[2] = (N2)? data1_i[2] : 
                     (N9)? data0_i[2] : 1'b0;
  assign N2 = sel_i[2];
  assign data_o[3] = (N3)? data1_i[3] : 
                     (N10)? data0_i[3] : 1'b0;
  assign N3 = sel_i[3];
  assign data_o[4] = (N4)? data1_i[4] : 
                     (N11)? data0_i[4] : 1'b0;
  assign N4 = sel_i[4];
  assign data_o[5] = (N5)? data1_i[5] : 
                     (N12)? data0_i[5] : 1'b0;
  assign N5 = sel_i[5];
  assign data_o[6] = (N6)? data1_i[6] : 
                     (N13)? data0_i[6] : 1'b0;
  assign N6 = sel_i[6];
  assign N7 = ~sel_i[0];
  assign N8 = ~sel_i[1];
  assign N9 = ~sel_i[2];
  assign N10 = ~sel_i[3];
  assign N11 = ~sel_i[4];
  assign N12 = ~sel_i[5];
  assign N13 = ~sel_i[6];

endmodule



module bsg_mux_bitwise_00000007
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [6:0] data0_i;
  input [6:0] data1_i;
  input [6:0] sel_i;
  output [6:0] data_o;
  wire [6:0] data_o;

  bsg_mux_segmented_00000007_1
  mux_segmented
  (
    .data0_i(data0_i),
    .data1_i(data1_i),
    .sel_i(sel_i),
    .data_o(data_o)
  );


endmodule



module bsg_mux_width_p1_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [1:0] data_i;
  input [0:0] sel_i;
  output [0:0] data_o;
  wire [0:0] data_o;
  wire N0,N1;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[1] : 1'b0;
  assign N0 = sel_i[0];
  assign N1 = ~sel_i[0];

endmodule



module bsg_mux_00000001_00000004
(
  data_i,
  sel_i,
  data_o
);

  input [3:0] data_i;
  input [1:0] sel_i;
  output [0:0] data_o;
  wire [0:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[1] : 
                     (N3)? data_i[2] : 
                     (N5)? data_i[3] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_lru_pseudo_tree_encode_00000008
(
  lru_i,
  way_id_o
);

  input [6:0] lru_i;
  output [2:0] way_id_o;
  wire [2:0] way_id_o;
  wire way_id_o_2_;
  assign way_id_o_2_ = lru_i[0];
  assign way_id_o[2] = way_id_o_2_;

  bsg_mux_width_p1_els_p2
  \lru.rank_1_.nz.mux 
  (
    .data_i(lru_i[2:1]),
    .sel_i(way_id_o_2_),
    .data_o(way_id_o[1])
  );


  bsg_mux_00000001_00000004
  \lru.rank_2_.nz.mux 
  (
    .data_i(lru_i[6:3]),
    .sel_i({ way_id_o_2_, way_id_o[1:1] }),
    .data_o(way_id_o[0])
  );


endmodule



module bsg_decode_00000008
(
  i,
  o
);

  input [2:0] i;
  output [7:0] o;
  wire [7:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_cache_miss_00000021_00000080_00000004_00000080_00000008_1
(
  clk_i,
  reset_i,
  miss_v_i,
  track_miss_i,
  decode_v_i,
  addr_v_i,
  mask_v_i,
  tag_v_i,
  valid_v_i,
  lock_v_i,
  tag_hit_v_i,
  tag_hit_way_id_i,
  tag_hit_found_i,
  sbuf_empty_i,
  tbuf_empty_i,
  dma_cmd_o,
  dma_way_o,
  dma_addr_o,
  dma_done_i,
  track_data_we_o,
  stat_info_i,
  stat_mem_v_o,
  stat_mem_w_o,
  stat_mem_addr_o,
  stat_mem_data_o,
  stat_mem_w_mask_o,
  tag_mem_v_o,
  tag_mem_w_o,
  tag_mem_addr_o,
  tag_mem_data_o,
  tag_mem_w_mask_o,
  track_mem_v_o,
  track_mem_w_o,
  track_mem_addr_o,
  track_mem_w_mask_o,
  track_mem_data_o,
  done_o,
  recover_o,
  chosen_way_o,
  select_snoop_data_r_o,
  ack_i
);

  input [20:0] decode_v_i;
  input [32:0] addr_v_i;
  input [15:0] mask_v_i;
  input [159:0] tag_v_i;
  input [7:0] valid_v_i;
  input [7:0] lock_v_i;
  input [7:0] tag_hit_v_i;
  input [2:0] tag_hit_way_id_i;
  output [3:0] dma_cmd_o;
  output [2:0] dma_way_o;
  output [32:0] dma_addr_o;
  input [14:0] stat_info_i;
  output [6:0] stat_mem_addr_o;
  output [14:0] stat_mem_data_o;
  output [14:0] stat_mem_w_mask_o;
  output [6:0] tag_mem_addr_o;
  output [175:0] tag_mem_data_o;
  output [175:0] tag_mem_w_mask_o;
  output [6:0] track_mem_addr_o;
  output [31:0] track_mem_w_mask_o;
  output [31:0] track_mem_data_o;
  output [2:0] chosen_way_o;
  input clk_i;
  input reset_i;
  input miss_v_i;
  input track_miss_i;
  input tag_hit_found_i;
  input sbuf_empty_i;
  input tbuf_empty_i;
  input dma_done_i;
  input ack_i;
  output track_data_we_o;
  output stat_mem_v_o;
  output stat_mem_w_o;
  output tag_mem_v_o;
  output tag_mem_w_o;
  output track_mem_v_o;
  output track_mem_w_o;
  output done_o;
  output recover_o;
  output select_snoop_data_r_o;
  wire [3:0] dma_cmd_o,miss_state_r,miss_state_n;
  wire [2:0] dma_way_o,chosen_way_o,invalid_way_id,flush_way_r,lru_way_id,chosen_way_n;
  wire [32:0] dma_addr_o;
  wire [6:0] stat_mem_addr_o,tag_mem_addr_o,track_mem_addr_o,chosen_way_lru_data,
  chosen_way_lru_mask,modify_mask_lo,modify_data_lo,modified_lru_bits;
  wire [14:0] stat_mem_data_o,stat_mem_w_mask_o;
  wire [175:0] tag_mem_data_o,tag_mem_w_mask_o;
  wire [31:0] track_mem_w_mask_o,track_mem_data_o;
  wire track_data_we_o,stat_mem_v_o,stat_mem_w_o,tag_mem_v_o,tag_mem_w_o,track_mem_v_o,
  track_mem_w_o,done_o,recover_o,select_snoop_data_r_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,
  N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,track_mem_data_o_7__3_,
  _0_net__7_,_0_net__6_,_0_net__5_,_0_net__4_,_0_net__3_,_0_net__2_,_0_net__1_,
  _0_net__0_,invalid_exist,goto_flush_op,goto_lock_op,N23,N24,full_word_op,
  st_tag_miss_op,N25,N26,select_snoop_data_n,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,
  N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,
  N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,
  N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,
  N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,
  N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
  N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,
  N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,
  N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,
  N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,
  N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,
  N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,
  N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
  N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,
  N355;
  wire [7:0] chosen_way_decode,addr_way_v_decode,flush_way_decode;
  reg track_data_we_o_sv2v_reg,miss_state_r_3_sv2v_reg,miss_state_r_2_sv2v_reg,
  miss_state_r_1_sv2v_reg,miss_state_r_0_sv2v_reg,chosen_way_o_2_sv2v_reg,
  chosen_way_o_1_sv2v_reg,chosen_way_o_0_sv2v_reg,flush_way_r_2_sv2v_reg,flush_way_r_1_sv2v_reg,
  flush_way_r_0_sv2v_reg,select_snoop_data_r_o_sv2v_reg;
  assign track_data_we_o = track_data_we_o_sv2v_reg;
  assign miss_state_r[3] = miss_state_r_3_sv2v_reg;
  assign miss_state_r[2] = miss_state_r_2_sv2v_reg;
  assign miss_state_r[1] = miss_state_r_1_sv2v_reg;
  assign miss_state_r[0] = miss_state_r_0_sv2v_reg;
  assign chosen_way_o[2] = chosen_way_o_2_sv2v_reg;
  assign chosen_way_o[1] = chosen_way_o_1_sv2v_reg;
  assign chosen_way_o[0] = chosen_way_o_0_sv2v_reg;
  assign flush_way_r[2] = flush_way_r_2_sv2v_reg;
  assign flush_way_r[1] = flush_way_r_1_sv2v_reg;
  assign flush_way_r[0] = flush_way_r_0_sv2v_reg;
  assign select_snoop_data_r_o = select_snoop_data_r_o_sv2v_reg;
  assign dma_addr_o[0] = 1'b0;
  assign dma_addr_o[1] = 1'b0;
  assign dma_addr_o[2] = 1'b0;
  assign dma_addr_o[3] = 1'b0;
  assign stat_mem_addr_o[6] = addr_v_i[12];
  assign track_mem_addr_o[6] = stat_mem_addr_o[6];
  assign tag_mem_addr_o[6] = stat_mem_addr_o[6];
  assign stat_mem_addr_o[5] = addr_v_i[11];
  assign track_mem_addr_o[5] = stat_mem_addr_o[5];
  assign tag_mem_addr_o[5] = stat_mem_addr_o[5];
  assign stat_mem_addr_o[4] = addr_v_i[10];
  assign track_mem_addr_o[4] = stat_mem_addr_o[4];
  assign tag_mem_addr_o[4] = stat_mem_addr_o[4];
  assign stat_mem_addr_o[3] = addr_v_i[9];
  assign track_mem_addr_o[3] = stat_mem_addr_o[3];
  assign tag_mem_addr_o[3] = stat_mem_addr_o[3];
  assign stat_mem_addr_o[2] = addr_v_i[8];
  assign track_mem_addr_o[2] = stat_mem_addr_o[2];
  assign tag_mem_addr_o[2] = stat_mem_addr_o[2];
  assign stat_mem_addr_o[1] = addr_v_i[7];
  assign track_mem_addr_o[1] = stat_mem_addr_o[1];
  assign tag_mem_addr_o[1] = stat_mem_addr_o[1];
  assign stat_mem_addr_o[0] = addr_v_i[6];
  assign track_mem_addr_o[0] = stat_mem_addr_o[0];
  assign tag_mem_addr_o[0] = stat_mem_addr_o[0];
  assign dma_cmd_o[2] = track_mem_data_o_7__3_;
  assign track_mem_data_o[0] = track_mem_data_o_7__3_;
  assign track_mem_data_o[1] = track_mem_data_o_7__3_;
  assign track_mem_data_o[2] = track_mem_data_o_7__3_;
  assign track_mem_data_o[3] = track_mem_data_o_7__3_;
  assign track_mem_data_o[4] = track_mem_data_o_7__3_;
  assign track_mem_data_o[5] = track_mem_data_o_7__3_;
  assign track_mem_data_o[6] = track_mem_data_o_7__3_;
  assign track_mem_data_o[7] = track_mem_data_o_7__3_;
  assign track_mem_data_o[8] = track_mem_data_o_7__3_;
  assign track_mem_data_o[9] = track_mem_data_o_7__3_;
  assign track_mem_data_o[10] = track_mem_data_o_7__3_;
  assign track_mem_data_o[11] = track_mem_data_o_7__3_;
  assign track_mem_data_o[12] = track_mem_data_o_7__3_;
  assign track_mem_data_o[13] = track_mem_data_o_7__3_;
  assign track_mem_data_o[14] = track_mem_data_o_7__3_;
  assign track_mem_data_o[15] = track_mem_data_o_7__3_;
  assign track_mem_data_o[16] = track_mem_data_o_7__3_;
  assign track_mem_data_o[17] = track_mem_data_o_7__3_;
  assign track_mem_data_o[18] = track_mem_data_o_7__3_;
  assign track_mem_data_o[19] = track_mem_data_o_7__3_;
  assign track_mem_data_o[20] = track_mem_data_o_7__3_;
  assign track_mem_data_o[21] = track_mem_data_o_7__3_;
  assign track_mem_data_o[22] = track_mem_data_o_7__3_;
  assign track_mem_data_o[23] = track_mem_data_o_7__3_;
  assign track_mem_data_o[24] = track_mem_data_o_7__3_;
  assign track_mem_data_o[25] = track_mem_data_o_7__3_;
  assign track_mem_data_o[26] = track_mem_data_o_7__3_;
  assign track_mem_data_o[27] = track_mem_data_o_7__3_;
  assign track_mem_data_o[28] = track_mem_data_o_7__3_;
  assign track_mem_data_o[29] = track_mem_data_o_7__3_;
  assign track_mem_data_o[30] = track_mem_data_o_7__3_;
  assign track_mem_data_o[31] = track_mem_data_o_7__3_;

  bsg_priority_encode_00000008_1
  invalid_way_pe
  (
    .i({ _0_net__7_, _0_net__6_, _0_net__5_, _0_net__4_, _0_net__3_, _0_net__2_, _0_net__1_, _0_net__0_ }),
    .addr_o(invalid_way_id),
    .v_o(invalid_exist)
  );


  bsg_lru_pseudo_tree_decode_00000008
  chosen_way_lru_decode
  (
    .way_id_i(chosen_way_o),
    .data_o(chosen_way_lru_data),
    .mask_o(chosen_way_lru_mask)
  );


  bsg_lru_pseudo_tree_backup_00000008
  backup_lru
  (
    .disabled_ways_i(lock_v_i),
    .modify_mask_o(modify_mask_lo),
    .modify_data_o(modify_data_lo)
  );


  bsg_mux_bitwise_00000007
  lru_bit_mux
  (
    .data0_i(stat_info_i[6:0]),
    .data1_i(modify_data_lo),
    .sel_i(modify_mask_lo),
    .data_o(modified_lru_bits)
  );


  bsg_lru_pseudo_tree_encode_00000008
  lru_encode
  (
    .lru_i(modified_lru_bits),
    .way_id_o(lru_way_id)
  );


  bsg_decode_00000008
  chosen_way_demux
  (
    .i(chosen_way_n),
    .o(chosen_way_decode)
  );


  bsg_decode_00000008
  addr_way_v_demux
  (
    .i(addr_v_i[15:13]),
    .o(addr_way_v_decode)
  );

  assign N31 = N27 & N28;
  assign N32 = N29 & N30;
  assign N33 = N31 & N32;
  assign N34 = miss_state_r[3] | N28;
  assign N35 = miss_state_r[1] | miss_state_r[0];
  assign N36 = N34 | N35;
  assign N38 = miss_state_r[3] | miss_state_r[2];
  assign N39 = miss_state_r[1] | N30;
  assign N40 = N38 | N39;
  assign N42 = miss_state_r[3] | miss_state_r[2];
  assign N43 = N29 | miss_state_r[0];
  assign N44 = N42 | N43;
  assign N46 = miss_state_r[3] | miss_state_r[2];
  assign N47 = N29 | N30;
  assign N48 = N46 | N47;
  assign N50 = miss_state_r[3] | N28;
  assign N51 = miss_state_r[1] | N30;
  assign N52 = N50 | N51;
  assign N54 = miss_state_r[3] | N28;
  assign N55 = N29 | miss_state_r[0];
  assign N56 = N54 | N55;
  assign N58 = miss_state_r[3] | N28;
  assign N59 = N29 | N30;
  assign N60 = N58 | N59;
  assign N62 = N27 | miss_state_r[2];
  assign N63 = miss_state_r[1] | miss_state_r[0];
  assign N64 = N62 | N63;
  assign N66 = N27 | miss_state_r[2];
  assign N67 = miss_state_r[1] | N30;
  assign N68 = N66 | N67;
  assign N70 = N27 | miss_state_r[2];
  assign N71 = N29 | miss_state_r[0];
  assign N72 = N70 | N71;
  assign N74 = miss_state_r[3] & miss_state_r[1];
  assign N75 = N74 & miss_state_r[0];
  assign N76 = miss_state_r[3] & miss_state_r[2];
  assign N109 = (N101)? stat_info_i[7] : 
                (N103)? stat_info_i[8] : 
                (N105)? stat_info_i[9] : 
                (N107)? stat_info_i[10] : 
                (N102)? stat_info_i[11] : 
                (N104)? stat_info_i[12] : 
                (N106)? stat_info_i[13] : 
                (N108)? stat_info_i[14] : 1'b0;
  assign N110 = (N101)? valid_v_i[0] : 
                (N103)? valid_v_i[1] : 
                (N105)? valid_v_i[2] : 
                (N107)? valid_v_i[3] : 
                (N102)? valid_v_i[4] : 
                (N104)? valid_v_i[5] : 
                (N106)? valid_v_i[6] : 
                (N108)? valid_v_i[7] : 1'b0;
  assign N149 = (N141)? stat_info_i[7] : 
                (N143)? stat_info_i[8] : 
                (N145)? stat_info_i[9] : 
                (N147)? stat_info_i[10] : 
                (N142)? stat_info_i[11] : 
                (N144)? stat_info_i[12] : 
                (N146)? stat_info_i[13] : 
                (N148)? stat_info_i[14] : 1'b0;
  assign N150 = (N141)? valid_v_i[0] : 
                (N143)? valid_v_i[1] : 
                (N145)? valid_v_i[2] : 
                (N147)? valid_v_i[3] : 
                (N142)? valid_v_i[4] : 
                (N144)? valid_v_i[5] : 
                (N146)? valid_v_i[6] : 
                (N148)? valid_v_i[7] : 1'b0;
  assign N168 = (N160)? tag_v_i[19] : 
                (N162)? tag_v_i[39] : 
                (N164)? tag_v_i[59] : 
                (N166)? tag_v_i[79] : 
                (N161)? tag_v_i[99] : 
                (N163)? tag_v_i[119] : 
                (N165)? tag_v_i[139] : 
                (N167)? tag_v_i[159] : 1'b0;
  assign N169 = (N160)? tag_v_i[18] : 
                (N162)? tag_v_i[38] : 
                (N164)? tag_v_i[58] : 
                (N166)? tag_v_i[78] : 
                (N161)? tag_v_i[98] : 
                (N163)? tag_v_i[118] : 
                (N165)? tag_v_i[138] : 
                (N167)? tag_v_i[158] : 1'b0;
  assign N170 = (N160)? tag_v_i[17] : 
                (N162)? tag_v_i[37] : 
                (N164)? tag_v_i[57] : 
                (N166)? tag_v_i[77] : 
                (N161)? tag_v_i[97] : 
                (N163)? tag_v_i[117] : 
                (N165)? tag_v_i[137] : 
                (N167)? tag_v_i[157] : 1'b0;
  assign N171 = (N160)? tag_v_i[16] : 
                (N162)? tag_v_i[36] : 
                (N164)? tag_v_i[56] : 
                (N166)? tag_v_i[76] : 
                (N161)? tag_v_i[96] : 
                (N163)? tag_v_i[116] : 
                (N165)? tag_v_i[136] : 
                (N167)? tag_v_i[156] : 1'b0;
  assign N172 = (N160)? tag_v_i[15] : 
                (N162)? tag_v_i[35] : 
                (N164)? tag_v_i[55] : 
                (N166)? tag_v_i[75] : 
                (N161)? tag_v_i[95] : 
                (N163)? tag_v_i[115] : 
                (N165)? tag_v_i[135] : 
                (N167)? tag_v_i[155] : 1'b0;
  assign N173 = (N160)? tag_v_i[14] : 
                (N162)? tag_v_i[34] : 
                (N164)? tag_v_i[54] : 
                (N166)? tag_v_i[74] : 
                (N161)? tag_v_i[94] : 
                (N163)? tag_v_i[114] : 
                (N165)? tag_v_i[134] : 
                (N167)? tag_v_i[154] : 1'b0;
  assign N174 = (N160)? tag_v_i[13] : 
                (N162)? tag_v_i[33] : 
                (N164)? tag_v_i[53] : 
                (N166)? tag_v_i[73] : 
                (N161)? tag_v_i[93] : 
                (N163)? tag_v_i[113] : 
                (N165)? tag_v_i[133] : 
                (N167)? tag_v_i[153] : 1'b0;
  assign N175 = (N160)? tag_v_i[12] : 
                (N162)? tag_v_i[32] : 
                (N164)? tag_v_i[52] : 
                (N166)? tag_v_i[72] : 
                (N161)? tag_v_i[92] : 
                (N163)? tag_v_i[112] : 
                (N165)? tag_v_i[132] : 
                (N167)? tag_v_i[152] : 1'b0;
  assign N176 = (N160)? tag_v_i[11] : 
                (N162)? tag_v_i[31] : 
                (N164)? tag_v_i[51] : 
                (N166)? tag_v_i[71] : 
                (N161)? tag_v_i[91] : 
                (N163)? tag_v_i[111] : 
                (N165)? tag_v_i[131] : 
                (N167)? tag_v_i[151] : 1'b0;
  assign N177 = (N160)? tag_v_i[10] : 
                (N162)? tag_v_i[30] : 
                (N164)? tag_v_i[50] : 
                (N166)? tag_v_i[70] : 
                (N161)? tag_v_i[90] : 
                (N163)? tag_v_i[110] : 
                (N165)? tag_v_i[130] : 
                (N167)? tag_v_i[150] : 1'b0;
  assign N178 = (N160)? tag_v_i[9] : 
                (N162)? tag_v_i[29] : 
                (N164)? tag_v_i[49] : 
                (N166)? tag_v_i[69] : 
                (N161)? tag_v_i[89] : 
                (N163)? tag_v_i[109] : 
                (N165)? tag_v_i[129] : 
                (N167)? tag_v_i[149] : 1'b0;
  assign N179 = (N160)? tag_v_i[8] : 
                (N162)? tag_v_i[28] : 
                (N164)? tag_v_i[48] : 
                (N166)? tag_v_i[68] : 
                (N161)? tag_v_i[88] : 
                (N163)? tag_v_i[108] : 
                (N165)? tag_v_i[128] : 
                (N167)? tag_v_i[148] : 1'b0;
  assign N180 = (N160)? tag_v_i[7] : 
                (N162)? tag_v_i[27] : 
                (N164)? tag_v_i[47] : 
                (N166)? tag_v_i[67] : 
                (N161)? tag_v_i[87] : 
                (N163)? tag_v_i[107] : 
                (N165)? tag_v_i[127] : 
                (N167)? tag_v_i[147] : 1'b0;
  assign N181 = (N160)? tag_v_i[6] : 
                (N162)? tag_v_i[26] : 
                (N164)? tag_v_i[46] : 
                (N166)? tag_v_i[66] : 
                (N161)? tag_v_i[86] : 
                (N163)? tag_v_i[106] : 
                (N165)? tag_v_i[126] : 
                (N167)? tag_v_i[146] : 1'b0;
  assign N182 = (N160)? tag_v_i[5] : 
                (N162)? tag_v_i[25] : 
                (N164)? tag_v_i[45] : 
                (N166)? tag_v_i[65] : 
                (N161)? tag_v_i[85] : 
                (N163)? tag_v_i[105] : 
                (N165)? tag_v_i[125] : 
                (N167)? tag_v_i[145] : 1'b0;
  assign N183 = (N160)? tag_v_i[4] : 
                (N162)? tag_v_i[24] : 
                (N164)? tag_v_i[44] : 
                (N166)? tag_v_i[64] : 
                (N161)? tag_v_i[84] : 
                (N163)? tag_v_i[104] : 
                (N165)? tag_v_i[124] : 
                (N167)? tag_v_i[144] : 1'b0;
  assign N184 = (N160)? tag_v_i[3] : 
                (N162)? tag_v_i[23] : 
                (N164)? tag_v_i[43] : 
                (N166)? tag_v_i[63] : 
                (N161)? tag_v_i[83] : 
                (N163)? tag_v_i[103] : 
                (N165)? tag_v_i[123] : 
                (N167)? tag_v_i[143] : 1'b0;
  assign N185 = (N160)? tag_v_i[2] : 
                (N162)? tag_v_i[22] : 
                (N164)? tag_v_i[42] : 
                (N166)? tag_v_i[62] : 
                (N161)? tag_v_i[82] : 
                (N163)? tag_v_i[102] : 
                (N165)? tag_v_i[122] : 
                (N167)? tag_v_i[142] : 1'b0;
  assign N186 = (N160)? tag_v_i[1] : 
                (N162)? tag_v_i[21] : 
                (N164)? tag_v_i[41] : 
                (N166)? tag_v_i[61] : 
                (N161)? tag_v_i[81] : 
                (N163)? tag_v_i[101] : 
                (N165)? tag_v_i[121] : 
                (N167)? tag_v_i[141] : 1'b0;
  assign N187 = (N160)? tag_v_i[0] : 
                (N162)? tag_v_i[20] : 
                (N164)? tag_v_i[40] : 
                (N166)? tag_v_i[60] : 
                (N161)? tag_v_i[80] : 
                (N163)? tag_v_i[100] : 
                (N165)? tag_v_i[120] : 
                (N167)? tag_v_i[140] : 1'b0;
  assign N201 = (N193)? tag_v_i[19] : 
                (N195)? tag_v_i[39] : 
                (N197)? tag_v_i[59] : 
                (N199)? tag_v_i[79] : 
                (N194)? tag_v_i[99] : 
                (N196)? tag_v_i[119] : 
                (N198)? tag_v_i[139] : 
                (N200)? tag_v_i[159] : 1'b0;
  assign N202 = (N193)? tag_v_i[18] : 
                (N195)? tag_v_i[38] : 
                (N197)? tag_v_i[58] : 
                (N199)? tag_v_i[78] : 
                (N194)? tag_v_i[98] : 
                (N196)? tag_v_i[118] : 
                (N198)? tag_v_i[138] : 
                (N200)? tag_v_i[158] : 1'b0;
  assign N203 = (N193)? tag_v_i[17] : 
                (N195)? tag_v_i[37] : 
                (N197)? tag_v_i[57] : 
                (N199)? tag_v_i[77] : 
                (N194)? tag_v_i[97] : 
                (N196)? tag_v_i[117] : 
                (N198)? tag_v_i[137] : 
                (N200)? tag_v_i[157] : 1'b0;
  assign N204 = (N193)? tag_v_i[16] : 
                (N195)? tag_v_i[36] : 
                (N197)? tag_v_i[56] : 
                (N199)? tag_v_i[76] : 
                (N194)? tag_v_i[96] : 
                (N196)? tag_v_i[116] : 
                (N198)? tag_v_i[136] : 
                (N200)? tag_v_i[156] : 1'b0;
  assign N205 = (N193)? tag_v_i[15] : 
                (N195)? tag_v_i[35] : 
                (N197)? tag_v_i[55] : 
                (N199)? tag_v_i[75] : 
                (N194)? tag_v_i[95] : 
                (N196)? tag_v_i[115] : 
                (N198)? tag_v_i[135] : 
                (N200)? tag_v_i[155] : 1'b0;
  assign N206 = (N193)? tag_v_i[14] : 
                (N195)? tag_v_i[34] : 
                (N197)? tag_v_i[54] : 
                (N199)? tag_v_i[74] : 
                (N194)? tag_v_i[94] : 
                (N196)? tag_v_i[114] : 
                (N198)? tag_v_i[134] : 
                (N200)? tag_v_i[154] : 1'b0;
  assign N207 = (N193)? tag_v_i[13] : 
                (N195)? tag_v_i[33] : 
                (N197)? tag_v_i[53] : 
                (N199)? tag_v_i[73] : 
                (N194)? tag_v_i[93] : 
                (N196)? tag_v_i[113] : 
                (N198)? tag_v_i[133] : 
                (N200)? tag_v_i[153] : 1'b0;
  assign N208 = (N193)? tag_v_i[12] : 
                (N195)? tag_v_i[32] : 
                (N197)? tag_v_i[52] : 
                (N199)? tag_v_i[72] : 
                (N194)? tag_v_i[92] : 
                (N196)? tag_v_i[112] : 
                (N198)? tag_v_i[132] : 
                (N200)? tag_v_i[152] : 1'b0;
  assign N209 = (N193)? tag_v_i[11] : 
                (N195)? tag_v_i[31] : 
                (N197)? tag_v_i[51] : 
                (N199)? tag_v_i[71] : 
                (N194)? tag_v_i[91] : 
                (N196)? tag_v_i[111] : 
                (N198)? tag_v_i[131] : 
                (N200)? tag_v_i[151] : 1'b0;
  assign N210 = (N193)? tag_v_i[10] : 
                (N195)? tag_v_i[30] : 
                (N197)? tag_v_i[50] : 
                (N199)? tag_v_i[70] : 
                (N194)? tag_v_i[90] : 
                (N196)? tag_v_i[110] : 
                (N198)? tag_v_i[130] : 
                (N200)? tag_v_i[150] : 1'b0;
  assign N211 = (N193)? tag_v_i[9] : 
                (N195)? tag_v_i[29] : 
                (N197)? tag_v_i[49] : 
                (N199)? tag_v_i[69] : 
                (N194)? tag_v_i[89] : 
                (N196)? tag_v_i[109] : 
                (N198)? tag_v_i[129] : 
                (N200)? tag_v_i[149] : 1'b0;
  assign N212 = (N193)? tag_v_i[8] : 
                (N195)? tag_v_i[28] : 
                (N197)? tag_v_i[48] : 
                (N199)? tag_v_i[68] : 
                (N194)? tag_v_i[88] : 
                (N196)? tag_v_i[108] : 
                (N198)? tag_v_i[128] : 
                (N200)? tag_v_i[148] : 1'b0;
  assign N213 = (N193)? tag_v_i[7] : 
                (N195)? tag_v_i[27] : 
                (N197)? tag_v_i[47] : 
                (N199)? tag_v_i[67] : 
                (N194)? tag_v_i[87] : 
                (N196)? tag_v_i[107] : 
                (N198)? tag_v_i[127] : 
                (N200)? tag_v_i[147] : 1'b0;
  assign N214 = (N193)? tag_v_i[6] : 
                (N195)? tag_v_i[26] : 
                (N197)? tag_v_i[46] : 
                (N199)? tag_v_i[66] : 
                (N194)? tag_v_i[86] : 
                (N196)? tag_v_i[106] : 
                (N198)? tag_v_i[126] : 
                (N200)? tag_v_i[146] : 1'b0;
  assign N215 = (N193)? tag_v_i[5] : 
                (N195)? tag_v_i[25] : 
                (N197)? tag_v_i[45] : 
                (N199)? tag_v_i[65] : 
                (N194)? tag_v_i[85] : 
                (N196)? tag_v_i[105] : 
                (N198)? tag_v_i[125] : 
                (N200)? tag_v_i[145] : 1'b0;
  assign N216 = (N193)? tag_v_i[4] : 
                (N195)? tag_v_i[24] : 
                (N197)? tag_v_i[44] : 
                (N199)? tag_v_i[64] : 
                (N194)? tag_v_i[84] : 
                (N196)? tag_v_i[104] : 
                (N198)? tag_v_i[124] : 
                (N200)? tag_v_i[144] : 1'b0;
  assign N217 = (N193)? tag_v_i[3] : 
                (N195)? tag_v_i[23] : 
                (N197)? tag_v_i[43] : 
                (N199)? tag_v_i[63] : 
                (N194)? tag_v_i[83] : 
                (N196)? tag_v_i[103] : 
                (N198)? tag_v_i[123] : 
                (N200)? tag_v_i[143] : 1'b0;
  assign N218 = (N193)? tag_v_i[2] : 
                (N195)? tag_v_i[22] : 
                (N197)? tag_v_i[42] : 
                (N199)? tag_v_i[62] : 
                (N194)? tag_v_i[82] : 
                (N196)? tag_v_i[102] : 
                (N198)? tag_v_i[122] : 
                (N200)? tag_v_i[142] : 1'b0;
  assign N219 = (N193)? tag_v_i[1] : 
                (N195)? tag_v_i[21] : 
                (N197)? tag_v_i[41] : 
                (N199)? tag_v_i[61] : 
                (N194)? tag_v_i[81] : 
                (N196)? tag_v_i[101] : 
                (N198)? tag_v_i[121] : 
                (N200)? tag_v_i[141] : 1'b0;
  assign N220 = (N193)? tag_v_i[0] : 
                (N195)? tag_v_i[20] : 
                (N197)? tag_v_i[40] : 
                (N199)? tag_v_i[60] : 
                (N194)? tag_v_i[80] : 
                (N196)? tag_v_i[100] : 
                (N198)? tag_v_i[120] : 
                (N200)? tag_v_i[140] : 1'b0;
  assign N258 = (N250)? stat_info_i[7] : 
                (N252)? stat_info_i[8] : 
                (N254)? stat_info_i[9] : 
                (N256)? stat_info_i[10] : 
                (N251)? stat_info_i[11] : 
                (N253)? stat_info_i[12] : 
                (N255)? stat_info_i[13] : 
                (N257)? stat_info_i[14] : 1'b0;
  assign N259 = (N250)? valid_v_i[0] : 
                (N252)? valid_v_i[1] : 
                (N254)? valid_v_i[2] : 
                (N256)? valid_v_i[3] : 
                (N251)? valid_v_i[4] : 
                (N253)? valid_v_i[5] : 
                (N255)? valid_v_i[6] : 
                (N257)? valid_v_i[7] : 1'b0;
  assign full_word_op = (N0)? N24 : 
                        (N23)? 1'b0 : 1'b0;
  assign N0 = decode_v_i[17];
  assign dma_way_o = (N1)? flush_way_r : 
                     (N2)? chosen_way_o : 1'b0;
  assign N1 = goto_flush_op;
  assign N2 = N25;
  assign flush_way_decode = (N3)? addr_way_v_decode : 
                            (N26)? tag_hit_v_i : 1'b0;
  assign N3 = decode_v_i[13];
  assign { N85, N84, N83 } = (N1)? { 1'b0, 1'b0, 1'b1 } : 
                             (N266)? { 1'b0, 1'b1, 1'b0 } : 
                             (N269)? { 1'b1, 1'b1, 1'b1 } : 
                             (N82)? { 1'b1, 1'b0, 1'b0 } : 1'b0;
  assign { N88, N87, N86 } = (N4)? { N85, N84, N83 } : 
                             (N79)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N4 = N78;
  assign { N93, N92, N91 } = (N5)? tag_hit_way_id_i : 
                             (N271)? invalid_way_id : 
                             (N90)? lru_way_id : 1'b0;
  assign N5 = track_miss_i;
  assign N112 = ~N111;
  assign { N114, N113 } = (N6)? { N112, N111 } : 
                          (N7)? { 1'b1, 1'b0 } : 1'b0;
  assign N6 = dma_done_i;
  assign N7 = N188;
  assign { N117, N116, N115 } = (N3)? addr_v_i[15:13] : 
                                (N26)? tag_hit_way_id_i : 1'b0;
  assign N152 = ~N151;
  assign N225 = ~N224;
  assign { N229, N228, N227, N226 } = (N6)? { N224, N225, N225, N224 } : 
                                      (N7)? { 1'b0, 1'b1, 1'b0, 1'b1 } : 1'b0;
  assign { N238, N237, N236, N235, N234, N233, N232, N231 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                              (N8)? chosen_way_decode : 1'b0;
  assign N8 = N333;
  assign { N242, N241, N240 } = (N9)? invalid_way_id : 
                                (N10)? lru_way_id : 1'b0;
  assign N9 = invalid_exist;
  assign N10 = N239;
  assign N261 = ~N260;
  assign stat_mem_v_o = (N11)? N78 : 
                        (N12)? 1'b0 : 
                        (N13)? 1'b1 : 
                        (N14)? 1'b0 : 
                        (N15)? 1'b0 : 
                        (N16)? N221 : 
                        (N17)? dma_done_i : 
                        (N18)? 1'b0 : 
                        (N19)? 1'b1 : 
                        (N20)? 1'b0 : 
                        (N21)? 1'b0 : 
                        (N22)? 1'b0 : 1'b0;
  assign N11 = N33;
  assign N12 = dma_cmd_o[0];
  assign N13 = N41;
  assign N14 = N45;
  assign N15 = dma_cmd_o[1];
  assign N16 = dma_cmd_o[3];
  assign N17 = track_mem_data_o_7__3_;
  assign N18 = N61;
  assign N19 = N65;
  assign N20 = N69;
  assign N21 = N73;
  assign N22 = N77;
  assign track_mem_v_o = (N11)? N78 : 
                         (N12)? 1'b0 : 
                         (N13)? 1'b0 : 
                         (N14)? 1'b0 : 
                         (N15)? 1'b0 : 
                         (N16)? N223 : 
                         (N17)? dma_done_i : 
                         (N18)? 1'b0 : 
                         (N19)? 1'b1 : 
                         (N20)? 1'b0 : 
                         (N21)? 1'b0 : 
                         (N22)? 1'b0 : 1'b0;
  assign miss_state_n = (N11)? { 1'b0, N88, N87, N86 } : 
                        (N12)? { 1'b0, N114, dma_done_i, N113 } : 
                        (N13)? { N152, 1'b0, N151, 1'b1 } : 
                        (N14)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                        (N15)? { 1'b0, dma_done_i, N188, 1'b1 } : 
                        (N16)? { N229, N228, N227, N226 } : 
                        (N17)? { dma_done_i, N188, N188, dma_done_i } : 
                        (N18)? { N261, 1'b0, N260, N260 } : 
                        (N19)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                        (N20)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                        (N21)? { N262, 1'b0, N262, 1'b0 } : 
                        (N22)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign chosen_way_n = (N11)? chosen_way_o : 
                        (N12)? { N93, N92, N91 } : 
                        (N13)? chosen_way_o : 
                        (N14)? chosen_way_o : 
                        (N15)? chosen_way_o : 
                        (N16)? chosen_way_o : 
                        (N17)? chosen_way_o : 
                        (N18)? { N242, N241, N240 } : 
                        (N19)? chosen_way_o : 
                        (N20)? chosen_way_o : 
                        (N21)? chosen_way_o : 
                        (N22)? chosen_way_o : 1'b0;
  assign dma_addr_o[5:4] = (N17)? addr_v_i[5:4] : 
                           (N264)? { 1'b0, 1'b0 } : 1'b0;
  assign dma_addr_o[32:6] = (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N12)? { addr_v_i[32:13], stat_mem_addr_o } : 
                            (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N15)? { N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, stat_mem_addr_o } : 
                            (N16)? { N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, stat_mem_addr_o } : 
                            (N17)? { addr_v_i[32:13], stat_mem_addr_o } : 
                            (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stat_mem_w_o = (N11)? 1'b0 : 
                        (N12)? 1'b0 : 
                        (N13)? 1'b1 : 
                        (N14)? 1'b0 : 
                        (N15)? 1'b0 : 
                        (N16)? 1'b1 : 
                        (N17)? 1'b1 : 
                        (N18)? 1'b0 : 
                        (N19)? 1'b1 : 
                        (N20)? 1'b0 : 
                        (N21)? 1'b0 : 
                        (N22)? 1'b0 : 1'b0;
  assign stat_mem_data_o = (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N16)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, chosen_way_lru_data } : 
                           (N17)? { N230, N230, N230, N230, N230, N230, N230, N230, chosen_way_lru_data } : 
                           (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N19)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, chosen_way_lru_data } : 
                           (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stat_mem_w_mask_o = (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N13)? { flush_way_decode, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N16)? { chosen_way_decode, chosen_way_lru_mask } : 
                             (N17)? { N238, N237, N236, N235, N234, N233, N232, N231, chosen_way_lru_mask } : 
                             (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N19)? { chosen_way_decode, chosen_way_lru_mask } : 
                             (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_mem_v_o = (N11)? 1'b0 : 
                       (N12)? 1'b0 : 
                       (N13)? 1'b1 : 
                       (N14)? 1'b1 : 
                       (N15)? 1'b0 : 
                       (N16)? N222 : 
                       (N17)? dma_done_i : 
                       (N18)? 1'b0 : 
                       (N19)? 1'b1 : 
                       (N20)? 1'b0 : 
                       (N21)? 1'b0 : 
                       (N22)? 1'b0 : 1'b0;
  assign tag_mem_w_o = (N11)? 1'b0 : 
                       (N12)? 1'b0 : 
                       (N13)? 1'b1 : 
                       (N14)? 1'b1 : 
                       (N15)? 1'b0 : 
                       (N16)? 1'b1 : 
                       (N17)? 1'b1 : 
                       (N18)? 1'b0 : 
                       (N19)? 1'b1 : 
                       (N20)? 1'b0 : 
                       (N21)? 1'b0 : 
                       (N22)? 1'b0 : 1'b0;
  assign tag_mem_w_mask_o = (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N13)? { N132, N133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N130, N131, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N128, N129, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N126, N127, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N124, N125, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N122, N123, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N120, N121, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N118, N119, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N14)? { 1'b0, tag_hit_v_i[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tag_hit_v_i[6:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tag_hit_v_i[5:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tag_hit_v_i[4:4], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tag_hit_v_i[3:3], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tag_hit_v_i[2:2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tag_hit_v_i[1:1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tag_hit_v_i[0:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N16)? { chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                            (N17)? { chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                            (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N19)? { chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                            (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_mem_data_o = (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N14)? { 1'b0, decode_v_i[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, decode_v_i[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, decode_v_i[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, decode_v_i[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, decode_v_i[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, decode_v_i[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, decode_v_i[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, decode_v_i[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N16)? { 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13] } : 
                          (N17)? { 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13] } : 
                          (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N19)? { 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13], 1'b1, decode_v_i[7:7], addr_v_i[32:13] } : 
                          (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign track_mem_w_o = (N11)? 1'b0 : 
                         (N12)? 1'b0 : 
                         (N13)? 1'b0 : 
                         (N14)? 1'b0 : 
                         (N15)? 1'b0 : 
                         (N16)? 1'b1 : 
                         (N17)? 1'b1 : 
                         (N18)? 1'b0 : 
                         (N19)? 1'b1 : 
                         (N20)? 1'b0 : 
                         (N21)? 1'b0 : 
                         (N22)? 1'b0 : 1'b0;
  assign track_mem_w_mask_o = (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N16)? { chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                              (N17)? { chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                              (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N19)? { chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:7], chosen_way_decode[7:6], chosen_way_decode[6:6], chosen_way_decode[6:6], chosen_way_decode[6:5], chosen_way_decode[5:5], chosen_way_decode[5:5], chosen_way_decode[5:4], chosen_way_decode[4:4], chosen_way_decode[4:4], chosen_way_decode[4:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                              (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign select_snoop_data_n = (N17)? 1'b1 : 
                               (N21)? 1'b0 : 1'b0;
  assign recover_o = (N11)? 1'b0 : 
                     (N12)? 1'b0 : 
                     (N13)? 1'b0 : 
                     (N14)? 1'b0 : 
                     (N15)? 1'b0 : 
                     (N16)? 1'b0 : 
                     (N17)? 1'b0 : 
                     (N18)? 1'b0 : 
                     (N19)? 1'b0 : 
                     (N20)? 1'b1 : 
                     (N21)? 1'b0 : 
                     (N22)? 1'b0 : 1'b0;
  assign done_o = (N11)? 1'b0 : 
                  (N12)? 1'b0 : 
                  (N13)? 1'b0 : 
                  (N14)? 1'b0 : 
                  (N15)? 1'b0 : 
                  (N16)? 1'b0 : 
                  (N17)? 1'b0 : 
                  (N18)? 1'b0 : 
                  (N19)? 1'b0 : 
                  (N20)? 1'b0 : 
                  (N21)? 1'b1 : 
                  (N22)? 1'b0 : 1'b0;
  assign _0_net__7_ = N297 & N298;
  assign N297 = ~valid_v_i[7];
  assign N298 = ~lock_v_i[7];
  assign _0_net__6_ = N299 & N300;
  assign N299 = ~valid_v_i[6];
  assign N300 = ~lock_v_i[6];
  assign _0_net__5_ = N301 & N302;
  assign N301 = ~valid_v_i[5];
  assign N302 = ~lock_v_i[5];
  assign _0_net__4_ = N303 & N304;
  assign N303 = ~valid_v_i[4];
  assign N304 = ~lock_v_i[4];
  assign _0_net__3_ = N305 & N306;
  assign N305 = ~valid_v_i[3];
  assign N306 = ~lock_v_i[3];
  assign _0_net__2_ = N307 & N308;
  assign N307 = ~valid_v_i[2];
  assign N308 = ~lock_v_i[2];
  assign _0_net__1_ = N309 & N310;
  assign N309 = ~valid_v_i[1];
  assign N310 = ~lock_v_i[1];
  assign _0_net__0_ = N311 & N312;
  assign N311 = ~valid_v_i[0];
  assign N312 = ~lock_v_i[0];
  assign goto_flush_op = N314 | decode_v_i[9];
  assign N314 = N313 | decode_v_i[10];
  assign N313 = decode_v_i[13] | decode_v_i[8];
  assign goto_lock_op = decode_v_i[6] | N315;
  assign N315 = decode_v_i[7] & tag_hit_found_i;
  assign N23 = ~decode_v_i[17];
  assign N24 = N329 & mask_v_i[0];
  assign N329 = N328 & mask_v_i[1];
  assign N328 = N327 & mask_v_i[2];
  assign N327 = N326 & mask_v_i[3];
  assign N326 = N325 & mask_v_i[4];
  assign N325 = N324 & mask_v_i[5];
  assign N324 = N323 & mask_v_i[6];
  assign N323 = N322 & mask_v_i[7];
  assign N322 = N321 & mask_v_i[8];
  assign N321 = N320 & mask_v_i[9];
  assign N320 = N319 & mask_v_i[10];
  assign N319 = N318 & mask_v_i[11];
  assign N318 = N317 & mask_v_i[12];
  assign N317 = N316 & mask_v_i[13];
  assign N316 = mask_v_i[15] & mask_v_i[14];
  assign st_tag_miss_op = N330 & N331;
  assign N330 = decode_v_i[15] & full_word_op;
  assign N331 = ~tag_hit_found_i;
  assign N25 = ~goto_flush_op;
  assign N26 = ~decode_v_i[13];
  assign N27 = ~miss_state_r[3];
  assign N28 = ~miss_state_r[2];
  assign N29 = ~miss_state_r[1];
  assign N30 = ~miss_state_r[0];
  assign N37 = ~N36;
  assign N41 = ~N40;
  assign N45 = ~N44;
  assign N49 = ~N48;
  assign N53 = ~N52;
  assign N57 = ~N56;
  assign N61 = ~N60;
  assign N65 = ~N64;
  assign N69 = ~N68;
  assign N73 = ~N72;
  assign N77 = N75 | N76;
  assign dma_cmd_o[0] = N37;
  assign dma_cmd_o[1] = N49;
  assign dma_cmd_o[3] = N53;
  assign track_mem_data_o_7__3_ = N57;
  assign N78 = N332 & tbuf_empty_i;
  assign N332 = miss_v_i & sbuf_empty_i;
  assign N79 = ~N78;
  assign N80 = goto_lock_op | goto_flush_op;
  assign N81 = st_tag_miss_op | N80;
  assign N82 = ~N81;
  assign N89 = invalid_exist | track_miss_i;
  assign N90 = ~N89;
  assign N94 = ~N91;
  assign N95 = ~N92;
  assign N96 = N94 & N95;
  assign N97 = N94 & N92;
  assign N98 = N91 & N95;
  assign N99 = N91 & N92;
  assign N100 = ~N93;
  assign N101 = N96 & N100;
  assign N102 = N96 & N93;
  assign N103 = N98 & N100;
  assign N104 = N98 & N93;
  assign N105 = N97 & N100;
  assign N106 = N97 & N93;
  assign N107 = N99 & N100;
  assign N108 = N99 & N93;
  assign N111 = N334 & N110;
  assign N334 = N333 & N109;
  assign N333 = ~track_miss_i;
  assign N118 = N335 & flush_way_decode[0];
  assign N335 = decode_v_i[8] | decode_v_i[9];
  assign N119 = N336 & flush_way_decode[0];
  assign N336 = decode_v_i[8] | decode_v_i[9];
  assign N120 = N337 & flush_way_decode[1];
  assign N337 = decode_v_i[8] | decode_v_i[9];
  assign N121 = N338 & flush_way_decode[1];
  assign N338 = decode_v_i[8] | decode_v_i[9];
  assign N122 = N339 & flush_way_decode[2];
  assign N339 = decode_v_i[8] | decode_v_i[9];
  assign N123 = N340 & flush_way_decode[2];
  assign N340 = decode_v_i[8] | decode_v_i[9];
  assign N124 = N341 & flush_way_decode[3];
  assign N341 = decode_v_i[8] | decode_v_i[9];
  assign N125 = N342 & flush_way_decode[3];
  assign N342 = decode_v_i[8] | decode_v_i[9];
  assign N126 = N343 & flush_way_decode[4];
  assign N343 = decode_v_i[8] | decode_v_i[9];
  assign N127 = N344 & flush_way_decode[4];
  assign N344 = decode_v_i[8] | decode_v_i[9];
  assign N128 = N345 & flush_way_decode[5];
  assign N345 = decode_v_i[8] | decode_v_i[9];
  assign N129 = N346 & flush_way_decode[5];
  assign N346 = decode_v_i[8] | decode_v_i[9];
  assign N130 = N347 & flush_way_decode[6];
  assign N347 = decode_v_i[8] | decode_v_i[9];
  assign N131 = N348 & flush_way_decode[6];
  assign N348 = decode_v_i[8] | decode_v_i[9];
  assign N132 = N349 & flush_way_decode[7];
  assign N349 = decode_v_i[8] | decode_v_i[9];
  assign N133 = N350 & flush_way_decode[7];
  assign N350 = decode_v_i[8] | decode_v_i[9];
  assign N134 = ~N115;
  assign N135 = ~N116;
  assign N136 = N134 & N135;
  assign N137 = N134 & N116;
  assign N138 = N115 & N135;
  assign N139 = N115 & N116;
  assign N140 = ~N117;
  assign N141 = N136 & N140;
  assign N142 = N136 & N117;
  assign N143 = N138 & N140;
  assign N144 = N138 & N117;
  assign N145 = N137 & N140;
  assign N146 = N137 & N117;
  assign N147 = N139 & N140;
  assign N148 = N139 & N117;
  assign N151 = N352 & N150;
  assign N352 = N351 & N149;
  assign N351 = ~decode_v_i[8];
  assign N153 = ~dma_way_o[0];
  assign N154 = ~dma_way_o[1];
  assign N155 = N153 & N154;
  assign N156 = N153 & dma_way_o[1];
  assign N157 = dma_way_o[0] & N154;
  assign N158 = dma_way_o[0] & dma_way_o[1];
  assign N159 = ~dma_way_o[2];
  assign N160 = N155 & N159;
  assign N161 = N155 & dma_way_o[2];
  assign N162 = N157 & N159;
  assign N163 = N157 & dma_way_o[2];
  assign N164 = N156 & N159;
  assign N165 = N156 & dma_way_o[2];
  assign N166 = N158 & N159;
  assign N167 = N158 & dma_way_o[2];
  assign N188 = ~dma_done_i;
  assign N189 = N153 & N154;
  assign N190 = N153 & dma_way_o[1];
  assign N191 = dma_way_o[0] & N154;
  assign N192 = dma_way_o[0] & dma_way_o[1];
  assign N193 = N189 & N159;
  assign N194 = N189 & dma_way_o[2];
  assign N195 = N191 & N159;
  assign N196 = N191 & dma_way_o[2];
  assign N197 = N190 & N159;
  assign N198 = N190 & dma_way_o[2];
  assign N199 = N192 & N159;
  assign N200 = N192 & dma_way_o[2];
  assign N221 = dma_done_i & st_tag_miss_op;
  assign N222 = dma_done_i & st_tag_miss_op;
  assign N223 = dma_done_i & st_tag_miss_op;
  assign N224 = N354 | st_tag_miss_op;
  assign N354 = N353 | decode_v_i[10];
  assign N353 = decode_v_i[13] | decode_v_i[9];
  assign N230 = decode_v_i[15] | decode_v_i[4];
  assign N239 = ~invalid_exist;
  assign N243 = ~N240;
  assign N244 = ~N241;
  assign N245 = N243 & N244;
  assign N246 = N243 & N241;
  assign N247 = N240 & N244;
  assign N248 = N240 & N241;
  assign N249 = ~N242;
  assign N250 = N245 & N249;
  assign N251 = N245 & N242;
  assign N252 = N247 & N249;
  assign N253 = N247 & N242;
  assign N254 = N246 & N249;
  assign N255 = N246 & N242;
  assign N256 = N248 & N249;
  assign N257 = N248 & N242;
  assign N260 = N258 & N259;
  assign N262 = ~ack_i;
  assign N263 = ~track_mem_data_o_7__3_;
  assign N264 = N263;
  assign N265 = ~goto_flush_op;
  assign N266 = goto_lock_op & N265;
  assign N267 = ~goto_lock_op;
  assign N268 = N265 & N267;
  assign N269 = st_tag_miss_op & N268;
  assign N270 = ~track_miss_i;
  assign N271 = invalid_exist & N270;
  assign N272 = track_mem_v_o & N355;
  assign N355 = ~track_mem_w_o;
  assign N273 = N33 | dma_cmd_o[0];
  assign N274 = N273 | N45;
  assign N275 = N274 | dma_cmd_o[1];
  assign N276 = N275 | dma_cmd_o[3];
  assign N277 = N276 | track_mem_data_o_7__3_;
  assign N278 = N277 | N61;
  assign N279 = N278 | N65;
  assign N280 = N279 | N69;
  assign N281 = N280 | N73;
  assign N282 = N281 | N77;
  assign N283 = ~N282;
  assign N284 = N273 | N41;
  assign N285 = N284 | N45;
  assign N286 = N285 | dma_cmd_o[1];
  assign N287 = N286 | dma_cmd_o[3];
  assign N288 = N188 & track_mem_data_o_7__3_;
  assign N289 = N287 | N288;
  assign N290 = N289 | N61;
  assign N291 = N290 | N65;
  assign N292 = N291 | N69;
  assign N293 = N262 & N73;
  assign N294 = N292 | N293;
  assign N295 = N294 | N77;
  assign N296 = ~N295;

  always @(posedge clk_i) begin
    if(reset_i) begin
      track_data_we_o_sv2v_reg <= 1'b0;
      miss_state_r_3_sv2v_reg <= 1'b0;
      miss_state_r_2_sv2v_reg <= 1'b0;
      miss_state_r_1_sv2v_reg <= 1'b0;
      miss_state_r_0_sv2v_reg <= 1'b0;
      chosen_way_o_2_sv2v_reg <= 1'b0;
      chosen_way_o_1_sv2v_reg <= 1'b0;
      chosen_way_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      track_data_we_o_sv2v_reg <= N272;
      miss_state_r_3_sv2v_reg <= miss_state_n[3];
      miss_state_r_2_sv2v_reg <= miss_state_n[2];
      miss_state_r_1_sv2v_reg <= miss_state_n[1];
      miss_state_r_0_sv2v_reg <= miss_state_n[0];
      chosen_way_o_2_sv2v_reg <= chosen_way_n[2];
      chosen_way_o_1_sv2v_reg <= chosen_way_n[1];
      chosen_way_o_0_sv2v_reg <= chosen_way_n[0];
    end 
    if(reset_i) begin
      flush_way_r_2_sv2v_reg <= 1'b0;
      flush_way_r_1_sv2v_reg <= 1'b0;
      flush_way_r_0_sv2v_reg <= 1'b0;
    end else if(N283) begin
      flush_way_r_2_sv2v_reg <= N117;
      flush_way_r_1_sv2v_reg <= N116;
      flush_way_r_0_sv2v_reg <= N115;
    end 
    if(reset_i) begin
      select_snoop_data_r_o_sv2v_reg <= 1'b0;
    end else if(N296) begin
      select_snoop_data_r_o_sv2v_reg <= select_snoop_data_n;
    end 
  end


endmodule



module bsg_counter_clear_up_00000004_0
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [2:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire [2:0] count_o;
  wire N0,N1,N4,N5,N6,N8,N9,N10,N11,N12,N13,N14,N15,N2,N3,N7,N30,N16;
  reg count_o_2_sv2v_reg,count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[2] = count_o_2_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign N16 = reset_i | clear_i;
  assign { N8, N6, N5 } = count_o + 1'b1;
  assign N9 = (N0)? 1'b1 : 
              (N7)? 1'b1 : 
              (N3)? 1'b0 : 1'b0;
  assign N0 = clear_i;
  assign N11 = (N1)? 1'b1 : 
               (N30)? 1'b0 : 1'b0;
  assign N1 = up_i;
  assign N10 = (N0)? up_i : 
               (N7)? N5 : 1'b0;
  assign N4 = N15;
  assign N12 = ~reset_i;
  assign N13 = ~clear_i;
  assign N14 = N12 & N13;
  assign N15 = up_i & N14;
  assign N2 = up_i | clear_i;
  assign N3 = ~N2;
  assign N7 = up_i & N13;
  assign N30 = ~up_i;

  always @(posedge clk_i) begin
    if(N16) begin
      count_o_2_sv2v_reg <= 1'b0;
      count_o_1_sv2v_reg <= 1'b0;
    end else if(N11) begin
      count_o_2_sv2v_reg <= N8;
      count_o_1_sv2v_reg <= N6;
    end 
    if(reset_i) begin
      count_o_0_sv2v_reg <= 1'b0;
    end else if(N9) begin
      count_o_0_sv2v_reg <= N10;
    end 
  end


endmodule



module bsg_fifo_1r1w_small_unhardened_00000080_00000004_0
(
  clk_i,
  reset_i,
  v_i,
  ready_param_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [127:0] data_i;
  output [127:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_param_o;
  output v_o;
  wire [127:0] data_o;
  wire ready_param_o,v_o,enque,full,empty,sv2v_dc_1,sv2v_dc_2;
  wire [1:0] wptr_r,rptr_r;

  bsg_fifo_tracker_00000004
  ft
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .enq_i(enque),
    .deq_i(yumi_i),
    .wptr_r_o(wptr_r),
    .rptr_r_o(rptr_r),
    .rptr_n_o({ sv2v_dc_1, sv2v_dc_2 }),
    .full_o(full),
    .empty_o(empty)
  );


  bsg_mem_1r1w
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enque),
    .w_addr_i(wptr_r),
    .w_data_i(data_i),
    .r_v_i(v_o),
    .r_addr_i(rptr_r),
    .r_data_o(data_o)
  );

  assign enque = v_i & ready_param_o;
  assign ready_param_o = ~full;
  assign v_o = ~empty;

endmodule



module bsg_fifo_1r1w_small_00000080_00000004
(
  clk_i,
  reset_i,
  v_i,
  ready_param_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [127:0] data_i;
  output [127:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_param_o;
  output v_o;
  wire [127:0] data_o;
  wire ready_param_o,v_o;

  bsg_fifo_1r1w_small_unhardened_00000080_00000004_0
  \unhardened.un.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_param_o(ready_param_o),
    .data_i(data_i),
    .v_o(v_o),
    .data_o(data_o),
    .yumi_i(yumi_i)
  );


endmodule



module bsg_two_fifo_00000080
(
  clk_i,
  reset_i,
  ready_param_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [127:0] data_i;
  output [127:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_param_o;
  output v_o;
  wire [127:0] data_o;
  wire ready_param_o,v_o,enq_i,tail_r,_0_net_,head_r,empty_r,full_r,N0,N1,N2,N3,N4,N5,
  N6,N7,N8,N9,N10,N11,N12,N13,N14;
  reg full_r_sv2v_reg,tail_r_sv2v_reg,head_r_sv2v_reg,empty_r_sv2v_reg;
  assign full_r = full_r_sv2v_reg;
  assign tail_r = tail_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign empty_r = empty_r_sv2v_reg;

  bsg_mem_1r1w
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign _0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_param_o = ~full_r;
  assign enq_i = v_i & N5;
  assign N5 = ~full_r;
  assign N1 = enq_i;
  assign N0 = ~tail_r;
  assign N2 = ~head_r;
  assign N3 = N7 | N9;
  assign N7 = empty_r & N6;
  assign N6 = ~enq_i;
  assign N9 = N8 & N6;
  assign N8 = N5 & yumi_i;
  assign N4 = N13 | N14;
  assign N13 = N11 & N12;
  assign N11 = N10 & enq_i;
  assign N10 = ~empty_r;
  assign N12 = ~yumi_i;
  assign N14 = full_r & N12;

  always @(posedge clk_i) begin
    if(reset_i) begin
      full_r_sv2v_reg <= 1'b0;
      empty_r_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      full_r_sv2v_reg <= N4;
      empty_r_sv2v_reg <= N3;
    end 
    if(reset_i) begin
      tail_r_sv2v_reg <= 1'b0;
    end else if(N1) begin
      tail_r_sv2v_reg <= N0;
    end 
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_expand_bitmask_00000008_00000010
(
  i,
  o
);

  input [7:0] i;
  output [127:0] o;
  wire [127:0] o;
  wire o_127_,o_111_,o_95_,o_79_,o_63_,o_47_,o_31_,o_15_;
  assign o_127_ = i[7];
  assign o[112] = o_127_;
  assign o[113] = o_127_;
  assign o[114] = o_127_;
  assign o[115] = o_127_;
  assign o[116] = o_127_;
  assign o[117] = o_127_;
  assign o[118] = o_127_;
  assign o[119] = o_127_;
  assign o[120] = o_127_;
  assign o[121] = o_127_;
  assign o[122] = o_127_;
  assign o[123] = o_127_;
  assign o[124] = o_127_;
  assign o[125] = o_127_;
  assign o[126] = o_127_;
  assign o[127] = o_127_;
  assign o_111_ = i[6];
  assign o[96] = o_111_;
  assign o[97] = o_111_;
  assign o[98] = o_111_;
  assign o[99] = o_111_;
  assign o[100] = o_111_;
  assign o[101] = o_111_;
  assign o[102] = o_111_;
  assign o[103] = o_111_;
  assign o[104] = o_111_;
  assign o[105] = o_111_;
  assign o[106] = o_111_;
  assign o[107] = o_111_;
  assign o[108] = o_111_;
  assign o[109] = o_111_;
  assign o[110] = o_111_;
  assign o[111] = o_111_;
  assign o_95_ = i[5];
  assign o[80] = o_95_;
  assign o[81] = o_95_;
  assign o[82] = o_95_;
  assign o[83] = o_95_;
  assign o[84] = o_95_;
  assign o[85] = o_95_;
  assign o[86] = o_95_;
  assign o[87] = o_95_;
  assign o[88] = o_95_;
  assign o[89] = o_95_;
  assign o[90] = o_95_;
  assign o[91] = o_95_;
  assign o[92] = o_95_;
  assign o[93] = o_95_;
  assign o[94] = o_95_;
  assign o[95] = o_95_;
  assign o_79_ = i[4];
  assign o[64] = o_79_;
  assign o[65] = o_79_;
  assign o[66] = o_79_;
  assign o[67] = o_79_;
  assign o[68] = o_79_;
  assign o[69] = o_79_;
  assign o[70] = o_79_;
  assign o[71] = o_79_;
  assign o[72] = o_79_;
  assign o[73] = o_79_;
  assign o[74] = o_79_;
  assign o[75] = o_79_;
  assign o[76] = o_79_;
  assign o[77] = o_79_;
  assign o[78] = o_79_;
  assign o[79] = o_79_;
  assign o_63_ = i[3];
  assign o[48] = o_63_;
  assign o[49] = o_63_;
  assign o[50] = o_63_;
  assign o[51] = o_63_;
  assign o[52] = o_63_;
  assign o[53] = o_63_;
  assign o[54] = o_63_;
  assign o[55] = o_63_;
  assign o[56] = o_63_;
  assign o[57] = o_63_;
  assign o[58] = o_63_;
  assign o[59] = o_63_;
  assign o[60] = o_63_;
  assign o[61] = o_63_;
  assign o[62] = o_63_;
  assign o[63] = o_63_;
  assign o_47_ = i[2];
  assign o[32] = o_47_;
  assign o[33] = o_47_;
  assign o[34] = o_47_;
  assign o[35] = o_47_;
  assign o[36] = o_47_;
  assign o[37] = o_47_;
  assign o[38] = o_47_;
  assign o[39] = o_47_;
  assign o[40] = o_47_;
  assign o[41] = o_47_;
  assign o[42] = o_47_;
  assign o[43] = o_47_;
  assign o[44] = o_47_;
  assign o[45] = o_47_;
  assign o[46] = o_47_;
  assign o[47] = o_47_;
  assign o_31_ = i[1];
  assign o[16] = o_31_;
  assign o[17] = o_31_;
  assign o[18] = o_31_;
  assign o[19] = o_31_;
  assign o[20] = o_31_;
  assign o[21] = o_31_;
  assign o[22] = o_31_;
  assign o[23] = o_31_;
  assign o[24] = o_31_;
  assign o[25] = o_31_;
  assign o[26] = o_31_;
  assign o[27] = o_31_;
  assign o[28] = o_31_;
  assign o[29] = o_31_;
  assign o[30] = o_31_;
  assign o[31] = o_31_;
  assign o_15_ = i[0];
  assign o[0] = o_15_;
  assign o[1] = o_15_;
  assign o[2] = o_15_;
  assign o[3] = o_15_;
  assign o[4] = o_15_;
  assign o[5] = o_15_;
  assign o[6] = o_15_;
  assign o[7] = o_15_;
  assign o[8] = o_15_;
  assign o[9] = o_15_;
  assign o[10] = o_15_;
  assign o[11] = o_15_;
  assign o[12] = o_15_;
  assign o[13] = o_15_;
  assign o[14] = o_15_;
  assign o[15] = o_15_;

endmodule



module bsg_mux_00000004_00000008
(
  data_i,
  sel_i,
  data_o
);

  input [31:0] data_i;
  input [2:0] sel_i;
  output [3:0] data_o;
  wire [3:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;
  assign data_o[3] = (N7)? data_i[3] : 
                     (N9)? data_i[7] : 
                     (N11)? data_i[11] : 
                     (N13)? data_i[15] : 
                     (N8)? data_i[19] : 
                     (N10)? data_i[23] : 
                     (N12)? data_i[27] : 
                     (N14)? data_i[31] : 1'b0;
  assign data_o[2] = (N7)? data_i[2] : 
                     (N9)? data_i[6] : 
                     (N11)? data_i[10] : 
                     (N13)? data_i[14] : 
                     (N8)? data_i[18] : 
                     (N10)? data_i[22] : 
                     (N12)? data_i[26] : 
                     (N14)? data_i[30] : 1'b0;
  assign data_o[1] = (N7)? data_i[1] : 
                     (N9)? data_i[5] : 
                     (N11)? data_i[9] : 
                     (N13)? data_i[13] : 
                     (N8)? data_i[17] : 
                     (N10)? data_i[21] : 
                     (N12)? data_i[25] : 
                     (N14)? data_i[29] : 1'b0;
  assign data_o[0] = (N7)? data_i[0] : 
                     (N9)? data_i[4] : 
                     (N11)? data_i[8] : 
                     (N13)? data_i[12] : 
                     (N8)? data_i[16] : 
                     (N10)? data_i[20] : 
                     (N12)? data_i[24] : 
                     (N14)? data_i[28] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];
  assign N6 = ~sel_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & sel_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & sel_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & sel_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & sel_i[2];

endmodule



module bsg_expand_bitmask_00000001_00000010
(
  i,
  o
);

  input [0:0] i;
  output [15:0] o;
  wire [15:0] o;
  wire o_15_;
  assign o_15_ = i[0];
  assign o[0] = o_15_;
  assign o[1] = o_15_;
  assign o[2] = o_15_;
  assign o[3] = o_15_;
  assign o[4] = o_15_;
  assign o[5] = o_15_;
  assign o[6] = o_15_;
  assign o[7] = o_15_;
  assign o[8] = o_15_;
  assign o[9] = o_15_;
  assign o[10] = o_15_;
  assign o[11] = o_15_;
  assign o[12] = o_15_;
  assign o[13] = o_15_;
  assign o[14] = o_15_;
  assign o[15] = o_15_;

endmodule



module bsg_mux_00000080_00000001
(
  data_i,
  sel_i,
  data_o
);

  input [127:0] data_i;
  input [0:0] sel_i;
  output [127:0] data_o;
  wire [127:0] data_o;
  assign data_o[127] = data_i[127];
  assign data_o[126] = data_i[126];
  assign data_o[125] = data_i[125];
  assign data_o[124] = data_i[124];
  assign data_o[123] = data_i[123];
  assign data_o[122] = data_i[122];
  assign data_o[121] = data_i[121];
  assign data_o[120] = data_i[120];
  assign data_o[119] = data_i[119];
  assign data_o[118] = data_i[118];
  assign data_o[117] = data_i[117];
  assign data_o[116] = data_i[116];
  assign data_o[115] = data_i[115];
  assign data_o[114] = data_i[114];
  assign data_o[113] = data_i[113];
  assign data_o[112] = data_i[112];
  assign data_o[111] = data_i[111];
  assign data_o[110] = data_i[110];
  assign data_o[109] = data_i[109];
  assign data_o[108] = data_i[108];
  assign data_o[107] = data_i[107];
  assign data_o[106] = data_i[106];
  assign data_o[105] = data_i[105];
  assign data_o[104] = data_i[104];
  assign data_o[103] = data_i[103];
  assign data_o[102] = data_i[102];
  assign data_o[101] = data_i[101];
  assign data_o[100] = data_i[100];
  assign data_o[99] = data_i[99];
  assign data_o[98] = data_i[98];
  assign data_o[97] = data_i[97];
  assign data_o[96] = data_i[96];
  assign data_o[95] = data_i[95];
  assign data_o[94] = data_i[94];
  assign data_o[93] = data_i[93];
  assign data_o[92] = data_i[92];
  assign data_o[91] = data_i[91];
  assign data_o[90] = data_i[90];
  assign data_o[89] = data_i[89];
  assign data_o[88] = data_i[88];
  assign data_o[87] = data_i[87];
  assign data_o[86] = data_i[86];
  assign data_o[85] = data_i[85];
  assign data_o[84] = data_i[84];
  assign data_o[83] = data_i[83];
  assign data_o[82] = data_i[82];
  assign data_o[81] = data_i[81];
  assign data_o[80] = data_i[80];
  assign data_o[79] = data_i[79];
  assign data_o[78] = data_i[78];
  assign data_o[77] = data_i[77];
  assign data_o[76] = data_i[76];
  assign data_o[75] = data_i[75];
  assign data_o[74] = data_i[74];
  assign data_o[73] = data_i[73];
  assign data_o[72] = data_i[72];
  assign data_o[71] = data_i[71];
  assign data_o[70] = data_i[70];
  assign data_o[69] = data_i[69];
  assign data_o[68] = data_i[68];
  assign data_o[67] = data_i[67];
  assign data_o[66] = data_i[66];
  assign data_o[65] = data_i[65];
  assign data_o[64] = data_i[64];
  assign data_o[63] = data_i[63];
  assign data_o[62] = data_i[62];
  assign data_o[61] = data_i[61];
  assign data_o[60] = data_i[60];
  assign data_o[59] = data_i[59];
  assign data_o[58] = data_i[58];
  assign data_o[57] = data_i[57];
  assign data_o[56] = data_i[56];
  assign data_o[55] = data_i[55];
  assign data_o[54] = data_i[54];
  assign data_o[53] = data_i[53];
  assign data_o[52] = data_i[52];
  assign data_o[51] = data_i[51];
  assign data_o[50] = data_i[50];
  assign data_o[49] = data_i[49];
  assign data_o[48] = data_i[48];
  assign data_o[47] = data_i[47];
  assign data_o[46] = data_i[46];
  assign data_o[45] = data_i[45];
  assign data_o[44] = data_i[44];
  assign data_o[43] = data_i[43];
  assign data_o[42] = data_i[42];
  assign data_o[41] = data_i[41];
  assign data_o[40] = data_i[40];
  assign data_o[39] = data_i[39];
  assign data_o[38] = data_i[38];
  assign data_o[37] = data_i[37];
  assign data_o[36] = data_i[36];
  assign data_o[35] = data_i[35];
  assign data_o[34] = data_i[34];
  assign data_o[33] = data_i[33];
  assign data_o[32] = data_i[32];
  assign data_o[31] = data_i[31];
  assign data_o[30] = data_i[30];
  assign data_o[29] = data_i[29];
  assign data_o[28] = data_i[28];
  assign data_o[27] = data_i[27];
  assign data_o[26] = data_i[26];
  assign data_o[25] = data_i[25];
  assign data_o[24] = data_i[24];
  assign data_o[23] = data_i[23];
  assign data_o[22] = data_i[22];
  assign data_o[21] = data_i[21];
  assign data_o[20] = data_i[20];
  assign data_o[19] = data_i[19];
  assign data_o[18] = data_i[18];
  assign data_o[17] = data_i[17];
  assign data_o[16] = data_i[16];
  assign data_o[15] = data_i[15];
  assign data_o[14] = data_i[14];
  assign data_o[13] = data_i[13];
  assign data_o[12] = data_i[12];
  assign data_o[11] = data_i[11];
  assign data_o[10] = data_i[10];
  assign data_o[9] = data_i[9];
  assign data_o[8] = data_i[8];
  assign data_o[7] = data_i[7];
  assign data_o[6] = data_i[6];
  assign data_o[5] = data_i[5];
  assign data_o[4] = data_i[4];
  assign data_o[3] = data_i[3];
  assign data_o[2] = data_i[2];
  assign data_o[1] = data_i[1];
  assign data_o[0] = data_i[0];

endmodule



module bsg_cache_dma_00000021_00000080_00000004_00000080_00000008_1_00000080_0
(
  clk_i,
  reset_i,
  dma_cmd_i,
  dma_way_i,
  dma_addr_i,
  done_o,
  track_data_we_i,
  snoop_word_o,
  dma_pkt_o,
  dma_pkt_v_o,
  dma_pkt_yumi_i,
  dma_data_i,
  dma_data_v_i,
  dma_data_ready_and_o,
  dma_data_o,
  dma_data_v_o,
  dma_data_yumi_i,
  data_mem_v_o,
  data_mem_w_o,
  data_mem_addr_o,
  data_mem_w_mask_o,
  data_mem_data_o,
  data_mem_data_i,
  track_miss_i,
  track_mem_data_i,
  dma_evict_o
);

  input [3:0] dma_cmd_i;
  input [2:0] dma_way_i;
  input [32:0] dma_addr_i;
  output [127:0] snoop_word_o;
  output [37:0] dma_pkt_o;
  input [127:0] dma_data_i;
  output [127:0] dma_data_o;
  output [8:0] data_mem_addr_o;
  output [127:0] data_mem_w_mask_o;
  output [1023:0] data_mem_data_o;
  input [1023:0] data_mem_data_i;
  input [31:0] track_mem_data_i;
  input clk_i;
  input reset_i;
  input track_data_we_i;
  input dma_pkt_yumi_i;
  input dma_data_v_i;
  input dma_data_yumi_i;
  input track_miss_i;
  output done_o;
  output dma_pkt_v_o;
  output dma_data_ready_and_o;
  output dma_data_v_o;
  output data_mem_v_o;
  output data_mem_w_o;
  output dma_evict_o;
  wire [127:0] snoop_word_o,dma_data_o,data_mem_w_mask_o,out_fifo_data_li,
  dma_way_mask_expanded,snoop_word_n;
  wire [37:0] dma_pkt_o;
  wire [8:0] data_mem_addr_o;
  wire [1023:0] data_mem_data_o;
  wire done_o,dma_pkt_v_o,dma_data_ready_and_o,dma_data_v_o,data_mem_v_o,data_mem_w_o,
  dma_evict_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,dma_pkt_o_36_,dma_pkt_o_35_,
  dma_pkt_o_34_,dma_pkt_o_33_,dma_pkt_o_32_,dma_pkt_o_31_,dma_pkt_o_30_,
  dma_pkt_o_29_,dma_pkt_o_28_,dma_pkt_o_27_,dma_pkt_o_26_,dma_pkt_o_25_,dma_pkt_o_24_,
  dma_pkt_o_23_,dma_pkt_o_22_,dma_pkt_o_21_,dma_pkt_o_20_,dma_pkt_o_19_,dma_pkt_o_18_,
  dma_pkt_o_17_,data_mem_addr_o_8_,data_mem_addr_o_7_,data_mem_addr_o_6_,
  data_mem_addr_o_5_,data_mem_addr_o_4_,data_mem_addr_o_3_,data_mem_addr_o_2_,
  data_mem_data_o_7__127_,data_mem_data_o_7__126_,data_mem_data_o_7__125_,data_mem_data_o_7__124_,
  data_mem_data_o_7__123_,data_mem_data_o_7__122_,data_mem_data_o_7__121_,
  data_mem_data_o_7__120_,data_mem_data_o_7__119_,data_mem_data_o_7__118_,
  data_mem_data_o_7__117_,data_mem_data_o_7__116_,data_mem_data_o_7__115_,data_mem_data_o_7__114_,
  data_mem_data_o_7__113_,data_mem_data_o_7__112_,data_mem_data_o_7__111_,
  data_mem_data_o_7__110_,data_mem_data_o_7__109_,data_mem_data_o_7__108_,
  data_mem_data_o_7__107_,data_mem_data_o_7__106_,data_mem_data_o_7__105_,data_mem_data_o_7__104_,
  data_mem_data_o_7__103_,data_mem_data_o_7__102_,data_mem_data_o_7__101_,
  data_mem_data_o_7__100_,data_mem_data_o_7__99_,data_mem_data_o_7__98_,
  data_mem_data_o_7__97_,data_mem_data_o_7__96_,data_mem_data_o_7__95_,data_mem_data_o_7__94_,
  data_mem_data_o_7__93_,data_mem_data_o_7__92_,data_mem_data_o_7__91_,
  data_mem_data_o_7__90_,data_mem_data_o_7__89_,data_mem_data_o_7__88_,data_mem_data_o_7__87_,
  data_mem_data_o_7__86_,data_mem_data_o_7__85_,data_mem_data_o_7__84_,
  data_mem_data_o_7__83_,data_mem_data_o_7__82_,data_mem_data_o_7__81_,data_mem_data_o_7__80_,
  data_mem_data_o_7__79_,data_mem_data_o_7__78_,data_mem_data_o_7__77_,
  data_mem_data_o_7__76_,data_mem_data_o_7__75_,data_mem_data_o_7__74_,data_mem_data_o_7__73_,
  data_mem_data_o_7__72_,data_mem_data_o_7__71_,data_mem_data_o_7__70_,
  data_mem_data_o_7__69_,data_mem_data_o_7__68_,data_mem_data_o_7__67_,data_mem_data_o_7__66_,
  data_mem_data_o_7__65_,data_mem_data_o_7__64_,data_mem_data_o_7__63_,
  data_mem_data_o_7__62_,data_mem_data_o_7__61_,data_mem_data_o_7__60_,data_mem_data_o_7__59_,
  data_mem_data_o_7__58_,data_mem_data_o_7__57_,data_mem_data_o_7__56_,
  data_mem_data_o_7__55_,data_mem_data_o_7__54_,data_mem_data_o_7__53_,data_mem_data_o_7__52_,
  data_mem_data_o_7__51_,data_mem_data_o_7__50_,data_mem_data_o_7__49_,
  data_mem_data_o_7__48_,data_mem_data_o_7__47_,data_mem_data_o_7__46_,data_mem_data_o_7__45_,
  data_mem_data_o_7__44_,data_mem_data_o_7__43_,data_mem_data_o_7__42_,
  data_mem_data_o_7__41_,data_mem_data_o_7__40_,data_mem_data_o_7__39_,data_mem_data_o_7__38_,
  data_mem_data_o_7__37_,data_mem_data_o_7__36_,data_mem_data_o_7__35_,
  data_mem_data_o_7__34_,data_mem_data_o_7__33_,data_mem_data_o_7__32_,
  data_mem_data_o_7__31_,data_mem_data_o_7__30_,data_mem_data_o_7__29_,data_mem_data_o_7__28_,
  data_mem_data_o_7__27_,data_mem_data_o_7__26_,data_mem_data_o_7__25_,
  data_mem_data_o_7__24_,data_mem_data_o_7__23_,data_mem_data_o_7__22_,data_mem_data_o_7__21_,
  data_mem_data_o_7__20_,data_mem_data_o_7__19_,data_mem_data_o_7__18_,
  data_mem_data_o_7__17_,data_mem_data_o_7__16_,data_mem_data_o_7__15_,data_mem_data_o_7__14_,
  data_mem_data_o_7__13_,data_mem_data_o_7__12_,data_mem_data_o_7__11_,
  data_mem_data_o_7__10_,data_mem_data_o_7__9_,data_mem_data_o_7__8_,data_mem_data_o_7__7_,
  data_mem_data_o_7__6_,data_mem_data_o_7__5_,data_mem_data_o_7__4_,data_mem_data_o_7__3_,
  data_mem_data_o_7__2_,data_mem_data_o_7__1_,data_mem_data_o_7__0_,counter_clear,
  counter_up,in_fifo_v_lo,in_fifo_yumi_li,out_fifo_v_li,out_fifo_ready_lo,N12,N13,
  N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,
  N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,
  N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,snoop_word_we,N84,N85,N86,N87,N88,N89,N90,
  N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102;
  wire [2:2] counter_r;
  wire [7:0] dma_way_mask;
  wire [31:0] track_mem_data_r;
  wire [3:0] track_data_way_picked;
  wire [0:0] track_bits_offset_picked;
  wire [15:0] track_bits_offset_picked_expanded,data_mem_w_mask_way_picked;
  wire [1:0] dma_state_r,dma_state_n;
  reg track_mem_data_r_31_sv2v_reg,track_mem_data_r_30_sv2v_reg,
  track_mem_data_r_29_sv2v_reg,track_mem_data_r_28_sv2v_reg,track_mem_data_r_27_sv2v_reg,
  track_mem_data_r_26_sv2v_reg,track_mem_data_r_25_sv2v_reg,track_mem_data_r_24_sv2v_reg,
  track_mem_data_r_23_sv2v_reg,track_mem_data_r_22_sv2v_reg,track_mem_data_r_21_sv2v_reg,
  track_mem_data_r_20_sv2v_reg,track_mem_data_r_19_sv2v_reg,
  track_mem_data_r_18_sv2v_reg,track_mem_data_r_17_sv2v_reg,track_mem_data_r_16_sv2v_reg,
  track_mem_data_r_15_sv2v_reg,track_mem_data_r_14_sv2v_reg,track_mem_data_r_13_sv2v_reg,
  track_mem_data_r_12_sv2v_reg,track_mem_data_r_11_sv2v_reg,track_mem_data_r_10_sv2v_reg,
  track_mem_data_r_9_sv2v_reg,track_mem_data_r_8_sv2v_reg,
  track_mem_data_r_7_sv2v_reg,track_mem_data_r_6_sv2v_reg,track_mem_data_r_5_sv2v_reg,
  track_mem_data_r_4_sv2v_reg,track_mem_data_r_3_sv2v_reg,track_mem_data_r_2_sv2v_reg,
  track_mem_data_r_1_sv2v_reg,track_mem_data_r_0_sv2v_reg,dma_state_r_1_sv2v_reg,
  dma_state_r_0_sv2v_reg,snoop_word_o_127_sv2v_reg,snoop_word_o_126_sv2v_reg,
  snoop_word_o_125_sv2v_reg,snoop_word_o_124_sv2v_reg,snoop_word_o_123_sv2v_reg,snoop_word_o_122_sv2v_reg,
  snoop_word_o_121_sv2v_reg,snoop_word_o_120_sv2v_reg,snoop_word_o_119_sv2v_reg,
  snoop_word_o_118_sv2v_reg,snoop_word_o_117_sv2v_reg,snoop_word_o_116_sv2v_reg,
  snoop_word_o_115_sv2v_reg,snoop_word_o_114_sv2v_reg,snoop_word_o_113_sv2v_reg,
  snoop_word_o_112_sv2v_reg,snoop_word_o_111_sv2v_reg,snoop_word_o_110_sv2v_reg,
  snoop_word_o_109_sv2v_reg,snoop_word_o_108_sv2v_reg,snoop_word_o_107_sv2v_reg,
  snoop_word_o_106_sv2v_reg,snoop_word_o_105_sv2v_reg,snoop_word_o_104_sv2v_reg,
  snoop_word_o_103_sv2v_reg,snoop_word_o_102_sv2v_reg,snoop_word_o_101_sv2v_reg,
  snoop_word_o_100_sv2v_reg,snoop_word_o_99_sv2v_reg,snoop_word_o_98_sv2v_reg,
  snoop_word_o_97_sv2v_reg,snoop_word_o_96_sv2v_reg,snoop_word_o_95_sv2v_reg,
  snoop_word_o_94_sv2v_reg,snoop_word_o_93_sv2v_reg,snoop_word_o_92_sv2v_reg,snoop_word_o_91_sv2v_reg,
  snoop_word_o_90_sv2v_reg,snoop_word_o_89_sv2v_reg,snoop_word_o_88_sv2v_reg,
  snoop_word_o_87_sv2v_reg,snoop_word_o_86_sv2v_reg,snoop_word_o_85_sv2v_reg,
  snoop_word_o_84_sv2v_reg,snoop_word_o_83_sv2v_reg,snoop_word_o_82_sv2v_reg,
  snoop_word_o_81_sv2v_reg,snoop_word_o_80_sv2v_reg,snoop_word_o_79_sv2v_reg,
  snoop_word_o_78_sv2v_reg,snoop_word_o_77_sv2v_reg,snoop_word_o_76_sv2v_reg,snoop_word_o_75_sv2v_reg,
  snoop_word_o_74_sv2v_reg,snoop_word_o_73_sv2v_reg,snoop_word_o_72_sv2v_reg,
  snoop_word_o_71_sv2v_reg,snoop_word_o_70_sv2v_reg,snoop_word_o_69_sv2v_reg,
  snoop_word_o_68_sv2v_reg,snoop_word_o_67_sv2v_reg,snoop_word_o_66_sv2v_reg,
  snoop_word_o_65_sv2v_reg,snoop_word_o_64_sv2v_reg,snoop_word_o_63_sv2v_reg,
  snoop_word_o_62_sv2v_reg,snoop_word_o_61_sv2v_reg,snoop_word_o_60_sv2v_reg,snoop_word_o_59_sv2v_reg,
  snoop_word_o_58_sv2v_reg,snoop_word_o_57_sv2v_reg,snoop_word_o_56_sv2v_reg,
  snoop_word_o_55_sv2v_reg,snoop_word_o_54_sv2v_reg,snoop_word_o_53_sv2v_reg,
  snoop_word_o_52_sv2v_reg,snoop_word_o_51_sv2v_reg,snoop_word_o_50_sv2v_reg,
  snoop_word_o_49_sv2v_reg,snoop_word_o_48_sv2v_reg,snoop_word_o_47_sv2v_reg,
  snoop_word_o_46_sv2v_reg,snoop_word_o_45_sv2v_reg,snoop_word_o_44_sv2v_reg,snoop_word_o_43_sv2v_reg,
  snoop_word_o_42_sv2v_reg,snoop_word_o_41_sv2v_reg,snoop_word_o_40_sv2v_reg,
  snoop_word_o_39_sv2v_reg,snoop_word_o_38_sv2v_reg,snoop_word_o_37_sv2v_reg,
  snoop_word_o_36_sv2v_reg,snoop_word_o_35_sv2v_reg,snoop_word_o_34_sv2v_reg,
  snoop_word_o_33_sv2v_reg,snoop_word_o_32_sv2v_reg,snoop_word_o_31_sv2v_reg,
  snoop_word_o_30_sv2v_reg,snoop_word_o_29_sv2v_reg,snoop_word_o_28_sv2v_reg,snoop_word_o_27_sv2v_reg,
  snoop_word_o_26_sv2v_reg,snoop_word_o_25_sv2v_reg,snoop_word_o_24_sv2v_reg,
  snoop_word_o_23_sv2v_reg,snoop_word_o_22_sv2v_reg,snoop_word_o_21_sv2v_reg,
  snoop_word_o_20_sv2v_reg,snoop_word_o_19_sv2v_reg,snoop_word_o_18_sv2v_reg,
  snoop_word_o_17_sv2v_reg,snoop_word_o_16_sv2v_reg,snoop_word_o_15_sv2v_reg,
  snoop_word_o_14_sv2v_reg,snoop_word_o_13_sv2v_reg,snoop_word_o_12_sv2v_reg,snoop_word_o_11_sv2v_reg,
  snoop_word_o_10_sv2v_reg,snoop_word_o_9_sv2v_reg,snoop_word_o_8_sv2v_reg,
  snoop_word_o_7_sv2v_reg,snoop_word_o_6_sv2v_reg,snoop_word_o_5_sv2v_reg,
  snoop_word_o_4_sv2v_reg,snoop_word_o_3_sv2v_reg,snoop_word_o_2_sv2v_reg,snoop_word_o_1_sv2v_reg,
  snoop_word_o_0_sv2v_reg;
  assign track_mem_data_r[31] = track_mem_data_r_31_sv2v_reg;
  assign track_mem_data_r[30] = track_mem_data_r_30_sv2v_reg;
  assign track_mem_data_r[29] = track_mem_data_r_29_sv2v_reg;
  assign track_mem_data_r[28] = track_mem_data_r_28_sv2v_reg;
  assign track_mem_data_r[27] = track_mem_data_r_27_sv2v_reg;
  assign track_mem_data_r[26] = track_mem_data_r_26_sv2v_reg;
  assign track_mem_data_r[25] = track_mem_data_r_25_sv2v_reg;
  assign track_mem_data_r[24] = track_mem_data_r_24_sv2v_reg;
  assign track_mem_data_r[23] = track_mem_data_r_23_sv2v_reg;
  assign track_mem_data_r[22] = track_mem_data_r_22_sv2v_reg;
  assign track_mem_data_r[21] = track_mem_data_r_21_sv2v_reg;
  assign track_mem_data_r[20] = track_mem_data_r_20_sv2v_reg;
  assign track_mem_data_r[19] = track_mem_data_r_19_sv2v_reg;
  assign track_mem_data_r[18] = track_mem_data_r_18_sv2v_reg;
  assign track_mem_data_r[17] = track_mem_data_r_17_sv2v_reg;
  assign track_mem_data_r[16] = track_mem_data_r_16_sv2v_reg;
  assign track_mem_data_r[15] = track_mem_data_r_15_sv2v_reg;
  assign track_mem_data_r[14] = track_mem_data_r_14_sv2v_reg;
  assign track_mem_data_r[13] = track_mem_data_r_13_sv2v_reg;
  assign track_mem_data_r[12] = track_mem_data_r_12_sv2v_reg;
  assign track_mem_data_r[11] = track_mem_data_r_11_sv2v_reg;
  assign track_mem_data_r[10] = track_mem_data_r_10_sv2v_reg;
  assign track_mem_data_r[9] = track_mem_data_r_9_sv2v_reg;
  assign track_mem_data_r[8] = track_mem_data_r_8_sv2v_reg;
  assign track_mem_data_r[7] = track_mem_data_r_7_sv2v_reg;
  assign track_mem_data_r[6] = track_mem_data_r_6_sv2v_reg;
  assign track_mem_data_r[5] = track_mem_data_r_5_sv2v_reg;
  assign track_mem_data_r[4] = track_mem_data_r_4_sv2v_reg;
  assign track_mem_data_r[3] = track_mem_data_r_3_sv2v_reg;
  assign track_mem_data_r[2] = track_mem_data_r_2_sv2v_reg;
  assign track_mem_data_r[1] = track_mem_data_r_1_sv2v_reg;
  assign track_mem_data_r[0] = track_mem_data_r_0_sv2v_reg;
  assign dma_state_r[1] = dma_state_r_1_sv2v_reg;
  assign dma_state_r[0] = dma_state_r_0_sv2v_reg;
  assign snoop_word_o[127] = snoop_word_o_127_sv2v_reg;
  assign snoop_word_o[126] = snoop_word_o_126_sv2v_reg;
  assign snoop_word_o[125] = snoop_word_o_125_sv2v_reg;
  assign snoop_word_o[124] = snoop_word_o_124_sv2v_reg;
  assign snoop_word_o[123] = snoop_word_o_123_sv2v_reg;
  assign snoop_word_o[122] = snoop_word_o_122_sv2v_reg;
  assign snoop_word_o[121] = snoop_word_o_121_sv2v_reg;
  assign snoop_word_o[120] = snoop_word_o_120_sv2v_reg;
  assign snoop_word_o[119] = snoop_word_o_119_sv2v_reg;
  assign snoop_word_o[118] = snoop_word_o_118_sv2v_reg;
  assign snoop_word_o[117] = snoop_word_o_117_sv2v_reg;
  assign snoop_word_o[116] = snoop_word_o_116_sv2v_reg;
  assign snoop_word_o[115] = snoop_word_o_115_sv2v_reg;
  assign snoop_word_o[114] = snoop_word_o_114_sv2v_reg;
  assign snoop_word_o[113] = snoop_word_o_113_sv2v_reg;
  assign snoop_word_o[112] = snoop_word_o_112_sv2v_reg;
  assign snoop_word_o[111] = snoop_word_o_111_sv2v_reg;
  assign snoop_word_o[110] = snoop_word_o_110_sv2v_reg;
  assign snoop_word_o[109] = snoop_word_o_109_sv2v_reg;
  assign snoop_word_o[108] = snoop_word_o_108_sv2v_reg;
  assign snoop_word_o[107] = snoop_word_o_107_sv2v_reg;
  assign snoop_word_o[106] = snoop_word_o_106_sv2v_reg;
  assign snoop_word_o[105] = snoop_word_o_105_sv2v_reg;
  assign snoop_word_o[104] = snoop_word_o_104_sv2v_reg;
  assign snoop_word_o[103] = snoop_word_o_103_sv2v_reg;
  assign snoop_word_o[102] = snoop_word_o_102_sv2v_reg;
  assign snoop_word_o[101] = snoop_word_o_101_sv2v_reg;
  assign snoop_word_o[100] = snoop_word_o_100_sv2v_reg;
  assign snoop_word_o[99] = snoop_word_o_99_sv2v_reg;
  assign snoop_word_o[98] = snoop_word_o_98_sv2v_reg;
  assign snoop_word_o[97] = snoop_word_o_97_sv2v_reg;
  assign snoop_word_o[96] = snoop_word_o_96_sv2v_reg;
  assign snoop_word_o[95] = snoop_word_o_95_sv2v_reg;
  assign snoop_word_o[94] = snoop_word_o_94_sv2v_reg;
  assign snoop_word_o[93] = snoop_word_o_93_sv2v_reg;
  assign snoop_word_o[92] = snoop_word_o_92_sv2v_reg;
  assign snoop_word_o[91] = snoop_word_o_91_sv2v_reg;
  assign snoop_word_o[90] = snoop_word_o_90_sv2v_reg;
  assign snoop_word_o[89] = snoop_word_o_89_sv2v_reg;
  assign snoop_word_o[88] = snoop_word_o_88_sv2v_reg;
  assign snoop_word_o[87] = snoop_word_o_87_sv2v_reg;
  assign snoop_word_o[86] = snoop_word_o_86_sv2v_reg;
  assign snoop_word_o[85] = snoop_word_o_85_sv2v_reg;
  assign snoop_word_o[84] = snoop_word_o_84_sv2v_reg;
  assign snoop_word_o[83] = snoop_word_o_83_sv2v_reg;
  assign snoop_word_o[82] = snoop_word_o_82_sv2v_reg;
  assign snoop_word_o[81] = snoop_word_o_81_sv2v_reg;
  assign snoop_word_o[80] = snoop_word_o_80_sv2v_reg;
  assign snoop_word_o[79] = snoop_word_o_79_sv2v_reg;
  assign snoop_word_o[78] = snoop_word_o_78_sv2v_reg;
  assign snoop_word_o[77] = snoop_word_o_77_sv2v_reg;
  assign snoop_word_o[76] = snoop_word_o_76_sv2v_reg;
  assign snoop_word_o[75] = snoop_word_o_75_sv2v_reg;
  assign snoop_word_o[74] = snoop_word_o_74_sv2v_reg;
  assign snoop_word_o[73] = snoop_word_o_73_sv2v_reg;
  assign snoop_word_o[72] = snoop_word_o_72_sv2v_reg;
  assign snoop_word_o[71] = snoop_word_o_71_sv2v_reg;
  assign snoop_word_o[70] = snoop_word_o_70_sv2v_reg;
  assign snoop_word_o[69] = snoop_word_o_69_sv2v_reg;
  assign snoop_word_o[68] = snoop_word_o_68_sv2v_reg;
  assign snoop_word_o[67] = snoop_word_o_67_sv2v_reg;
  assign snoop_word_o[66] = snoop_word_o_66_sv2v_reg;
  assign snoop_word_o[65] = snoop_word_o_65_sv2v_reg;
  assign snoop_word_o[64] = snoop_word_o_64_sv2v_reg;
  assign snoop_word_o[63] = snoop_word_o_63_sv2v_reg;
  assign snoop_word_o[62] = snoop_word_o_62_sv2v_reg;
  assign snoop_word_o[61] = snoop_word_o_61_sv2v_reg;
  assign snoop_word_o[60] = snoop_word_o_60_sv2v_reg;
  assign snoop_word_o[59] = snoop_word_o_59_sv2v_reg;
  assign snoop_word_o[58] = snoop_word_o_58_sv2v_reg;
  assign snoop_word_o[57] = snoop_word_o_57_sv2v_reg;
  assign snoop_word_o[56] = snoop_word_o_56_sv2v_reg;
  assign snoop_word_o[55] = snoop_word_o_55_sv2v_reg;
  assign snoop_word_o[54] = snoop_word_o_54_sv2v_reg;
  assign snoop_word_o[53] = snoop_word_o_53_sv2v_reg;
  assign snoop_word_o[52] = snoop_word_o_52_sv2v_reg;
  assign snoop_word_o[51] = snoop_word_o_51_sv2v_reg;
  assign snoop_word_o[50] = snoop_word_o_50_sv2v_reg;
  assign snoop_word_o[49] = snoop_word_o_49_sv2v_reg;
  assign snoop_word_o[48] = snoop_word_o_48_sv2v_reg;
  assign snoop_word_o[47] = snoop_word_o_47_sv2v_reg;
  assign snoop_word_o[46] = snoop_word_o_46_sv2v_reg;
  assign snoop_word_o[45] = snoop_word_o_45_sv2v_reg;
  assign snoop_word_o[44] = snoop_word_o_44_sv2v_reg;
  assign snoop_word_o[43] = snoop_word_o_43_sv2v_reg;
  assign snoop_word_o[42] = snoop_word_o_42_sv2v_reg;
  assign snoop_word_o[41] = snoop_word_o_41_sv2v_reg;
  assign snoop_word_o[40] = snoop_word_o_40_sv2v_reg;
  assign snoop_word_o[39] = snoop_word_o_39_sv2v_reg;
  assign snoop_word_o[38] = snoop_word_o_38_sv2v_reg;
  assign snoop_word_o[37] = snoop_word_o_37_sv2v_reg;
  assign snoop_word_o[36] = snoop_word_o_36_sv2v_reg;
  assign snoop_word_o[35] = snoop_word_o_35_sv2v_reg;
  assign snoop_word_o[34] = snoop_word_o_34_sv2v_reg;
  assign snoop_word_o[33] = snoop_word_o_33_sv2v_reg;
  assign snoop_word_o[32] = snoop_word_o_32_sv2v_reg;
  assign snoop_word_o[31] = snoop_word_o_31_sv2v_reg;
  assign snoop_word_o[30] = snoop_word_o_30_sv2v_reg;
  assign snoop_word_o[29] = snoop_word_o_29_sv2v_reg;
  assign snoop_word_o[28] = snoop_word_o_28_sv2v_reg;
  assign snoop_word_o[27] = snoop_word_o_27_sv2v_reg;
  assign snoop_word_o[26] = snoop_word_o_26_sv2v_reg;
  assign snoop_word_o[25] = snoop_word_o_25_sv2v_reg;
  assign snoop_word_o[24] = snoop_word_o_24_sv2v_reg;
  assign snoop_word_o[23] = snoop_word_o_23_sv2v_reg;
  assign snoop_word_o[22] = snoop_word_o_22_sv2v_reg;
  assign snoop_word_o[21] = snoop_word_o_21_sv2v_reg;
  assign snoop_word_o[20] = snoop_word_o_20_sv2v_reg;
  assign snoop_word_o[19] = snoop_word_o_19_sv2v_reg;
  assign snoop_word_o[18] = snoop_word_o_18_sv2v_reg;
  assign snoop_word_o[17] = snoop_word_o_17_sv2v_reg;
  assign snoop_word_o[16] = snoop_word_o_16_sv2v_reg;
  assign snoop_word_o[15] = snoop_word_o_15_sv2v_reg;
  assign snoop_word_o[14] = snoop_word_o_14_sv2v_reg;
  assign snoop_word_o[13] = snoop_word_o_13_sv2v_reg;
  assign snoop_word_o[12] = snoop_word_o_12_sv2v_reg;
  assign snoop_word_o[11] = snoop_word_o_11_sv2v_reg;
  assign snoop_word_o[10] = snoop_word_o_10_sv2v_reg;
  assign snoop_word_o[9] = snoop_word_o_9_sv2v_reg;
  assign snoop_word_o[8] = snoop_word_o_8_sv2v_reg;
  assign snoop_word_o[7] = snoop_word_o_7_sv2v_reg;
  assign snoop_word_o[6] = snoop_word_o_6_sv2v_reg;
  assign snoop_word_o[5] = snoop_word_o_5_sv2v_reg;
  assign snoop_word_o[4] = snoop_word_o_4_sv2v_reg;
  assign snoop_word_o[3] = snoop_word_o_3_sv2v_reg;
  assign snoop_word_o[2] = snoop_word_o_2_sv2v_reg;
  assign snoop_word_o[1] = snoop_word_o_1_sv2v_reg;
  assign snoop_word_o[0] = snoop_word_o_0_sv2v_reg;
  assign dma_pkt_o[4] = 1'b0;
  assign dma_pkt_o[5] = 1'b0;
  assign dma_pkt_o[6] = 1'b0;
  assign dma_pkt_o[7] = 1'b0;
  assign dma_pkt_o[8] = 1'b0;
  assign dma_pkt_o[9] = 1'b0;
  assign dma_pkt_o_36_ = dma_addr_i[32];
  assign dma_pkt_o[36] = dma_pkt_o_36_;
  assign dma_pkt_o_35_ = dma_addr_i[31];
  assign dma_pkt_o[35] = dma_pkt_o_35_;
  assign dma_pkt_o_34_ = dma_addr_i[30];
  assign dma_pkt_o[34] = dma_pkt_o_34_;
  assign dma_pkt_o_33_ = dma_addr_i[29];
  assign dma_pkt_o[33] = dma_pkt_o_33_;
  assign dma_pkt_o_32_ = dma_addr_i[28];
  assign dma_pkt_o[32] = dma_pkt_o_32_;
  assign dma_pkt_o_31_ = dma_addr_i[27];
  assign dma_pkt_o[31] = dma_pkt_o_31_;
  assign dma_pkt_o_30_ = dma_addr_i[26];
  assign dma_pkt_o[30] = dma_pkt_o_30_;
  assign dma_pkt_o_29_ = dma_addr_i[25];
  assign dma_pkt_o[29] = dma_pkt_o_29_;
  assign dma_pkt_o_28_ = dma_addr_i[24];
  assign dma_pkt_o[28] = dma_pkt_o_28_;
  assign dma_pkt_o_27_ = dma_addr_i[23];
  assign dma_pkt_o[27] = dma_pkt_o_27_;
  assign dma_pkt_o_26_ = dma_addr_i[22];
  assign dma_pkt_o[26] = dma_pkt_o_26_;
  assign dma_pkt_o_25_ = dma_addr_i[21];
  assign dma_pkt_o[25] = dma_pkt_o_25_;
  assign dma_pkt_o_24_ = dma_addr_i[20];
  assign dma_pkt_o[24] = dma_pkt_o_24_;
  assign dma_pkt_o_23_ = dma_addr_i[19];
  assign dma_pkt_o[23] = dma_pkt_o_23_;
  assign dma_pkt_o_22_ = dma_addr_i[18];
  assign dma_pkt_o[22] = dma_pkt_o_22_;
  assign dma_pkt_o_21_ = dma_addr_i[17];
  assign dma_pkt_o[21] = dma_pkt_o_21_;
  assign dma_pkt_o_20_ = dma_addr_i[16];
  assign dma_pkt_o[20] = dma_pkt_o_20_;
  assign dma_pkt_o_19_ = dma_addr_i[15];
  assign dma_pkt_o[19] = dma_pkt_o_19_;
  assign dma_pkt_o_18_ = dma_addr_i[14];
  assign dma_pkt_o[18] = dma_pkt_o_18_;
  assign dma_pkt_o_17_ = dma_addr_i[13];
  assign dma_pkt_o[17] = dma_pkt_o_17_;
  assign data_mem_addr_o_8_ = dma_addr_i[12];
  assign dma_pkt_o[16] = data_mem_addr_o_8_;
  assign data_mem_addr_o[8] = data_mem_addr_o_8_;
  assign data_mem_addr_o_7_ = dma_addr_i[11];
  assign dma_pkt_o[15] = data_mem_addr_o_7_;
  assign data_mem_addr_o[7] = data_mem_addr_o_7_;
  assign data_mem_addr_o_6_ = dma_addr_i[10];
  assign dma_pkt_o[14] = data_mem_addr_o_6_;
  assign data_mem_addr_o[6] = data_mem_addr_o_6_;
  assign data_mem_addr_o_5_ = dma_addr_i[9];
  assign dma_pkt_o[13] = data_mem_addr_o_5_;
  assign data_mem_addr_o[5] = data_mem_addr_o_5_;
  assign data_mem_addr_o_4_ = dma_addr_i[8];
  assign dma_pkt_o[12] = data_mem_addr_o_4_;
  assign data_mem_addr_o[4] = data_mem_addr_o_4_;
  assign data_mem_addr_o_3_ = dma_addr_i[7];
  assign dma_pkt_o[11] = data_mem_addr_o_3_;
  assign data_mem_addr_o[3] = data_mem_addr_o_3_;
  assign data_mem_addr_o_2_ = dma_addr_i[6];
  assign dma_pkt_o[10] = data_mem_addr_o_2_;
  assign data_mem_addr_o[2] = data_mem_addr_o_2_;
  assign data_mem_data_o[127] = data_mem_data_o_7__127_;
  assign data_mem_data_o[255] = data_mem_data_o_7__127_;
  assign data_mem_data_o[383] = data_mem_data_o_7__127_;
  assign data_mem_data_o[511] = data_mem_data_o_7__127_;
  assign data_mem_data_o[639] = data_mem_data_o_7__127_;
  assign data_mem_data_o[767] = data_mem_data_o_7__127_;
  assign data_mem_data_o[895] = data_mem_data_o_7__127_;
  assign data_mem_data_o[1023] = data_mem_data_o_7__127_;
  assign data_mem_data_o[126] = data_mem_data_o_7__126_;
  assign data_mem_data_o[254] = data_mem_data_o_7__126_;
  assign data_mem_data_o[382] = data_mem_data_o_7__126_;
  assign data_mem_data_o[510] = data_mem_data_o_7__126_;
  assign data_mem_data_o[638] = data_mem_data_o_7__126_;
  assign data_mem_data_o[766] = data_mem_data_o_7__126_;
  assign data_mem_data_o[894] = data_mem_data_o_7__126_;
  assign data_mem_data_o[1022] = data_mem_data_o_7__126_;
  assign data_mem_data_o[125] = data_mem_data_o_7__125_;
  assign data_mem_data_o[253] = data_mem_data_o_7__125_;
  assign data_mem_data_o[381] = data_mem_data_o_7__125_;
  assign data_mem_data_o[509] = data_mem_data_o_7__125_;
  assign data_mem_data_o[637] = data_mem_data_o_7__125_;
  assign data_mem_data_o[765] = data_mem_data_o_7__125_;
  assign data_mem_data_o[893] = data_mem_data_o_7__125_;
  assign data_mem_data_o[1021] = data_mem_data_o_7__125_;
  assign data_mem_data_o[124] = data_mem_data_o_7__124_;
  assign data_mem_data_o[252] = data_mem_data_o_7__124_;
  assign data_mem_data_o[380] = data_mem_data_o_7__124_;
  assign data_mem_data_o[508] = data_mem_data_o_7__124_;
  assign data_mem_data_o[636] = data_mem_data_o_7__124_;
  assign data_mem_data_o[764] = data_mem_data_o_7__124_;
  assign data_mem_data_o[892] = data_mem_data_o_7__124_;
  assign data_mem_data_o[1020] = data_mem_data_o_7__124_;
  assign data_mem_data_o[123] = data_mem_data_o_7__123_;
  assign data_mem_data_o[251] = data_mem_data_o_7__123_;
  assign data_mem_data_o[379] = data_mem_data_o_7__123_;
  assign data_mem_data_o[507] = data_mem_data_o_7__123_;
  assign data_mem_data_o[635] = data_mem_data_o_7__123_;
  assign data_mem_data_o[763] = data_mem_data_o_7__123_;
  assign data_mem_data_o[891] = data_mem_data_o_7__123_;
  assign data_mem_data_o[1019] = data_mem_data_o_7__123_;
  assign data_mem_data_o[122] = data_mem_data_o_7__122_;
  assign data_mem_data_o[250] = data_mem_data_o_7__122_;
  assign data_mem_data_o[378] = data_mem_data_o_7__122_;
  assign data_mem_data_o[506] = data_mem_data_o_7__122_;
  assign data_mem_data_o[634] = data_mem_data_o_7__122_;
  assign data_mem_data_o[762] = data_mem_data_o_7__122_;
  assign data_mem_data_o[890] = data_mem_data_o_7__122_;
  assign data_mem_data_o[1018] = data_mem_data_o_7__122_;
  assign data_mem_data_o[121] = data_mem_data_o_7__121_;
  assign data_mem_data_o[249] = data_mem_data_o_7__121_;
  assign data_mem_data_o[377] = data_mem_data_o_7__121_;
  assign data_mem_data_o[505] = data_mem_data_o_7__121_;
  assign data_mem_data_o[633] = data_mem_data_o_7__121_;
  assign data_mem_data_o[761] = data_mem_data_o_7__121_;
  assign data_mem_data_o[889] = data_mem_data_o_7__121_;
  assign data_mem_data_o[1017] = data_mem_data_o_7__121_;
  assign data_mem_data_o[120] = data_mem_data_o_7__120_;
  assign data_mem_data_o[248] = data_mem_data_o_7__120_;
  assign data_mem_data_o[376] = data_mem_data_o_7__120_;
  assign data_mem_data_o[504] = data_mem_data_o_7__120_;
  assign data_mem_data_o[632] = data_mem_data_o_7__120_;
  assign data_mem_data_o[760] = data_mem_data_o_7__120_;
  assign data_mem_data_o[888] = data_mem_data_o_7__120_;
  assign data_mem_data_o[1016] = data_mem_data_o_7__120_;
  assign data_mem_data_o[119] = data_mem_data_o_7__119_;
  assign data_mem_data_o[247] = data_mem_data_o_7__119_;
  assign data_mem_data_o[375] = data_mem_data_o_7__119_;
  assign data_mem_data_o[503] = data_mem_data_o_7__119_;
  assign data_mem_data_o[631] = data_mem_data_o_7__119_;
  assign data_mem_data_o[759] = data_mem_data_o_7__119_;
  assign data_mem_data_o[887] = data_mem_data_o_7__119_;
  assign data_mem_data_o[1015] = data_mem_data_o_7__119_;
  assign data_mem_data_o[118] = data_mem_data_o_7__118_;
  assign data_mem_data_o[246] = data_mem_data_o_7__118_;
  assign data_mem_data_o[374] = data_mem_data_o_7__118_;
  assign data_mem_data_o[502] = data_mem_data_o_7__118_;
  assign data_mem_data_o[630] = data_mem_data_o_7__118_;
  assign data_mem_data_o[758] = data_mem_data_o_7__118_;
  assign data_mem_data_o[886] = data_mem_data_o_7__118_;
  assign data_mem_data_o[1014] = data_mem_data_o_7__118_;
  assign data_mem_data_o[117] = data_mem_data_o_7__117_;
  assign data_mem_data_o[245] = data_mem_data_o_7__117_;
  assign data_mem_data_o[373] = data_mem_data_o_7__117_;
  assign data_mem_data_o[501] = data_mem_data_o_7__117_;
  assign data_mem_data_o[629] = data_mem_data_o_7__117_;
  assign data_mem_data_o[757] = data_mem_data_o_7__117_;
  assign data_mem_data_o[885] = data_mem_data_o_7__117_;
  assign data_mem_data_o[1013] = data_mem_data_o_7__117_;
  assign data_mem_data_o[116] = data_mem_data_o_7__116_;
  assign data_mem_data_o[244] = data_mem_data_o_7__116_;
  assign data_mem_data_o[372] = data_mem_data_o_7__116_;
  assign data_mem_data_o[500] = data_mem_data_o_7__116_;
  assign data_mem_data_o[628] = data_mem_data_o_7__116_;
  assign data_mem_data_o[756] = data_mem_data_o_7__116_;
  assign data_mem_data_o[884] = data_mem_data_o_7__116_;
  assign data_mem_data_o[1012] = data_mem_data_o_7__116_;
  assign data_mem_data_o[115] = data_mem_data_o_7__115_;
  assign data_mem_data_o[243] = data_mem_data_o_7__115_;
  assign data_mem_data_o[371] = data_mem_data_o_7__115_;
  assign data_mem_data_o[499] = data_mem_data_o_7__115_;
  assign data_mem_data_o[627] = data_mem_data_o_7__115_;
  assign data_mem_data_o[755] = data_mem_data_o_7__115_;
  assign data_mem_data_o[883] = data_mem_data_o_7__115_;
  assign data_mem_data_o[1011] = data_mem_data_o_7__115_;
  assign data_mem_data_o[114] = data_mem_data_o_7__114_;
  assign data_mem_data_o[242] = data_mem_data_o_7__114_;
  assign data_mem_data_o[370] = data_mem_data_o_7__114_;
  assign data_mem_data_o[498] = data_mem_data_o_7__114_;
  assign data_mem_data_o[626] = data_mem_data_o_7__114_;
  assign data_mem_data_o[754] = data_mem_data_o_7__114_;
  assign data_mem_data_o[882] = data_mem_data_o_7__114_;
  assign data_mem_data_o[1010] = data_mem_data_o_7__114_;
  assign data_mem_data_o[113] = data_mem_data_o_7__113_;
  assign data_mem_data_o[241] = data_mem_data_o_7__113_;
  assign data_mem_data_o[369] = data_mem_data_o_7__113_;
  assign data_mem_data_o[497] = data_mem_data_o_7__113_;
  assign data_mem_data_o[625] = data_mem_data_o_7__113_;
  assign data_mem_data_o[753] = data_mem_data_o_7__113_;
  assign data_mem_data_o[881] = data_mem_data_o_7__113_;
  assign data_mem_data_o[1009] = data_mem_data_o_7__113_;
  assign data_mem_data_o[112] = data_mem_data_o_7__112_;
  assign data_mem_data_o[240] = data_mem_data_o_7__112_;
  assign data_mem_data_o[368] = data_mem_data_o_7__112_;
  assign data_mem_data_o[496] = data_mem_data_o_7__112_;
  assign data_mem_data_o[624] = data_mem_data_o_7__112_;
  assign data_mem_data_o[752] = data_mem_data_o_7__112_;
  assign data_mem_data_o[880] = data_mem_data_o_7__112_;
  assign data_mem_data_o[1008] = data_mem_data_o_7__112_;
  assign data_mem_data_o[111] = data_mem_data_o_7__111_;
  assign data_mem_data_o[239] = data_mem_data_o_7__111_;
  assign data_mem_data_o[367] = data_mem_data_o_7__111_;
  assign data_mem_data_o[495] = data_mem_data_o_7__111_;
  assign data_mem_data_o[623] = data_mem_data_o_7__111_;
  assign data_mem_data_o[751] = data_mem_data_o_7__111_;
  assign data_mem_data_o[879] = data_mem_data_o_7__111_;
  assign data_mem_data_o[1007] = data_mem_data_o_7__111_;
  assign data_mem_data_o[110] = data_mem_data_o_7__110_;
  assign data_mem_data_o[238] = data_mem_data_o_7__110_;
  assign data_mem_data_o[366] = data_mem_data_o_7__110_;
  assign data_mem_data_o[494] = data_mem_data_o_7__110_;
  assign data_mem_data_o[622] = data_mem_data_o_7__110_;
  assign data_mem_data_o[750] = data_mem_data_o_7__110_;
  assign data_mem_data_o[878] = data_mem_data_o_7__110_;
  assign data_mem_data_o[1006] = data_mem_data_o_7__110_;
  assign data_mem_data_o[109] = data_mem_data_o_7__109_;
  assign data_mem_data_o[237] = data_mem_data_o_7__109_;
  assign data_mem_data_o[365] = data_mem_data_o_7__109_;
  assign data_mem_data_o[493] = data_mem_data_o_7__109_;
  assign data_mem_data_o[621] = data_mem_data_o_7__109_;
  assign data_mem_data_o[749] = data_mem_data_o_7__109_;
  assign data_mem_data_o[877] = data_mem_data_o_7__109_;
  assign data_mem_data_o[1005] = data_mem_data_o_7__109_;
  assign data_mem_data_o[108] = data_mem_data_o_7__108_;
  assign data_mem_data_o[236] = data_mem_data_o_7__108_;
  assign data_mem_data_o[364] = data_mem_data_o_7__108_;
  assign data_mem_data_o[492] = data_mem_data_o_7__108_;
  assign data_mem_data_o[620] = data_mem_data_o_7__108_;
  assign data_mem_data_o[748] = data_mem_data_o_7__108_;
  assign data_mem_data_o[876] = data_mem_data_o_7__108_;
  assign data_mem_data_o[1004] = data_mem_data_o_7__108_;
  assign data_mem_data_o[107] = data_mem_data_o_7__107_;
  assign data_mem_data_o[235] = data_mem_data_o_7__107_;
  assign data_mem_data_o[363] = data_mem_data_o_7__107_;
  assign data_mem_data_o[491] = data_mem_data_o_7__107_;
  assign data_mem_data_o[619] = data_mem_data_o_7__107_;
  assign data_mem_data_o[747] = data_mem_data_o_7__107_;
  assign data_mem_data_o[875] = data_mem_data_o_7__107_;
  assign data_mem_data_o[1003] = data_mem_data_o_7__107_;
  assign data_mem_data_o[106] = data_mem_data_o_7__106_;
  assign data_mem_data_o[234] = data_mem_data_o_7__106_;
  assign data_mem_data_o[362] = data_mem_data_o_7__106_;
  assign data_mem_data_o[490] = data_mem_data_o_7__106_;
  assign data_mem_data_o[618] = data_mem_data_o_7__106_;
  assign data_mem_data_o[746] = data_mem_data_o_7__106_;
  assign data_mem_data_o[874] = data_mem_data_o_7__106_;
  assign data_mem_data_o[1002] = data_mem_data_o_7__106_;
  assign data_mem_data_o[105] = data_mem_data_o_7__105_;
  assign data_mem_data_o[233] = data_mem_data_o_7__105_;
  assign data_mem_data_o[361] = data_mem_data_o_7__105_;
  assign data_mem_data_o[489] = data_mem_data_o_7__105_;
  assign data_mem_data_o[617] = data_mem_data_o_7__105_;
  assign data_mem_data_o[745] = data_mem_data_o_7__105_;
  assign data_mem_data_o[873] = data_mem_data_o_7__105_;
  assign data_mem_data_o[1001] = data_mem_data_o_7__105_;
  assign data_mem_data_o[104] = data_mem_data_o_7__104_;
  assign data_mem_data_o[232] = data_mem_data_o_7__104_;
  assign data_mem_data_o[360] = data_mem_data_o_7__104_;
  assign data_mem_data_o[488] = data_mem_data_o_7__104_;
  assign data_mem_data_o[616] = data_mem_data_o_7__104_;
  assign data_mem_data_o[744] = data_mem_data_o_7__104_;
  assign data_mem_data_o[872] = data_mem_data_o_7__104_;
  assign data_mem_data_o[1000] = data_mem_data_o_7__104_;
  assign data_mem_data_o[103] = data_mem_data_o_7__103_;
  assign data_mem_data_o[231] = data_mem_data_o_7__103_;
  assign data_mem_data_o[359] = data_mem_data_o_7__103_;
  assign data_mem_data_o[487] = data_mem_data_o_7__103_;
  assign data_mem_data_o[615] = data_mem_data_o_7__103_;
  assign data_mem_data_o[743] = data_mem_data_o_7__103_;
  assign data_mem_data_o[871] = data_mem_data_o_7__103_;
  assign data_mem_data_o[999] = data_mem_data_o_7__103_;
  assign data_mem_data_o[102] = data_mem_data_o_7__102_;
  assign data_mem_data_o[230] = data_mem_data_o_7__102_;
  assign data_mem_data_o[358] = data_mem_data_o_7__102_;
  assign data_mem_data_o[486] = data_mem_data_o_7__102_;
  assign data_mem_data_o[614] = data_mem_data_o_7__102_;
  assign data_mem_data_o[742] = data_mem_data_o_7__102_;
  assign data_mem_data_o[870] = data_mem_data_o_7__102_;
  assign data_mem_data_o[998] = data_mem_data_o_7__102_;
  assign data_mem_data_o[101] = data_mem_data_o_7__101_;
  assign data_mem_data_o[229] = data_mem_data_o_7__101_;
  assign data_mem_data_o[357] = data_mem_data_o_7__101_;
  assign data_mem_data_o[485] = data_mem_data_o_7__101_;
  assign data_mem_data_o[613] = data_mem_data_o_7__101_;
  assign data_mem_data_o[741] = data_mem_data_o_7__101_;
  assign data_mem_data_o[869] = data_mem_data_o_7__101_;
  assign data_mem_data_o[997] = data_mem_data_o_7__101_;
  assign data_mem_data_o[100] = data_mem_data_o_7__100_;
  assign data_mem_data_o[228] = data_mem_data_o_7__100_;
  assign data_mem_data_o[356] = data_mem_data_o_7__100_;
  assign data_mem_data_o[484] = data_mem_data_o_7__100_;
  assign data_mem_data_o[612] = data_mem_data_o_7__100_;
  assign data_mem_data_o[740] = data_mem_data_o_7__100_;
  assign data_mem_data_o[868] = data_mem_data_o_7__100_;
  assign data_mem_data_o[996] = data_mem_data_o_7__100_;
  assign data_mem_data_o[99] = data_mem_data_o_7__99_;
  assign data_mem_data_o[227] = data_mem_data_o_7__99_;
  assign data_mem_data_o[355] = data_mem_data_o_7__99_;
  assign data_mem_data_o[483] = data_mem_data_o_7__99_;
  assign data_mem_data_o[611] = data_mem_data_o_7__99_;
  assign data_mem_data_o[739] = data_mem_data_o_7__99_;
  assign data_mem_data_o[867] = data_mem_data_o_7__99_;
  assign data_mem_data_o[995] = data_mem_data_o_7__99_;
  assign data_mem_data_o[98] = data_mem_data_o_7__98_;
  assign data_mem_data_o[226] = data_mem_data_o_7__98_;
  assign data_mem_data_o[354] = data_mem_data_o_7__98_;
  assign data_mem_data_o[482] = data_mem_data_o_7__98_;
  assign data_mem_data_o[610] = data_mem_data_o_7__98_;
  assign data_mem_data_o[738] = data_mem_data_o_7__98_;
  assign data_mem_data_o[866] = data_mem_data_o_7__98_;
  assign data_mem_data_o[994] = data_mem_data_o_7__98_;
  assign data_mem_data_o[97] = data_mem_data_o_7__97_;
  assign data_mem_data_o[225] = data_mem_data_o_7__97_;
  assign data_mem_data_o[353] = data_mem_data_o_7__97_;
  assign data_mem_data_o[481] = data_mem_data_o_7__97_;
  assign data_mem_data_o[609] = data_mem_data_o_7__97_;
  assign data_mem_data_o[737] = data_mem_data_o_7__97_;
  assign data_mem_data_o[865] = data_mem_data_o_7__97_;
  assign data_mem_data_o[993] = data_mem_data_o_7__97_;
  assign data_mem_data_o[96] = data_mem_data_o_7__96_;
  assign data_mem_data_o[224] = data_mem_data_o_7__96_;
  assign data_mem_data_o[352] = data_mem_data_o_7__96_;
  assign data_mem_data_o[480] = data_mem_data_o_7__96_;
  assign data_mem_data_o[608] = data_mem_data_o_7__96_;
  assign data_mem_data_o[736] = data_mem_data_o_7__96_;
  assign data_mem_data_o[864] = data_mem_data_o_7__96_;
  assign data_mem_data_o[992] = data_mem_data_o_7__96_;
  assign data_mem_data_o[95] = data_mem_data_o_7__95_;
  assign data_mem_data_o[223] = data_mem_data_o_7__95_;
  assign data_mem_data_o[351] = data_mem_data_o_7__95_;
  assign data_mem_data_o[479] = data_mem_data_o_7__95_;
  assign data_mem_data_o[607] = data_mem_data_o_7__95_;
  assign data_mem_data_o[735] = data_mem_data_o_7__95_;
  assign data_mem_data_o[863] = data_mem_data_o_7__95_;
  assign data_mem_data_o[991] = data_mem_data_o_7__95_;
  assign data_mem_data_o[94] = data_mem_data_o_7__94_;
  assign data_mem_data_o[222] = data_mem_data_o_7__94_;
  assign data_mem_data_o[350] = data_mem_data_o_7__94_;
  assign data_mem_data_o[478] = data_mem_data_o_7__94_;
  assign data_mem_data_o[606] = data_mem_data_o_7__94_;
  assign data_mem_data_o[734] = data_mem_data_o_7__94_;
  assign data_mem_data_o[862] = data_mem_data_o_7__94_;
  assign data_mem_data_o[990] = data_mem_data_o_7__94_;
  assign data_mem_data_o[93] = data_mem_data_o_7__93_;
  assign data_mem_data_o[221] = data_mem_data_o_7__93_;
  assign data_mem_data_o[349] = data_mem_data_o_7__93_;
  assign data_mem_data_o[477] = data_mem_data_o_7__93_;
  assign data_mem_data_o[605] = data_mem_data_o_7__93_;
  assign data_mem_data_o[733] = data_mem_data_o_7__93_;
  assign data_mem_data_o[861] = data_mem_data_o_7__93_;
  assign data_mem_data_o[989] = data_mem_data_o_7__93_;
  assign data_mem_data_o[92] = data_mem_data_o_7__92_;
  assign data_mem_data_o[220] = data_mem_data_o_7__92_;
  assign data_mem_data_o[348] = data_mem_data_o_7__92_;
  assign data_mem_data_o[476] = data_mem_data_o_7__92_;
  assign data_mem_data_o[604] = data_mem_data_o_7__92_;
  assign data_mem_data_o[732] = data_mem_data_o_7__92_;
  assign data_mem_data_o[860] = data_mem_data_o_7__92_;
  assign data_mem_data_o[988] = data_mem_data_o_7__92_;
  assign data_mem_data_o[91] = data_mem_data_o_7__91_;
  assign data_mem_data_o[219] = data_mem_data_o_7__91_;
  assign data_mem_data_o[347] = data_mem_data_o_7__91_;
  assign data_mem_data_o[475] = data_mem_data_o_7__91_;
  assign data_mem_data_o[603] = data_mem_data_o_7__91_;
  assign data_mem_data_o[731] = data_mem_data_o_7__91_;
  assign data_mem_data_o[859] = data_mem_data_o_7__91_;
  assign data_mem_data_o[987] = data_mem_data_o_7__91_;
  assign data_mem_data_o[90] = data_mem_data_o_7__90_;
  assign data_mem_data_o[218] = data_mem_data_o_7__90_;
  assign data_mem_data_o[346] = data_mem_data_o_7__90_;
  assign data_mem_data_o[474] = data_mem_data_o_7__90_;
  assign data_mem_data_o[602] = data_mem_data_o_7__90_;
  assign data_mem_data_o[730] = data_mem_data_o_7__90_;
  assign data_mem_data_o[858] = data_mem_data_o_7__90_;
  assign data_mem_data_o[986] = data_mem_data_o_7__90_;
  assign data_mem_data_o[89] = data_mem_data_o_7__89_;
  assign data_mem_data_o[217] = data_mem_data_o_7__89_;
  assign data_mem_data_o[345] = data_mem_data_o_7__89_;
  assign data_mem_data_o[473] = data_mem_data_o_7__89_;
  assign data_mem_data_o[601] = data_mem_data_o_7__89_;
  assign data_mem_data_o[729] = data_mem_data_o_7__89_;
  assign data_mem_data_o[857] = data_mem_data_o_7__89_;
  assign data_mem_data_o[985] = data_mem_data_o_7__89_;
  assign data_mem_data_o[88] = data_mem_data_o_7__88_;
  assign data_mem_data_o[216] = data_mem_data_o_7__88_;
  assign data_mem_data_o[344] = data_mem_data_o_7__88_;
  assign data_mem_data_o[472] = data_mem_data_o_7__88_;
  assign data_mem_data_o[600] = data_mem_data_o_7__88_;
  assign data_mem_data_o[728] = data_mem_data_o_7__88_;
  assign data_mem_data_o[856] = data_mem_data_o_7__88_;
  assign data_mem_data_o[984] = data_mem_data_o_7__88_;
  assign data_mem_data_o[87] = data_mem_data_o_7__87_;
  assign data_mem_data_o[215] = data_mem_data_o_7__87_;
  assign data_mem_data_o[343] = data_mem_data_o_7__87_;
  assign data_mem_data_o[471] = data_mem_data_o_7__87_;
  assign data_mem_data_o[599] = data_mem_data_o_7__87_;
  assign data_mem_data_o[727] = data_mem_data_o_7__87_;
  assign data_mem_data_o[855] = data_mem_data_o_7__87_;
  assign data_mem_data_o[983] = data_mem_data_o_7__87_;
  assign data_mem_data_o[86] = data_mem_data_o_7__86_;
  assign data_mem_data_o[214] = data_mem_data_o_7__86_;
  assign data_mem_data_o[342] = data_mem_data_o_7__86_;
  assign data_mem_data_o[470] = data_mem_data_o_7__86_;
  assign data_mem_data_o[598] = data_mem_data_o_7__86_;
  assign data_mem_data_o[726] = data_mem_data_o_7__86_;
  assign data_mem_data_o[854] = data_mem_data_o_7__86_;
  assign data_mem_data_o[982] = data_mem_data_o_7__86_;
  assign data_mem_data_o[85] = data_mem_data_o_7__85_;
  assign data_mem_data_o[213] = data_mem_data_o_7__85_;
  assign data_mem_data_o[341] = data_mem_data_o_7__85_;
  assign data_mem_data_o[469] = data_mem_data_o_7__85_;
  assign data_mem_data_o[597] = data_mem_data_o_7__85_;
  assign data_mem_data_o[725] = data_mem_data_o_7__85_;
  assign data_mem_data_o[853] = data_mem_data_o_7__85_;
  assign data_mem_data_o[981] = data_mem_data_o_7__85_;
  assign data_mem_data_o[84] = data_mem_data_o_7__84_;
  assign data_mem_data_o[212] = data_mem_data_o_7__84_;
  assign data_mem_data_o[340] = data_mem_data_o_7__84_;
  assign data_mem_data_o[468] = data_mem_data_o_7__84_;
  assign data_mem_data_o[596] = data_mem_data_o_7__84_;
  assign data_mem_data_o[724] = data_mem_data_o_7__84_;
  assign data_mem_data_o[852] = data_mem_data_o_7__84_;
  assign data_mem_data_o[980] = data_mem_data_o_7__84_;
  assign data_mem_data_o[83] = data_mem_data_o_7__83_;
  assign data_mem_data_o[211] = data_mem_data_o_7__83_;
  assign data_mem_data_o[339] = data_mem_data_o_7__83_;
  assign data_mem_data_o[467] = data_mem_data_o_7__83_;
  assign data_mem_data_o[595] = data_mem_data_o_7__83_;
  assign data_mem_data_o[723] = data_mem_data_o_7__83_;
  assign data_mem_data_o[851] = data_mem_data_o_7__83_;
  assign data_mem_data_o[979] = data_mem_data_o_7__83_;
  assign data_mem_data_o[82] = data_mem_data_o_7__82_;
  assign data_mem_data_o[210] = data_mem_data_o_7__82_;
  assign data_mem_data_o[338] = data_mem_data_o_7__82_;
  assign data_mem_data_o[466] = data_mem_data_o_7__82_;
  assign data_mem_data_o[594] = data_mem_data_o_7__82_;
  assign data_mem_data_o[722] = data_mem_data_o_7__82_;
  assign data_mem_data_o[850] = data_mem_data_o_7__82_;
  assign data_mem_data_o[978] = data_mem_data_o_7__82_;
  assign data_mem_data_o[81] = data_mem_data_o_7__81_;
  assign data_mem_data_o[209] = data_mem_data_o_7__81_;
  assign data_mem_data_o[337] = data_mem_data_o_7__81_;
  assign data_mem_data_o[465] = data_mem_data_o_7__81_;
  assign data_mem_data_o[593] = data_mem_data_o_7__81_;
  assign data_mem_data_o[721] = data_mem_data_o_7__81_;
  assign data_mem_data_o[849] = data_mem_data_o_7__81_;
  assign data_mem_data_o[977] = data_mem_data_o_7__81_;
  assign data_mem_data_o[80] = data_mem_data_o_7__80_;
  assign data_mem_data_o[208] = data_mem_data_o_7__80_;
  assign data_mem_data_o[336] = data_mem_data_o_7__80_;
  assign data_mem_data_o[464] = data_mem_data_o_7__80_;
  assign data_mem_data_o[592] = data_mem_data_o_7__80_;
  assign data_mem_data_o[720] = data_mem_data_o_7__80_;
  assign data_mem_data_o[848] = data_mem_data_o_7__80_;
  assign data_mem_data_o[976] = data_mem_data_o_7__80_;
  assign data_mem_data_o[79] = data_mem_data_o_7__79_;
  assign data_mem_data_o[207] = data_mem_data_o_7__79_;
  assign data_mem_data_o[335] = data_mem_data_o_7__79_;
  assign data_mem_data_o[463] = data_mem_data_o_7__79_;
  assign data_mem_data_o[591] = data_mem_data_o_7__79_;
  assign data_mem_data_o[719] = data_mem_data_o_7__79_;
  assign data_mem_data_o[847] = data_mem_data_o_7__79_;
  assign data_mem_data_o[975] = data_mem_data_o_7__79_;
  assign data_mem_data_o[78] = data_mem_data_o_7__78_;
  assign data_mem_data_o[206] = data_mem_data_o_7__78_;
  assign data_mem_data_o[334] = data_mem_data_o_7__78_;
  assign data_mem_data_o[462] = data_mem_data_o_7__78_;
  assign data_mem_data_o[590] = data_mem_data_o_7__78_;
  assign data_mem_data_o[718] = data_mem_data_o_7__78_;
  assign data_mem_data_o[846] = data_mem_data_o_7__78_;
  assign data_mem_data_o[974] = data_mem_data_o_7__78_;
  assign data_mem_data_o[77] = data_mem_data_o_7__77_;
  assign data_mem_data_o[205] = data_mem_data_o_7__77_;
  assign data_mem_data_o[333] = data_mem_data_o_7__77_;
  assign data_mem_data_o[461] = data_mem_data_o_7__77_;
  assign data_mem_data_o[589] = data_mem_data_o_7__77_;
  assign data_mem_data_o[717] = data_mem_data_o_7__77_;
  assign data_mem_data_o[845] = data_mem_data_o_7__77_;
  assign data_mem_data_o[973] = data_mem_data_o_7__77_;
  assign data_mem_data_o[76] = data_mem_data_o_7__76_;
  assign data_mem_data_o[204] = data_mem_data_o_7__76_;
  assign data_mem_data_o[332] = data_mem_data_o_7__76_;
  assign data_mem_data_o[460] = data_mem_data_o_7__76_;
  assign data_mem_data_o[588] = data_mem_data_o_7__76_;
  assign data_mem_data_o[716] = data_mem_data_o_7__76_;
  assign data_mem_data_o[844] = data_mem_data_o_7__76_;
  assign data_mem_data_o[972] = data_mem_data_o_7__76_;
  assign data_mem_data_o[75] = data_mem_data_o_7__75_;
  assign data_mem_data_o[203] = data_mem_data_o_7__75_;
  assign data_mem_data_o[331] = data_mem_data_o_7__75_;
  assign data_mem_data_o[459] = data_mem_data_o_7__75_;
  assign data_mem_data_o[587] = data_mem_data_o_7__75_;
  assign data_mem_data_o[715] = data_mem_data_o_7__75_;
  assign data_mem_data_o[843] = data_mem_data_o_7__75_;
  assign data_mem_data_o[971] = data_mem_data_o_7__75_;
  assign data_mem_data_o[74] = data_mem_data_o_7__74_;
  assign data_mem_data_o[202] = data_mem_data_o_7__74_;
  assign data_mem_data_o[330] = data_mem_data_o_7__74_;
  assign data_mem_data_o[458] = data_mem_data_o_7__74_;
  assign data_mem_data_o[586] = data_mem_data_o_7__74_;
  assign data_mem_data_o[714] = data_mem_data_o_7__74_;
  assign data_mem_data_o[842] = data_mem_data_o_7__74_;
  assign data_mem_data_o[970] = data_mem_data_o_7__74_;
  assign data_mem_data_o[73] = data_mem_data_o_7__73_;
  assign data_mem_data_o[201] = data_mem_data_o_7__73_;
  assign data_mem_data_o[329] = data_mem_data_o_7__73_;
  assign data_mem_data_o[457] = data_mem_data_o_7__73_;
  assign data_mem_data_o[585] = data_mem_data_o_7__73_;
  assign data_mem_data_o[713] = data_mem_data_o_7__73_;
  assign data_mem_data_o[841] = data_mem_data_o_7__73_;
  assign data_mem_data_o[969] = data_mem_data_o_7__73_;
  assign data_mem_data_o[72] = data_mem_data_o_7__72_;
  assign data_mem_data_o[200] = data_mem_data_o_7__72_;
  assign data_mem_data_o[328] = data_mem_data_o_7__72_;
  assign data_mem_data_o[456] = data_mem_data_o_7__72_;
  assign data_mem_data_o[584] = data_mem_data_o_7__72_;
  assign data_mem_data_o[712] = data_mem_data_o_7__72_;
  assign data_mem_data_o[840] = data_mem_data_o_7__72_;
  assign data_mem_data_o[968] = data_mem_data_o_7__72_;
  assign data_mem_data_o[71] = data_mem_data_o_7__71_;
  assign data_mem_data_o[199] = data_mem_data_o_7__71_;
  assign data_mem_data_o[327] = data_mem_data_o_7__71_;
  assign data_mem_data_o[455] = data_mem_data_o_7__71_;
  assign data_mem_data_o[583] = data_mem_data_o_7__71_;
  assign data_mem_data_o[711] = data_mem_data_o_7__71_;
  assign data_mem_data_o[839] = data_mem_data_o_7__71_;
  assign data_mem_data_o[967] = data_mem_data_o_7__71_;
  assign data_mem_data_o[70] = data_mem_data_o_7__70_;
  assign data_mem_data_o[198] = data_mem_data_o_7__70_;
  assign data_mem_data_o[326] = data_mem_data_o_7__70_;
  assign data_mem_data_o[454] = data_mem_data_o_7__70_;
  assign data_mem_data_o[582] = data_mem_data_o_7__70_;
  assign data_mem_data_o[710] = data_mem_data_o_7__70_;
  assign data_mem_data_o[838] = data_mem_data_o_7__70_;
  assign data_mem_data_o[966] = data_mem_data_o_7__70_;
  assign data_mem_data_o[69] = data_mem_data_o_7__69_;
  assign data_mem_data_o[197] = data_mem_data_o_7__69_;
  assign data_mem_data_o[325] = data_mem_data_o_7__69_;
  assign data_mem_data_o[453] = data_mem_data_o_7__69_;
  assign data_mem_data_o[581] = data_mem_data_o_7__69_;
  assign data_mem_data_o[709] = data_mem_data_o_7__69_;
  assign data_mem_data_o[837] = data_mem_data_o_7__69_;
  assign data_mem_data_o[965] = data_mem_data_o_7__69_;
  assign data_mem_data_o[68] = data_mem_data_o_7__68_;
  assign data_mem_data_o[196] = data_mem_data_o_7__68_;
  assign data_mem_data_o[324] = data_mem_data_o_7__68_;
  assign data_mem_data_o[452] = data_mem_data_o_7__68_;
  assign data_mem_data_o[580] = data_mem_data_o_7__68_;
  assign data_mem_data_o[708] = data_mem_data_o_7__68_;
  assign data_mem_data_o[836] = data_mem_data_o_7__68_;
  assign data_mem_data_o[964] = data_mem_data_o_7__68_;
  assign data_mem_data_o[67] = data_mem_data_o_7__67_;
  assign data_mem_data_o[195] = data_mem_data_o_7__67_;
  assign data_mem_data_o[323] = data_mem_data_o_7__67_;
  assign data_mem_data_o[451] = data_mem_data_o_7__67_;
  assign data_mem_data_o[579] = data_mem_data_o_7__67_;
  assign data_mem_data_o[707] = data_mem_data_o_7__67_;
  assign data_mem_data_o[835] = data_mem_data_o_7__67_;
  assign data_mem_data_o[963] = data_mem_data_o_7__67_;
  assign data_mem_data_o[66] = data_mem_data_o_7__66_;
  assign data_mem_data_o[194] = data_mem_data_o_7__66_;
  assign data_mem_data_o[322] = data_mem_data_o_7__66_;
  assign data_mem_data_o[450] = data_mem_data_o_7__66_;
  assign data_mem_data_o[578] = data_mem_data_o_7__66_;
  assign data_mem_data_o[706] = data_mem_data_o_7__66_;
  assign data_mem_data_o[834] = data_mem_data_o_7__66_;
  assign data_mem_data_o[962] = data_mem_data_o_7__66_;
  assign data_mem_data_o[65] = data_mem_data_o_7__65_;
  assign data_mem_data_o[193] = data_mem_data_o_7__65_;
  assign data_mem_data_o[321] = data_mem_data_o_7__65_;
  assign data_mem_data_o[449] = data_mem_data_o_7__65_;
  assign data_mem_data_o[577] = data_mem_data_o_7__65_;
  assign data_mem_data_o[705] = data_mem_data_o_7__65_;
  assign data_mem_data_o[833] = data_mem_data_o_7__65_;
  assign data_mem_data_o[961] = data_mem_data_o_7__65_;
  assign data_mem_data_o[64] = data_mem_data_o_7__64_;
  assign data_mem_data_o[192] = data_mem_data_o_7__64_;
  assign data_mem_data_o[320] = data_mem_data_o_7__64_;
  assign data_mem_data_o[448] = data_mem_data_o_7__64_;
  assign data_mem_data_o[576] = data_mem_data_o_7__64_;
  assign data_mem_data_o[704] = data_mem_data_o_7__64_;
  assign data_mem_data_o[832] = data_mem_data_o_7__64_;
  assign data_mem_data_o[960] = data_mem_data_o_7__64_;
  assign data_mem_data_o[63] = data_mem_data_o_7__63_;
  assign data_mem_data_o[191] = data_mem_data_o_7__63_;
  assign data_mem_data_o[319] = data_mem_data_o_7__63_;
  assign data_mem_data_o[447] = data_mem_data_o_7__63_;
  assign data_mem_data_o[575] = data_mem_data_o_7__63_;
  assign data_mem_data_o[703] = data_mem_data_o_7__63_;
  assign data_mem_data_o[831] = data_mem_data_o_7__63_;
  assign data_mem_data_o[959] = data_mem_data_o_7__63_;
  assign data_mem_data_o[62] = data_mem_data_o_7__62_;
  assign data_mem_data_o[190] = data_mem_data_o_7__62_;
  assign data_mem_data_o[318] = data_mem_data_o_7__62_;
  assign data_mem_data_o[446] = data_mem_data_o_7__62_;
  assign data_mem_data_o[574] = data_mem_data_o_7__62_;
  assign data_mem_data_o[702] = data_mem_data_o_7__62_;
  assign data_mem_data_o[830] = data_mem_data_o_7__62_;
  assign data_mem_data_o[958] = data_mem_data_o_7__62_;
  assign data_mem_data_o[61] = data_mem_data_o_7__61_;
  assign data_mem_data_o[189] = data_mem_data_o_7__61_;
  assign data_mem_data_o[317] = data_mem_data_o_7__61_;
  assign data_mem_data_o[445] = data_mem_data_o_7__61_;
  assign data_mem_data_o[573] = data_mem_data_o_7__61_;
  assign data_mem_data_o[701] = data_mem_data_o_7__61_;
  assign data_mem_data_o[829] = data_mem_data_o_7__61_;
  assign data_mem_data_o[957] = data_mem_data_o_7__61_;
  assign data_mem_data_o[60] = data_mem_data_o_7__60_;
  assign data_mem_data_o[188] = data_mem_data_o_7__60_;
  assign data_mem_data_o[316] = data_mem_data_o_7__60_;
  assign data_mem_data_o[444] = data_mem_data_o_7__60_;
  assign data_mem_data_o[572] = data_mem_data_o_7__60_;
  assign data_mem_data_o[700] = data_mem_data_o_7__60_;
  assign data_mem_data_o[828] = data_mem_data_o_7__60_;
  assign data_mem_data_o[956] = data_mem_data_o_7__60_;
  assign data_mem_data_o[59] = data_mem_data_o_7__59_;
  assign data_mem_data_o[187] = data_mem_data_o_7__59_;
  assign data_mem_data_o[315] = data_mem_data_o_7__59_;
  assign data_mem_data_o[443] = data_mem_data_o_7__59_;
  assign data_mem_data_o[571] = data_mem_data_o_7__59_;
  assign data_mem_data_o[699] = data_mem_data_o_7__59_;
  assign data_mem_data_o[827] = data_mem_data_o_7__59_;
  assign data_mem_data_o[955] = data_mem_data_o_7__59_;
  assign data_mem_data_o[58] = data_mem_data_o_7__58_;
  assign data_mem_data_o[186] = data_mem_data_o_7__58_;
  assign data_mem_data_o[314] = data_mem_data_o_7__58_;
  assign data_mem_data_o[442] = data_mem_data_o_7__58_;
  assign data_mem_data_o[570] = data_mem_data_o_7__58_;
  assign data_mem_data_o[698] = data_mem_data_o_7__58_;
  assign data_mem_data_o[826] = data_mem_data_o_7__58_;
  assign data_mem_data_o[954] = data_mem_data_o_7__58_;
  assign data_mem_data_o[57] = data_mem_data_o_7__57_;
  assign data_mem_data_o[185] = data_mem_data_o_7__57_;
  assign data_mem_data_o[313] = data_mem_data_o_7__57_;
  assign data_mem_data_o[441] = data_mem_data_o_7__57_;
  assign data_mem_data_o[569] = data_mem_data_o_7__57_;
  assign data_mem_data_o[697] = data_mem_data_o_7__57_;
  assign data_mem_data_o[825] = data_mem_data_o_7__57_;
  assign data_mem_data_o[953] = data_mem_data_o_7__57_;
  assign data_mem_data_o[56] = data_mem_data_o_7__56_;
  assign data_mem_data_o[184] = data_mem_data_o_7__56_;
  assign data_mem_data_o[312] = data_mem_data_o_7__56_;
  assign data_mem_data_o[440] = data_mem_data_o_7__56_;
  assign data_mem_data_o[568] = data_mem_data_o_7__56_;
  assign data_mem_data_o[696] = data_mem_data_o_7__56_;
  assign data_mem_data_o[824] = data_mem_data_o_7__56_;
  assign data_mem_data_o[952] = data_mem_data_o_7__56_;
  assign data_mem_data_o[55] = data_mem_data_o_7__55_;
  assign data_mem_data_o[183] = data_mem_data_o_7__55_;
  assign data_mem_data_o[311] = data_mem_data_o_7__55_;
  assign data_mem_data_o[439] = data_mem_data_o_7__55_;
  assign data_mem_data_o[567] = data_mem_data_o_7__55_;
  assign data_mem_data_o[695] = data_mem_data_o_7__55_;
  assign data_mem_data_o[823] = data_mem_data_o_7__55_;
  assign data_mem_data_o[951] = data_mem_data_o_7__55_;
  assign data_mem_data_o[54] = data_mem_data_o_7__54_;
  assign data_mem_data_o[182] = data_mem_data_o_7__54_;
  assign data_mem_data_o[310] = data_mem_data_o_7__54_;
  assign data_mem_data_o[438] = data_mem_data_o_7__54_;
  assign data_mem_data_o[566] = data_mem_data_o_7__54_;
  assign data_mem_data_o[694] = data_mem_data_o_7__54_;
  assign data_mem_data_o[822] = data_mem_data_o_7__54_;
  assign data_mem_data_o[950] = data_mem_data_o_7__54_;
  assign data_mem_data_o[53] = data_mem_data_o_7__53_;
  assign data_mem_data_o[181] = data_mem_data_o_7__53_;
  assign data_mem_data_o[309] = data_mem_data_o_7__53_;
  assign data_mem_data_o[437] = data_mem_data_o_7__53_;
  assign data_mem_data_o[565] = data_mem_data_o_7__53_;
  assign data_mem_data_o[693] = data_mem_data_o_7__53_;
  assign data_mem_data_o[821] = data_mem_data_o_7__53_;
  assign data_mem_data_o[949] = data_mem_data_o_7__53_;
  assign data_mem_data_o[52] = data_mem_data_o_7__52_;
  assign data_mem_data_o[180] = data_mem_data_o_7__52_;
  assign data_mem_data_o[308] = data_mem_data_o_7__52_;
  assign data_mem_data_o[436] = data_mem_data_o_7__52_;
  assign data_mem_data_o[564] = data_mem_data_o_7__52_;
  assign data_mem_data_o[692] = data_mem_data_o_7__52_;
  assign data_mem_data_o[820] = data_mem_data_o_7__52_;
  assign data_mem_data_o[948] = data_mem_data_o_7__52_;
  assign data_mem_data_o[51] = data_mem_data_o_7__51_;
  assign data_mem_data_o[179] = data_mem_data_o_7__51_;
  assign data_mem_data_o[307] = data_mem_data_o_7__51_;
  assign data_mem_data_o[435] = data_mem_data_o_7__51_;
  assign data_mem_data_o[563] = data_mem_data_o_7__51_;
  assign data_mem_data_o[691] = data_mem_data_o_7__51_;
  assign data_mem_data_o[819] = data_mem_data_o_7__51_;
  assign data_mem_data_o[947] = data_mem_data_o_7__51_;
  assign data_mem_data_o[50] = data_mem_data_o_7__50_;
  assign data_mem_data_o[178] = data_mem_data_o_7__50_;
  assign data_mem_data_o[306] = data_mem_data_o_7__50_;
  assign data_mem_data_o[434] = data_mem_data_o_7__50_;
  assign data_mem_data_o[562] = data_mem_data_o_7__50_;
  assign data_mem_data_o[690] = data_mem_data_o_7__50_;
  assign data_mem_data_o[818] = data_mem_data_o_7__50_;
  assign data_mem_data_o[946] = data_mem_data_o_7__50_;
  assign data_mem_data_o[49] = data_mem_data_o_7__49_;
  assign data_mem_data_o[177] = data_mem_data_o_7__49_;
  assign data_mem_data_o[305] = data_mem_data_o_7__49_;
  assign data_mem_data_o[433] = data_mem_data_o_7__49_;
  assign data_mem_data_o[561] = data_mem_data_o_7__49_;
  assign data_mem_data_o[689] = data_mem_data_o_7__49_;
  assign data_mem_data_o[817] = data_mem_data_o_7__49_;
  assign data_mem_data_o[945] = data_mem_data_o_7__49_;
  assign data_mem_data_o[48] = data_mem_data_o_7__48_;
  assign data_mem_data_o[176] = data_mem_data_o_7__48_;
  assign data_mem_data_o[304] = data_mem_data_o_7__48_;
  assign data_mem_data_o[432] = data_mem_data_o_7__48_;
  assign data_mem_data_o[560] = data_mem_data_o_7__48_;
  assign data_mem_data_o[688] = data_mem_data_o_7__48_;
  assign data_mem_data_o[816] = data_mem_data_o_7__48_;
  assign data_mem_data_o[944] = data_mem_data_o_7__48_;
  assign data_mem_data_o[47] = data_mem_data_o_7__47_;
  assign data_mem_data_o[175] = data_mem_data_o_7__47_;
  assign data_mem_data_o[303] = data_mem_data_o_7__47_;
  assign data_mem_data_o[431] = data_mem_data_o_7__47_;
  assign data_mem_data_o[559] = data_mem_data_o_7__47_;
  assign data_mem_data_o[687] = data_mem_data_o_7__47_;
  assign data_mem_data_o[815] = data_mem_data_o_7__47_;
  assign data_mem_data_o[943] = data_mem_data_o_7__47_;
  assign data_mem_data_o[46] = data_mem_data_o_7__46_;
  assign data_mem_data_o[174] = data_mem_data_o_7__46_;
  assign data_mem_data_o[302] = data_mem_data_o_7__46_;
  assign data_mem_data_o[430] = data_mem_data_o_7__46_;
  assign data_mem_data_o[558] = data_mem_data_o_7__46_;
  assign data_mem_data_o[686] = data_mem_data_o_7__46_;
  assign data_mem_data_o[814] = data_mem_data_o_7__46_;
  assign data_mem_data_o[942] = data_mem_data_o_7__46_;
  assign data_mem_data_o[45] = data_mem_data_o_7__45_;
  assign data_mem_data_o[173] = data_mem_data_o_7__45_;
  assign data_mem_data_o[301] = data_mem_data_o_7__45_;
  assign data_mem_data_o[429] = data_mem_data_o_7__45_;
  assign data_mem_data_o[557] = data_mem_data_o_7__45_;
  assign data_mem_data_o[685] = data_mem_data_o_7__45_;
  assign data_mem_data_o[813] = data_mem_data_o_7__45_;
  assign data_mem_data_o[941] = data_mem_data_o_7__45_;
  assign data_mem_data_o[44] = data_mem_data_o_7__44_;
  assign data_mem_data_o[172] = data_mem_data_o_7__44_;
  assign data_mem_data_o[300] = data_mem_data_o_7__44_;
  assign data_mem_data_o[428] = data_mem_data_o_7__44_;
  assign data_mem_data_o[556] = data_mem_data_o_7__44_;
  assign data_mem_data_o[684] = data_mem_data_o_7__44_;
  assign data_mem_data_o[812] = data_mem_data_o_7__44_;
  assign data_mem_data_o[940] = data_mem_data_o_7__44_;
  assign data_mem_data_o[43] = data_mem_data_o_7__43_;
  assign data_mem_data_o[171] = data_mem_data_o_7__43_;
  assign data_mem_data_o[299] = data_mem_data_o_7__43_;
  assign data_mem_data_o[427] = data_mem_data_o_7__43_;
  assign data_mem_data_o[555] = data_mem_data_o_7__43_;
  assign data_mem_data_o[683] = data_mem_data_o_7__43_;
  assign data_mem_data_o[811] = data_mem_data_o_7__43_;
  assign data_mem_data_o[939] = data_mem_data_o_7__43_;
  assign data_mem_data_o[42] = data_mem_data_o_7__42_;
  assign data_mem_data_o[170] = data_mem_data_o_7__42_;
  assign data_mem_data_o[298] = data_mem_data_o_7__42_;
  assign data_mem_data_o[426] = data_mem_data_o_7__42_;
  assign data_mem_data_o[554] = data_mem_data_o_7__42_;
  assign data_mem_data_o[682] = data_mem_data_o_7__42_;
  assign data_mem_data_o[810] = data_mem_data_o_7__42_;
  assign data_mem_data_o[938] = data_mem_data_o_7__42_;
  assign data_mem_data_o[41] = data_mem_data_o_7__41_;
  assign data_mem_data_o[169] = data_mem_data_o_7__41_;
  assign data_mem_data_o[297] = data_mem_data_o_7__41_;
  assign data_mem_data_o[425] = data_mem_data_o_7__41_;
  assign data_mem_data_o[553] = data_mem_data_o_7__41_;
  assign data_mem_data_o[681] = data_mem_data_o_7__41_;
  assign data_mem_data_o[809] = data_mem_data_o_7__41_;
  assign data_mem_data_o[937] = data_mem_data_o_7__41_;
  assign data_mem_data_o[40] = data_mem_data_o_7__40_;
  assign data_mem_data_o[168] = data_mem_data_o_7__40_;
  assign data_mem_data_o[296] = data_mem_data_o_7__40_;
  assign data_mem_data_o[424] = data_mem_data_o_7__40_;
  assign data_mem_data_o[552] = data_mem_data_o_7__40_;
  assign data_mem_data_o[680] = data_mem_data_o_7__40_;
  assign data_mem_data_o[808] = data_mem_data_o_7__40_;
  assign data_mem_data_o[936] = data_mem_data_o_7__40_;
  assign data_mem_data_o[39] = data_mem_data_o_7__39_;
  assign data_mem_data_o[167] = data_mem_data_o_7__39_;
  assign data_mem_data_o[295] = data_mem_data_o_7__39_;
  assign data_mem_data_o[423] = data_mem_data_o_7__39_;
  assign data_mem_data_o[551] = data_mem_data_o_7__39_;
  assign data_mem_data_o[679] = data_mem_data_o_7__39_;
  assign data_mem_data_o[807] = data_mem_data_o_7__39_;
  assign data_mem_data_o[935] = data_mem_data_o_7__39_;
  assign data_mem_data_o[38] = data_mem_data_o_7__38_;
  assign data_mem_data_o[166] = data_mem_data_o_7__38_;
  assign data_mem_data_o[294] = data_mem_data_o_7__38_;
  assign data_mem_data_o[422] = data_mem_data_o_7__38_;
  assign data_mem_data_o[550] = data_mem_data_o_7__38_;
  assign data_mem_data_o[678] = data_mem_data_o_7__38_;
  assign data_mem_data_o[806] = data_mem_data_o_7__38_;
  assign data_mem_data_o[934] = data_mem_data_o_7__38_;
  assign data_mem_data_o[37] = data_mem_data_o_7__37_;
  assign data_mem_data_o[165] = data_mem_data_o_7__37_;
  assign data_mem_data_o[293] = data_mem_data_o_7__37_;
  assign data_mem_data_o[421] = data_mem_data_o_7__37_;
  assign data_mem_data_o[549] = data_mem_data_o_7__37_;
  assign data_mem_data_o[677] = data_mem_data_o_7__37_;
  assign data_mem_data_o[805] = data_mem_data_o_7__37_;
  assign data_mem_data_o[933] = data_mem_data_o_7__37_;
  assign data_mem_data_o[36] = data_mem_data_o_7__36_;
  assign data_mem_data_o[164] = data_mem_data_o_7__36_;
  assign data_mem_data_o[292] = data_mem_data_o_7__36_;
  assign data_mem_data_o[420] = data_mem_data_o_7__36_;
  assign data_mem_data_o[548] = data_mem_data_o_7__36_;
  assign data_mem_data_o[676] = data_mem_data_o_7__36_;
  assign data_mem_data_o[804] = data_mem_data_o_7__36_;
  assign data_mem_data_o[932] = data_mem_data_o_7__36_;
  assign data_mem_data_o[35] = data_mem_data_o_7__35_;
  assign data_mem_data_o[163] = data_mem_data_o_7__35_;
  assign data_mem_data_o[291] = data_mem_data_o_7__35_;
  assign data_mem_data_o[419] = data_mem_data_o_7__35_;
  assign data_mem_data_o[547] = data_mem_data_o_7__35_;
  assign data_mem_data_o[675] = data_mem_data_o_7__35_;
  assign data_mem_data_o[803] = data_mem_data_o_7__35_;
  assign data_mem_data_o[931] = data_mem_data_o_7__35_;
  assign data_mem_data_o[34] = data_mem_data_o_7__34_;
  assign data_mem_data_o[162] = data_mem_data_o_7__34_;
  assign data_mem_data_o[290] = data_mem_data_o_7__34_;
  assign data_mem_data_o[418] = data_mem_data_o_7__34_;
  assign data_mem_data_o[546] = data_mem_data_o_7__34_;
  assign data_mem_data_o[674] = data_mem_data_o_7__34_;
  assign data_mem_data_o[802] = data_mem_data_o_7__34_;
  assign data_mem_data_o[930] = data_mem_data_o_7__34_;
  assign data_mem_data_o[33] = data_mem_data_o_7__33_;
  assign data_mem_data_o[161] = data_mem_data_o_7__33_;
  assign data_mem_data_o[289] = data_mem_data_o_7__33_;
  assign data_mem_data_o[417] = data_mem_data_o_7__33_;
  assign data_mem_data_o[545] = data_mem_data_o_7__33_;
  assign data_mem_data_o[673] = data_mem_data_o_7__33_;
  assign data_mem_data_o[801] = data_mem_data_o_7__33_;
  assign data_mem_data_o[929] = data_mem_data_o_7__33_;
  assign data_mem_data_o[32] = data_mem_data_o_7__32_;
  assign data_mem_data_o[160] = data_mem_data_o_7__32_;
  assign data_mem_data_o[288] = data_mem_data_o_7__32_;
  assign data_mem_data_o[416] = data_mem_data_o_7__32_;
  assign data_mem_data_o[544] = data_mem_data_o_7__32_;
  assign data_mem_data_o[672] = data_mem_data_o_7__32_;
  assign data_mem_data_o[800] = data_mem_data_o_7__32_;
  assign data_mem_data_o[928] = data_mem_data_o_7__32_;
  assign data_mem_data_o[31] = data_mem_data_o_7__31_;
  assign data_mem_data_o[159] = data_mem_data_o_7__31_;
  assign data_mem_data_o[287] = data_mem_data_o_7__31_;
  assign data_mem_data_o[415] = data_mem_data_o_7__31_;
  assign data_mem_data_o[543] = data_mem_data_o_7__31_;
  assign data_mem_data_o[671] = data_mem_data_o_7__31_;
  assign data_mem_data_o[799] = data_mem_data_o_7__31_;
  assign data_mem_data_o[927] = data_mem_data_o_7__31_;
  assign data_mem_data_o[30] = data_mem_data_o_7__30_;
  assign data_mem_data_o[158] = data_mem_data_o_7__30_;
  assign data_mem_data_o[286] = data_mem_data_o_7__30_;
  assign data_mem_data_o[414] = data_mem_data_o_7__30_;
  assign data_mem_data_o[542] = data_mem_data_o_7__30_;
  assign data_mem_data_o[670] = data_mem_data_o_7__30_;
  assign data_mem_data_o[798] = data_mem_data_o_7__30_;
  assign data_mem_data_o[926] = data_mem_data_o_7__30_;
  assign data_mem_data_o[29] = data_mem_data_o_7__29_;
  assign data_mem_data_o[157] = data_mem_data_o_7__29_;
  assign data_mem_data_o[285] = data_mem_data_o_7__29_;
  assign data_mem_data_o[413] = data_mem_data_o_7__29_;
  assign data_mem_data_o[541] = data_mem_data_o_7__29_;
  assign data_mem_data_o[669] = data_mem_data_o_7__29_;
  assign data_mem_data_o[797] = data_mem_data_o_7__29_;
  assign data_mem_data_o[925] = data_mem_data_o_7__29_;
  assign data_mem_data_o[28] = data_mem_data_o_7__28_;
  assign data_mem_data_o[156] = data_mem_data_o_7__28_;
  assign data_mem_data_o[284] = data_mem_data_o_7__28_;
  assign data_mem_data_o[412] = data_mem_data_o_7__28_;
  assign data_mem_data_o[540] = data_mem_data_o_7__28_;
  assign data_mem_data_o[668] = data_mem_data_o_7__28_;
  assign data_mem_data_o[796] = data_mem_data_o_7__28_;
  assign data_mem_data_o[924] = data_mem_data_o_7__28_;
  assign data_mem_data_o[27] = data_mem_data_o_7__27_;
  assign data_mem_data_o[155] = data_mem_data_o_7__27_;
  assign data_mem_data_o[283] = data_mem_data_o_7__27_;
  assign data_mem_data_o[411] = data_mem_data_o_7__27_;
  assign data_mem_data_o[539] = data_mem_data_o_7__27_;
  assign data_mem_data_o[667] = data_mem_data_o_7__27_;
  assign data_mem_data_o[795] = data_mem_data_o_7__27_;
  assign data_mem_data_o[923] = data_mem_data_o_7__27_;
  assign data_mem_data_o[26] = data_mem_data_o_7__26_;
  assign data_mem_data_o[154] = data_mem_data_o_7__26_;
  assign data_mem_data_o[282] = data_mem_data_o_7__26_;
  assign data_mem_data_o[410] = data_mem_data_o_7__26_;
  assign data_mem_data_o[538] = data_mem_data_o_7__26_;
  assign data_mem_data_o[666] = data_mem_data_o_7__26_;
  assign data_mem_data_o[794] = data_mem_data_o_7__26_;
  assign data_mem_data_o[922] = data_mem_data_o_7__26_;
  assign data_mem_data_o[25] = data_mem_data_o_7__25_;
  assign data_mem_data_o[153] = data_mem_data_o_7__25_;
  assign data_mem_data_o[281] = data_mem_data_o_7__25_;
  assign data_mem_data_o[409] = data_mem_data_o_7__25_;
  assign data_mem_data_o[537] = data_mem_data_o_7__25_;
  assign data_mem_data_o[665] = data_mem_data_o_7__25_;
  assign data_mem_data_o[793] = data_mem_data_o_7__25_;
  assign data_mem_data_o[921] = data_mem_data_o_7__25_;
  assign data_mem_data_o[24] = data_mem_data_o_7__24_;
  assign data_mem_data_o[152] = data_mem_data_o_7__24_;
  assign data_mem_data_o[280] = data_mem_data_o_7__24_;
  assign data_mem_data_o[408] = data_mem_data_o_7__24_;
  assign data_mem_data_o[536] = data_mem_data_o_7__24_;
  assign data_mem_data_o[664] = data_mem_data_o_7__24_;
  assign data_mem_data_o[792] = data_mem_data_o_7__24_;
  assign data_mem_data_o[920] = data_mem_data_o_7__24_;
  assign data_mem_data_o[23] = data_mem_data_o_7__23_;
  assign data_mem_data_o[151] = data_mem_data_o_7__23_;
  assign data_mem_data_o[279] = data_mem_data_o_7__23_;
  assign data_mem_data_o[407] = data_mem_data_o_7__23_;
  assign data_mem_data_o[535] = data_mem_data_o_7__23_;
  assign data_mem_data_o[663] = data_mem_data_o_7__23_;
  assign data_mem_data_o[791] = data_mem_data_o_7__23_;
  assign data_mem_data_o[919] = data_mem_data_o_7__23_;
  assign data_mem_data_o[22] = data_mem_data_o_7__22_;
  assign data_mem_data_o[150] = data_mem_data_o_7__22_;
  assign data_mem_data_o[278] = data_mem_data_o_7__22_;
  assign data_mem_data_o[406] = data_mem_data_o_7__22_;
  assign data_mem_data_o[534] = data_mem_data_o_7__22_;
  assign data_mem_data_o[662] = data_mem_data_o_7__22_;
  assign data_mem_data_o[790] = data_mem_data_o_7__22_;
  assign data_mem_data_o[918] = data_mem_data_o_7__22_;
  assign data_mem_data_o[21] = data_mem_data_o_7__21_;
  assign data_mem_data_o[149] = data_mem_data_o_7__21_;
  assign data_mem_data_o[277] = data_mem_data_o_7__21_;
  assign data_mem_data_o[405] = data_mem_data_o_7__21_;
  assign data_mem_data_o[533] = data_mem_data_o_7__21_;
  assign data_mem_data_o[661] = data_mem_data_o_7__21_;
  assign data_mem_data_o[789] = data_mem_data_o_7__21_;
  assign data_mem_data_o[917] = data_mem_data_o_7__21_;
  assign data_mem_data_o[20] = data_mem_data_o_7__20_;
  assign data_mem_data_o[148] = data_mem_data_o_7__20_;
  assign data_mem_data_o[276] = data_mem_data_o_7__20_;
  assign data_mem_data_o[404] = data_mem_data_o_7__20_;
  assign data_mem_data_o[532] = data_mem_data_o_7__20_;
  assign data_mem_data_o[660] = data_mem_data_o_7__20_;
  assign data_mem_data_o[788] = data_mem_data_o_7__20_;
  assign data_mem_data_o[916] = data_mem_data_o_7__20_;
  assign data_mem_data_o[19] = data_mem_data_o_7__19_;
  assign data_mem_data_o[147] = data_mem_data_o_7__19_;
  assign data_mem_data_o[275] = data_mem_data_o_7__19_;
  assign data_mem_data_o[403] = data_mem_data_o_7__19_;
  assign data_mem_data_o[531] = data_mem_data_o_7__19_;
  assign data_mem_data_o[659] = data_mem_data_o_7__19_;
  assign data_mem_data_o[787] = data_mem_data_o_7__19_;
  assign data_mem_data_o[915] = data_mem_data_o_7__19_;
  assign data_mem_data_o[18] = data_mem_data_o_7__18_;
  assign data_mem_data_o[146] = data_mem_data_o_7__18_;
  assign data_mem_data_o[274] = data_mem_data_o_7__18_;
  assign data_mem_data_o[402] = data_mem_data_o_7__18_;
  assign data_mem_data_o[530] = data_mem_data_o_7__18_;
  assign data_mem_data_o[658] = data_mem_data_o_7__18_;
  assign data_mem_data_o[786] = data_mem_data_o_7__18_;
  assign data_mem_data_o[914] = data_mem_data_o_7__18_;
  assign data_mem_data_o[17] = data_mem_data_o_7__17_;
  assign data_mem_data_o[145] = data_mem_data_o_7__17_;
  assign data_mem_data_o[273] = data_mem_data_o_7__17_;
  assign data_mem_data_o[401] = data_mem_data_o_7__17_;
  assign data_mem_data_o[529] = data_mem_data_o_7__17_;
  assign data_mem_data_o[657] = data_mem_data_o_7__17_;
  assign data_mem_data_o[785] = data_mem_data_o_7__17_;
  assign data_mem_data_o[913] = data_mem_data_o_7__17_;
  assign data_mem_data_o[16] = data_mem_data_o_7__16_;
  assign data_mem_data_o[144] = data_mem_data_o_7__16_;
  assign data_mem_data_o[272] = data_mem_data_o_7__16_;
  assign data_mem_data_o[400] = data_mem_data_o_7__16_;
  assign data_mem_data_o[528] = data_mem_data_o_7__16_;
  assign data_mem_data_o[656] = data_mem_data_o_7__16_;
  assign data_mem_data_o[784] = data_mem_data_o_7__16_;
  assign data_mem_data_o[912] = data_mem_data_o_7__16_;
  assign data_mem_data_o[15] = data_mem_data_o_7__15_;
  assign data_mem_data_o[143] = data_mem_data_o_7__15_;
  assign data_mem_data_o[271] = data_mem_data_o_7__15_;
  assign data_mem_data_o[399] = data_mem_data_o_7__15_;
  assign data_mem_data_o[527] = data_mem_data_o_7__15_;
  assign data_mem_data_o[655] = data_mem_data_o_7__15_;
  assign data_mem_data_o[783] = data_mem_data_o_7__15_;
  assign data_mem_data_o[911] = data_mem_data_o_7__15_;
  assign data_mem_data_o[14] = data_mem_data_o_7__14_;
  assign data_mem_data_o[142] = data_mem_data_o_7__14_;
  assign data_mem_data_o[270] = data_mem_data_o_7__14_;
  assign data_mem_data_o[398] = data_mem_data_o_7__14_;
  assign data_mem_data_o[526] = data_mem_data_o_7__14_;
  assign data_mem_data_o[654] = data_mem_data_o_7__14_;
  assign data_mem_data_o[782] = data_mem_data_o_7__14_;
  assign data_mem_data_o[910] = data_mem_data_o_7__14_;
  assign data_mem_data_o[13] = data_mem_data_o_7__13_;
  assign data_mem_data_o[141] = data_mem_data_o_7__13_;
  assign data_mem_data_o[269] = data_mem_data_o_7__13_;
  assign data_mem_data_o[397] = data_mem_data_o_7__13_;
  assign data_mem_data_o[525] = data_mem_data_o_7__13_;
  assign data_mem_data_o[653] = data_mem_data_o_7__13_;
  assign data_mem_data_o[781] = data_mem_data_o_7__13_;
  assign data_mem_data_o[909] = data_mem_data_o_7__13_;
  assign data_mem_data_o[12] = data_mem_data_o_7__12_;
  assign data_mem_data_o[140] = data_mem_data_o_7__12_;
  assign data_mem_data_o[268] = data_mem_data_o_7__12_;
  assign data_mem_data_o[396] = data_mem_data_o_7__12_;
  assign data_mem_data_o[524] = data_mem_data_o_7__12_;
  assign data_mem_data_o[652] = data_mem_data_o_7__12_;
  assign data_mem_data_o[780] = data_mem_data_o_7__12_;
  assign data_mem_data_o[908] = data_mem_data_o_7__12_;
  assign data_mem_data_o[11] = data_mem_data_o_7__11_;
  assign data_mem_data_o[139] = data_mem_data_o_7__11_;
  assign data_mem_data_o[267] = data_mem_data_o_7__11_;
  assign data_mem_data_o[395] = data_mem_data_o_7__11_;
  assign data_mem_data_o[523] = data_mem_data_o_7__11_;
  assign data_mem_data_o[651] = data_mem_data_o_7__11_;
  assign data_mem_data_o[779] = data_mem_data_o_7__11_;
  assign data_mem_data_o[907] = data_mem_data_o_7__11_;
  assign data_mem_data_o[10] = data_mem_data_o_7__10_;
  assign data_mem_data_o[138] = data_mem_data_o_7__10_;
  assign data_mem_data_o[266] = data_mem_data_o_7__10_;
  assign data_mem_data_o[394] = data_mem_data_o_7__10_;
  assign data_mem_data_o[522] = data_mem_data_o_7__10_;
  assign data_mem_data_o[650] = data_mem_data_o_7__10_;
  assign data_mem_data_o[778] = data_mem_data_o_7__10_;
  assign data_mem_data_o[906] = data_mem_data_o_7__10_;
  assign data_mem_data_o[9] = data_mem_data_o_7__9_;
  assign data_mem_data_o[137] = data_mem_data_o_7__9_;
  assign data_mem_data_o[265] = data_mem_data_o_7__9_;
  assign data_mem_data_o[393] = data_mem_data_o_7__9_;
  assign data_mem_data_o[521] = data_mem_data_o_7__9_;
  assign data_mem_data_o[649] = data_mem_data_o_7__9_;
  assign data_mem_data_o[777] = data_mem_data_o_7__9_;
  assign data_mem_data_o[905] = data_mem_data_o_7__9_;
  assign data_mem_data_o[8] = data_mem_data_o_7__8_;
  assign data_mem_data_o[136] = data_mem_data_o_7__8_;
  assign data_mem_data_o[264] = data_mem_data_o_7__8_;
  assign data_mem_data_o[392] = data_mem_data_o_7__8_;
  assign data_mem_data_o[520] = data_mem_data_o_7__8_;
  assign data_mem_data_o[648] = data_mem_data_o_7__8_;
  assign data_mem_data_o[776] = data_mem_data_o_7__8_;
  assign data_mem_data_o[904] = data_mem_data_o_7__8_;
  assign data_mem_data_o[7] = data_mem_data_o_7__7_;
  assign data_mem_data_o[135] = data_mem_data_o_7__7_;
  assign data_mem_data_o[263] = data_mem_data_o_7__7_;
  assign data_mem_data_o[391] = data_mem_data_o_7__7_;
  assign data_mem_data_o[519] = data_mem_data_o_7__7_;
  assign data_mem_data_o[647] = data_mem_data_o_7__7_;
  assign data_mem_data_o[775] = data_mem_data_o_7__7_;
  assign data_mem_data_o[903] = data_mem_data_o_7__7_;
  assign data_mem_data_o[6] = data_mem_data_o_7__6_;
  assign data_mem_data_o[134] = data_mem_data_o_7__6_;
  assign data_mem_data_o[262] = data_mem_data_o_7__6_;
  assign data_mem_data_o[390] = data_mem_data_o_7__6_;
  assign data_mem_data_o[518] = data_mem_data_o_7__6_;
  assign data_mem_data_o[646] = data_mem_data_o_7__6_;
  assign data_mem_data_o[774] = data_mem_data_o_7__6_;
  assign data_mem_data_o[902] = data_mem_data_o_7__6_;
  assign data_mem_data_o[5] = data_mem_data_o_7__5_;
  assign data_mem_data_o[133] = data_mem_data_o_7__5_;
  assign data_mem_data_o[261] = data_mem_data_o_7__5_;
  assign data_mem_data_o[389] = data_mem_data_o_7__5_;
  assign data_mem_data_o[517] = data_mem_data_o_7__5_;
  assign data_mem_data_o[645] = data_mem_data_o_7__5_;
  assign data_mem_data_o[773] = data_mem_data_o_7__5_;
  assign data_mem_data_o[901] = data_mem_data_o_7__5_;
  assign data_mem_data_o[4] = data_mem_data_o_7__4_;
  assign data_mem_data_o[132] = data_mem_data_o_7__4_;
  assign data_mem_data_o[260] = data_mem_data_o_7__4_;
  assign data_mem_data_o[388] = data_mem_data_o_7__4_;
  assign data_mem_data_o[516] = data_mem_data_o_7__4_;
  assign data_mem_data_o[644] = data_mem_data_o_7__4_;
  assign data_mem_data_o[772] = data_mem_data_o_7__4_;
  assign data_mem_data_o[900] = data_mem_data_o_7__4_;
  assign data_mem_data_o[3] = data_mem_data_o_7__3_;
  assign data_mem_data_o[131] = data_mem_data_o_7__3_;
  assign data_mem_data_o[259] = data_mem_data_o_7__3_;
  assign data_mem_data_o[387] = data_mem_data_o_7__3_;
  assign data_mem_data_o[515] = data_mem_data_o_7__3_;
  assign data_mem_data_o[643] = data_mem_data_o_7__3_;
  assign data_mem_data_o[771] = data_mem_data_o_7__3_;
  assign data_mem_data_o[899] = data_mem_data_o_7__3_;
  assign data_mem_data_o[2] = data_mem_data_o_7__2_;
  assign data_mem_data_o[130] = data_mem_data_o_7__2_;
  assign data_mem_data_o[258] = data_mem_data_o_7__2_;
  assign data_mem_data_o[386] = data_mem_data_o_7__2_;
  assign data_mem_data_o[514] = data_mem_data_o_7__2_;
  assign data_mem_data_o[642] = data_mem_data_o_7__2_;
  assign data_mem_data_o[770] = data_mem_data_o_7__2_;
  assign data_mem_data_o[898] = data_mem_data_o_7__2_;
  assign data_mem_data_o[1] = data_mem_data_o_7__1_;
  assign data_mem_data_o[129] = data_mem_data_o_7__1_;
  assign data_mem_data_o[257] = data_mem_data_o_7__1_;
  assign data_mem_data_o[385] = data_mem_data_o_7__1_;
  assign data_mem_data_o[513] = data_mem_data_o_7__1_;
  assign data_mem_data_o[641] = data_mem_data_o_7__1_;
  assign data_mem_data_o[769] = data_mem_data_o_7__1_;
  assign data_mem_data_o[897] = data_mem_data_o_7__1_;
  assign data_mem_data_o[0] = data_mem_data_o_7__0_;
  assign data_mem_data_o[128] = data_mem_data_o_7__0_;
  assign data_mem_data_o[256] = data_mem_data_o_7__0_;
  assign data_mem_data_o[384] = data_mem_data_o_7__0_;
  assign data_mem_data_o[512] = data_mem_data_o_7__0_;
  assign data_mem_data_o[640] = data_mem_data_o_7__0_;
  assign data_mem_data_o[768] = data_mem_data_o_7__0_;
  assign data_mem_data_o[896] = data_mem_data_o_7__0_;

  bsg_counter_clear_up_00000004_0
  dma_counter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(counter_clear),
    .up_i(counter_up),
    .count_o({ counter_r[2:2], data_mem_addr_o[1:0] })
  );


  bsg_fifo_1r1w_small_00000080_00000004
  in_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(dma_data_v_i),
    .ready_param_o(dma_data_ready_and_o),
    .data_i(dma_data_i),
    .v_o(in_fifo_v_lo),
    .data_o({ data_mem_data_o_7__127_, data_mem_data_o_7__126_, data_mem_data_o_7__125_, data_mem_data_o_7__124_, data_mem_data_o_7__123_, data_mem_data_o_7__122_, data_mem_data_o_7__121_, data_mem_data_o_7__120_, data_mem_data_o_7__119_, data_mem_data_o_7__118_, data_mem_data_o_7__117_, data_mem_data_o_7__116_, data_mem_data_o_7__115_, data_mem_data_o_7__114_, data_mem_data_o_7__113_, data_mem_data_o_7__112_, data_mem_data_o_7__111_, data_mem_data_o_7__110_, data_mem_data_o_7__109_, data_mem_data_o_7__108_, data_mem_data_o_7__107_, data_mem_data_o_7__106_, data_mem_data_o_7__105_, data_mem_data_o_7__104_, data_mem_data_o_7__103_, data_mem_data_o_7__102_, data_mem_data_o_7__101_, data_mem_data_o_7__100_, data_mem_data_o_7__99_, data_mem_data_o_7__98_, data_mem_data_o_7__97_, data_mem_data_o_7__96_, data_mem_data_o_7__95_, data_mem_data_o_7__94_, data_mem_data_o_7__93_, data_mem_data_o_7__92_, data_mem_data_o_7__91_, data_mem_data_o_7__90_, data_mem_data_o_7__89_, data_mem_data_o_7__88_, data_mem_data_o_7__87_, data_mem_data_o_7__86_, data_mem_data_o_7__85_, data_mem_data_o_7__84_, data_mem_data_o_7__83_, data_mem_data_o_7__82_, data_mem_data_o_7__81_, data_mem_data_o_7__80_, data_mem_data_o_7__79_, data_mem_data_o_7__78_, data_mem_data_o_7__77_, data_mem_data_o_7__76_, data_mem_data_o_7__75_, data_mem_data_o_7__74_, data_mem_data_o_7__73_, data_mem_data_o_7__72_, data_mem_data_o_7__71_, data_mem_data_o_7__70_, data_mem_data_o_7__69_, data_mem_data_o_7__68_, data_mem_data_o_7__67_, data_mem_data_o_7__66_, data_mem_data_o_7__65_, data_mem_data_o_7__64_, data_mem_data_o_7__63_, data_mem_data_o_7__62_, data_mem_data_o_7__61_, data_mem_data_o_7__60_, data_mem_data_o_7__59_, data_mem_data_o_7__58_, data_mem_data_o_7__57_, data_mem_data_o_7__56_, data_mem_data_o_7__55_, data_mem_data_o_7__54_, data_mem_data_o_7__53_, data_mem_data_o_7__52_, data_mem_data_o_7__51_, data_mem_data_o_7__50_, data_mem_data_o_7__49_, data_mem_data_o_7__48_, data_mem_data_o_7__47_, data_mem_data_o_7__46_, data_mem_data_o_7__45_, data_mem_data_o_7__44_, data_mem_data_o_7__43_, data_mem_data_o_7__42_, data_mem_data_o_7__41_, data_mem_data_o_7__40_, data_mem_data_o_7__39_, data_mem_data_o_7__38_, data_mem_data_o_7__37_, data_mem_data_o_7__36_, data_mem_data_o_7__35_, data_mem_data_o_7__34_, data_mem_data_o_7__33_, data_mem_data_o_7__32_, data_mem_data_o_7__31_, data_mem_data_o_7__30_, data_mem_data_o_7__29_, data_mem_data_o_7__28_, data_mem_data_o_7__27_, data_mem_data_o_7__26_, data_mem_data_o_7__25_, data_mem_data_o_7__24_, data_mem_data_o_7__23_, data_mem_data_o_7__22_, data_mem_data_o_7__21_, data_mem_data_o_7__20_, data_mem_data_o_7__19_, data_mem_data_o_7__18_, data_mem_data_o_7__17_, data_mem_data_o_7__16_, data_mem_data_o_7__15_, data_mem_data_o_7__14_, data_mem_data_o_7__13_, data_mem_data_o_7__12_, data_mem_data_o_7__11_, data_mem_data_o_7__10_, data_mem_data_o_7__9_, data_mem_data_o_7__8_, data_mem_data_o_7__7_, data_mem_data_o_7__6_, data_mem_data_o_7__5_, data_mem_data_o_7__4_, data_mem_data_o_7__3_, data_mem_data_o_7__2_, data_mem_data_o_7__1_, data_mem_data_o_7__0_ }),
    .yumi_i(in_fifo_yumi_li)
  );


  bsg_two_fifo_00000080
  out_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_param_o(out_fifo_ready_lo),
    .data_i(out_fifo_data_li),
    .v_i(out_fifo_v_li),
    .v_o(dma_data_v_o),
    .data_o(dma_data_o),
    .yumi_i(dma_data_yumi_i)
  );


  bsg_decode_00000008
  dma_way_demux
  (
    .i(dma_way_i),
    .o(dma_way_mask)
  );


  bsg_expand_bitmask_00000008_00000010
  expand0
  (
    .i(dma_way_mask),
    .o(dma_way_mask_expanded)
  );


  bsg_mux_00000004_00000008
  track_way_mux
  (
    .data_i(track_mem_data_r),
    .sel_i(dma_way_i),
    .data_o(track_data_way_picked)
  );


  bsg_mux_00000001_00000004
  track_offset_mux
  (
    .data_i(track_data_way_picked),
    .sel_i(data_mem_addr_o[1:0]),
    .data_o(track_bits_offset_picked[0])
  );


  bsg_expand_bitmask_00000001_00000010
  expand1
  (
    .i(track_bits_offset_picked[0]),
    .o(track_bits_offset_picked_expanded)
  );


  bsg_mux_00000080_00000008
  write_data_mux
  (
    .data_i(data_mem_data_i),
    .sel_i(dma_way_i),
    .data_o(out_fifo_data_li)
  );

  assign N30 = N29 & N98;
  assign N31 = dma_state_r[1] | N98;
  assign N33 = N29 | dma_state_r[0];
  assign N35 = dma_state_r[1] & dma_state_r[0];
  assign N36 = dma_cmd_i[1] | N53;
  assign N37 = N39 | N36;
  assign N39 = dma_cmd_i[3] | dma_cmd_i[2];
  assign N40 = N52 | dma_cmd_i[0];
  assign N41 = N39 | N40;
  assign N43 = dma_cmd_i[3] | N51;
  assign N44 = N43 | N47;
  assign N46 = N50 | dma_cmd_i[2];
  assign N47 = dma_cmd_i[1] | dma_cmd_i[0];
  assign N48 = N46 | N47;
  assign N54 = N50 & N51;
  assign N55 = N52 & N53;
  assign N56 = N54 & N55;
  assign N83 = data_mem_addr_o[1:0] == dma_addr_i[5:4];

  bsg_mux_00000080_00000001
  snoop_mux0
  (
    .data_i({ data_mem_data_o_7__127_, data_mem_data_o_7__126_, data_mem_data_o_7__125_, data_mem_data_o_7__124_, data_mem_data_o_7__123_, data_mem_data_o_7__122_, data_mem_data_o_7__121_, data_mem_data_o_7__120_, data_mem_data_o_7__119_, data_mem_data_o_7__118_, data_mem_data_o_7__117_, data_mem_data_o_7__116_, data_mem_data_o_7__115_, data_mem_data_o_7__114_, data_mem_data_o_7__113_, data_mem_data_o_7__112_, data_mem_data_o_7__111_, data_mem_data_o_7__110_, data_mem_data_o_7__109_, data_mem_data_o_7__108_, data_mem_data_o_7__107_, data_mem_data_o_7__106_, data_mem_data_o_7__105_, data_mem_data_o_7__104_, data_mem_data_o_7__103_, data_mem_data_o_7__102_, data_mem_data_o_7__101_, data_mem_data_o_7__100_, data_mem_data_o_7__99_, data_mem_data_o_7__98_, data_mem_data_o_7__97_, data_mem_data_o_7__96_, data_mem_data_o_7__95_, data_mem_data_o_7__94_, data_mem_data_o_7__93_, data_mem_data_o_7__92_, data_mem_data_o_7__91_, data_mem_data_o_7__90_, data_mem_data_o_7__89_, data_mem_data_o_7__88_, data_mem_data_o_7__87_, data_mem_data_o_7__86_, data_mem_data_o_7__85_, data_mem_data_o_7__84_, data_mem_data_o_7__83_, data_mem_data_o_7__82_, data_mem_data_o_7__81_, data_mem_data_o_7__80_, data_mem_data_o_7__79_, data_mem_data_o_7__78_, data_mem_data_o_7__77_, data_mem_data_o_7__76_, data_mem_data_o_7__75_, data_mem_data_o_7__74_, data_mem_data_o_7__73_, data_mem_data_o_7__72_, data_mem_data_o_7__71_, data_mem_data_o_7__70_, data_mem_data_o_7__69_, data_mem_data_o_7__68_, data_mem_data_o_7__67_, data_mem_data_o_7__66_, data_mem_data_o_7__65_, data_mem_data_o_7__64_, data_mem_data_o_7__63_, data_mem_data_o_7__62_, data_mem_data_o_7__61_, data_mem_data_o_7__60_, data_mem_data_o_7__59_, data_mem_data_o_7__58_, data_mem_data_o_7__57_, data_mem_data_o_7__56_, data_mem_data_o_7__55_, data_mem_data_o_7__54_, data_mem_data_o_7__53_, data_mem_data_o_7__52_, data_mem_data_o_7__51_, data_mem_data_o_7__50_, data_mem_data_o_7__49_, data_mem_data_o_7__48_, data_mem_data_o_7__47_, data_mem_data_o_7__46_, data_mem_data_o_7__45_, data_mem_data_o_7__44_, data_mem_data_o_7__43_, data_mem_data_o_7__42_, data_mem_data_o_7__41_, data_mem_data_o_7__40_, data_mem_data_o_7__39_, data_mem_data_o_7__38_, data_mem_data_o_7__37_, data_mem_data_o_7__36_, data_mem_data_o_7__35_, data_mem_data_o_7__34_, data_mem_data_o_7__33_, data_mem_data_o_7__32_, data_mem_data_o_7__31_, data_mem_data_o_7__30_, data_mem_data_o_7__29_, data_mem_data_o_7__28_, data_mem_data_o_7__27_, data_mem_data_o_7__26_, data_mem_data_o_7__25_, data_mem_data_o_7__24_, data_mem_data_o_7__23_, data_mem_data_o_7__22_, data_mem_data_o_7__21_, data_mem_data_o_7__20_, data_mem_data_o_7__19_, data_mem_data_o_7__18_, data_mem_data_o_7__17_, data_mem_data_o_7__16_, data_mem_data_o_7__15_, data_mem_data_o_7__14_, data_mem_data_o_7__13_, data_mem_data_o_7__12_, data_mem_data_o_7__11_, data_mem_data_o_7__10_, data_mem_data_o_7__9_, data_mem_data_o_7__8_, data_mem_data_o_7__7_, data_mem_data_o_7__6_, data_mem_data_o_7__5_, data_mem_data_o_7__4_, data_mem_data_o_7__3_, data_mem_data_o_7__2_, data_mem_data_o_7__1_, data_mem_data_o_7__0_ }),
    .sel_i(dma_addr_i[4]),
    .data_o(snoop_word_n)
  );

  assign N89 = ~counter_r[2];
  assign N90 = data_mem_addr_o[1] | N89;
  assign N91 = data_mem_addr_o[0] | N90;
  assign N92 = ~N91;
  assign N93 = ~data_mem_addr_o[1];
  assign N94 = ~data_mem_addr_o[0];
  assign N95 = N93 | counter_r[2];
  assign N96 = N94 | N95;
  assign N97 = ~N96;
  assign N98 = ~dma_state_r[0];
  assign N99 = N98 | dma_state_r[1];
  assign N100 = ~N99;
  assign data_mem_w_mask_way_picked = (N0)? { N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28 } : 
                                      (N12)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N0 = track_miss_i;
  assign N62 = (N1)? 1'b1 : 
               (N2)? 1'b1 : 
               (N3)? 1'b0 : 
               (N4)? 1'b0 : 
               (N5)? 1'b0 : 
               (N61)? 1'b0 : 1'b0;
  assign N1 = N38;
  assign N2 = N42;
  assign N3 = N45;
  assign N4 = N49;
  assign N5 = N56;
  assign { N67, N66, N65, N64, N63 } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                       (N2)? { 1'b1, track_data_way_picked } : 
                                       (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                       (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                       (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                       (N61)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N68 = (N1)? dma_pkt_yumi_i : 
               (N2)? dma_pkt_yumi_i : 
               (N3)? 1'b0 : 
               (N4)? 1'b0 : 
               (N5)? 1'b0 : 
               (N61)? 1'b0 : 1'b0;
  assign N69 = (N1)? 1'b0 : 
               (N2)? 1'b0 : 
               (N3)? 1'b1 : 
               (N4)? 1'b1 : 
               (N5)? 1'b0 : 
               (N61)? 1'b0 : 1'b0;
  assign N70 = (N1)? 1'b0 : 
               (N2)? 1'b0 : 
               (N3)? 1'b0 : 
               (N4)? 1'b1 : 
               (N5)? 1'b0 : 
               (N61)? 1'b0 : 1'b0;
  assign N71 = (N1)? 1'b0 : 
               (N2)? 1'b0 : 
               (N3)? 1'b0 : 
               (N4)? track_bits_offset_picked[0] : 
               (N5)? 1'b0 : 
               (N61)? 1'b0 : 1'b0;
  assign N73 = ~N72;
  assign N78 = ~N77;
  assign counter_clear = (N6)? N69 : 
                         (N7)? N75 : 
                         (N8)? N80 : 
                         (N9)? 1'b0 : 1'b0;
  assign N6 = N30;
  assign N7 = N32;
  assign N8 = N34;
  assign N9 = N35;
  assign counter_up = (N6)? N70 : 
                      (N7)? N74 : 
                      (N8)? N79 : 
                      (N9)? 1'b0 : 1'b0;
  assign data_mem_v_o = (N6)? N71 : 
                        (N7)? in_fifo_v_lo : 
                        (N8)? N81 : 
                        (N9)? 1'b0 : 1'b0;
  assign dma_pkt_v_o = (N6)? N62 : 
                       (N7)? 1'b0 : 
                       (N8)? 1'b0 : 
                       (N9)? 1'b0 : 1'b0;
  assign { dma_pkt_o[37:37], dma_pkt_o[3:0] } = (N6)? { N67, N66, N65, N64, N63 } : 
                                                (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign done_o = (N6)? N68 : 
                  (N7)? N76 : 
                  (N8)? N82 : 
                  (N9)? 1'b0 : 1'b0;
  assign dma_state_n = (N6)? { N49, N45 } : 
                       (N7)? { 1'b0, N73 } : 
                       (N8)? { N78, 1'b0 } : 
                       (N9)? { 1'b0, 1'b0 } : 1'b0;
  assign data_mem_w_o = (N6)? 1'b0 : 
                        (N7)? in_fifo_v_lo : 
                        (N8)? 1'b0 : 
                        (N9)? 1'b0 : 1'b0;
  assign in_fifo_yumi_li = (N6)? 1'b0 : 
                           (N7)? in_fifo_v_lo : 
                           (N8)? 1'b0 : 
                           (N9)? 1'b0 : 1'b0;
  assign out_fifo_v_li = (N6)? 1'b0 : 
                         (N7)? 1'b0 : 
                         (N8)? 1'b1 : 
                         (N9)? 1'b0 : 1'b0;
  assign dma_evict_o = (N6)? 1'b0 : 
                       (N7)? 1'b0 : 
                       (N8)? 1'b1 : 
                       (N9)? 1'b0 : 1'b0;
  assign { N87, N86 } = (N10)? { 1'b0, 1'b0 } : 
                        (N11)? { snoop_word_we, snoop_word_we } : 1'b0;
  assign N10 = N85;
  assign N11 = N84;
  assign N88 = (N10)? 1'b0 : 
               (N11)? track_data_we_i : 1'b0;
  assign N12 = ~track_miss_i;
  assign N13 = ~track_bits_offset_picked_expanded[15];
  assign N14 = ~track_bits_offset_picked_expanded[14];
  assign N15 = ~track_bits_offset_picked_expanded[13];
  assign N16 = ~track_bits_offset_picked_expanded[12];
  assign N17 = ~track_bits_offset_picked_expanded[11];
  assign N18 = ~track_bits_offset_picked_expanded[10];
  assign N19 = ~track_bits_offset_picked_expanded[9];
  assign N20 = ~track_bits_offset_picked_expanded[8];
  assign N21 = ~track_bits_offset_picked_expanded[7];
  assign N22 = ~track_bits_offset_picked_expanded[6];
  assign N23 = ~track_bits_offset_picked_expanded[5];
  assign N24 = ~track_bits_offset_picked_expanded[4];
  assign N25 = ~track_bits_offset_picked_expanded[3];
  assign N26 = ~track_bits_offset_picked_expanded[2];
  assign N27 = ~track_bits_offset_picked_expanded[1];
  assign N28 = ~track_bits_offset_picked_expanded[0];
  assign data_mem_w_mask_o[127] = dma_way_mask_expanded[127] & data_mem_w_mask_way_picked[15];
  assign data_mem_w_mask_o[126] = dma_way_mask_expanded[126] & data_mem_w_mask_way_picked[14];
  assign data_mem_w_mask_o[125] = dma_way_mask_expanded[125] & data_mem_w_mask_way_picked[13];
  assign data_mem_w_mask_o[124] = dma_way_mask_expanded[124] & data_mem_w_mask_way_picked[12];
  assign data_mem_w_mask_o[123] = dma_way_mask_expanded[123] & data_mem_w_mask_way_picked[11];
  assign data_mem_w_mask_o[122] = dma_way_mask_expanded[122] & data_mem_w_mask_way_picked[10];
  assign data_mem_w_mask_o[121] = dma_way_mask_expanded[121] & data_mem_w_mask_way_picked[9];
  assign data_mem_w_mask_o[120] = dma_way_mask_expanded[120] & data_mem_w_mask_way_picked[8];
  assign data_mem_w_mask_o[119] = dma_way_mask_expanded[119] & data_mem_w_mask_way_picked[7];
  assign data_mem_w_mask_o[118] = dma_way_mask_expanded[118] & data_mem_w_mask_way_picked[6];
  assign data_mem_w_mask_o[117] = dma_way_mask_expanded[117] & data_mem_w_mask_way_picked[5];
  assign data_mem_w_mask_o[116] = dma_way_mask_expanded[116] & data_mem_w_mask_way_picked[4];
  assign data_mem_w_mask_o[115] = dma_way_mask_expanded[115] & data_mem_w_mask_way_picked[3];
  assign data_mem_w_mask_o[114] = dma_way_mask_expanded[114] & data_mem_w_mask_way_picked[2];
  assign data_mem_w_mask_o[113] = dma_way_mask_expanded[113] & data_mem_w_mask_way_picked[1];
  assign data_mem_w_mask_o[112] = dma_way_mask_expanded[112] & data_mem_w_mask_way_picked[0];
  assign data_mem_w_mask_o[111] = dma_way_mask_expanded[111] & data_mem_w_mask_way_picked[15];
  assign data_mem_w_mask_o[110] = dma_way_mask_expanded[110] & data_mem_w_mask_way_picked[14];
  assign data_mem_w_mask_o[109] = dma_way_mask_expanded[109] & data_mem_w_mask_way_picked[13];
  assign data_mem_w_mask_o[108] = dma_way_mask_expanded[108] & data_mem_w_mask_way_picked[12];
  assign data_mem_w_mask_o[107] = dma_way_mask_expanded[107] & data_mem_w_mask_way_picked[11];
  assign data_mem_w_mask_o[106] = dma_way_mask_expanded[106] & data_mem_w_mask_way_picked[10];
  assign data_mem_w_mask_o[105] = dma_way_mask_expanded[105] & data_mem_w_mask_way_picked[9];
  assign data_mem_w_mask_o[104] = dma_way_mask_expanded[104] & data_mem_w_mask_way_picked[8];
  assign data_mem_w_mask_o[103] = dma_way_mask_expanded[103] & data_mem_w_mask_way_picked[7];
  assign data_mem_w_mask_o[102] = dma_way_mask_expanded[102] & data_mem_w_mask_way_picked[6];
  assign data_mem_w_mask_o[101] = dma_way_mask_expanded[101] & data_mem_w_mask_way_picked[5];
  assign data_mem_w_mask_o[100] = dma_way_mask_expanded[100] & data_mem_w_mask_way_picked[4];
  assign data_mem_w_mask_o[99] = dma_way_mask_expanded[99] & data_mem_w_mask_way_picked[3];
  assign data_mem_w_mask_o[98] = dma_way_mask_expanded[98] & data_mem_w_mask_way_picked[2];
  assign data_mem_w_mask_o[97] = dma_way_mask_expanded[97] & data_mem_w_mask_way_picked[1];
  assign data_mem_w_mask_o[96] = dma_way_mask_expanded[96] & data_mem_w_mask_way_picked[0];
  assign data_mem_w_mask_o[95] = dma_way_mask_expanded[95] & data_mem_w_mask_way_picked[15];
  assign data_mem_w_mask_o[94] = dma_way_mask_expanded[94] & data_mem_w_mask_way_picked[14];
  assign data_mem_w_mask_o[93] = dma_way_mask_expanded[93] & data_mem_w_mask_way_picked[13];
  assign data_mem_w_mask_o[92] = dma_way_mask_expanded[92] & data_mem_w_mask_way_picked[12];
  assign data_mem_w_mask_o[91] = dma_way_mask_expanded[91] & data_mem_w_mask_way_picked[11];
  assign data_mem_w_mask_o[90] = dma_way_mask_expanded[90] & data_mem_w_mask_way_picked[10];
  assign data_mem_w_mask_o[89] = dma_way_mask_expanded[89] & data_mem_w_mask_way_picked[9];
  assign data_mem_w_mask_o[88] = dma_way_mask_expanded[88] & data_mem_w_mask_way_picked[8];
  assign data_mem_w_mask_o[87] = dma_way_mask_expanded[87] & data_mem_w_mask_way_picked[7];
  assign data_mem_w_mask_o[86] = dma_way_mask_expanded[86] & data_mem_w_mask_way_picked[6];
  assign data_mem_w_mask_o[85] = dma_way_mask_expanded[85] & data_mem_w_mask_way_picked[5];
  assign data_mem_w_mask_o[84] = dma_way_mask_expanded[84] & data_mem_w_mask_way_picked[4];
  assign data_mem_w_mask_o[83] = dma_way_mask_expanded[83] & data_mem_w_mask_way_picked[3];
  assign data_mem_w_mask_o[82] = dma_way_mask_expanded[82] & data_mem_w_mask_way_picked[2];
  assign data_mem_w_mask_o[81] = dma_way_mask_expanded[81] & data_mem_w_mask_way_picked[1];
  assign data_mem_w_mask_o[80] = dma_way_mask_expanded[80] & data_mem_w_mask_way_picked[0];
  assign data_mem_w_mask_o[79] = dma_way_mask_expanded[79] & data_mem_w_mask_way_picked[15];
  assign data_mem_w_mask_o[78] = dma_way_mask_expanded[78] & data_mem_w_mask_way_picked[14];
  assign data_mem_w_mask_o[77] = dma_way_mask_expanded[77] & data_mem_w_mask_way_picked[13];
  assign data_mem_w_mask_o[76] = dma_way_mask_expanded[76] & data_mem_w_mask_way_picked[12];
  assign data_mem_w_mask_o[75] = dma_way_mask_expanded[75] & data_mem_w_mask_way_picked[11];
  assign data_mem_w_mask_o[74] = dma_way_mask_expanded[74] & data_mem_w_mask_way_picked[10];
  assign data_mem_w_mask_o[73] = dma_way_mask_expanded[73] & data_mem_w_mask_way_picked[9];
  assign data_mem_w_mask_o[72] = dma_way_mask_expanded[72] & data_mem_w_mask_way_picked[8];
  assign data_mem_w_mask_o[71] = dma_way_mask_expanded[71] & data_mem_w_mask_way_picked[7];
  assign data_mem_w_mask_o[70] = dma_way_mask_expanded[70] & data_mem_w_mask_way_picked[6];
  assign data_mem_w_mask_o[69] = dma_way_mask_expanded[69] & data_mem_w_mask_way_picked[5];
  assign data_mem_w_mask_o[68] = dma_way_mask_expanded[68] & data_mem_w_mask_way_picked[4];
  assign data_mem_w_mask_o[67] = dma_way_mask_expanded[67] & data_mem_w_mask_way_picked[3];
  assign data_mem_w_mask_o[66] = dma_way_mask_expanded[66] & data_mem_w_mask_way_picked[2];
  assign data_mem_w_mask_o[65] = dma_way_mask_expanded[65] & data_mem_w_mask_way_picked[1];
  assign data_mem_w_mask_o[64] = dma_way_mask_expanded[64] & data_mem_w_mask_way_picked[0];
  assign data_mem_w_mask_o[63] = dma_way_mask_expanded[63] & data_mem_w_mask_way_picked[15];
  assign data_mem_w_mask_o[62] = dma_way_mask_expanded[62] & data_mem_w_mask_way_picked[14];
  assign data_mem_w_mask_o[61] = dma_way_mask_expanded[61] & data_mem_w_mask_way_picked[13];
  assign data_mem_w_mask_o[60] = dma_way_mask_expanded[60] & data_mem_w_mask_way_picked[12];
  assign data_mem_w_mask_o[59] = dma_way_mask_expanded[59] & data_mem_w_mask_way_picked[11];
  assign data_mem_w_mask_o[58] = dma_way_mask_expanded[58] & data_mem_w_mask_way_picked[10];
  assign data_mem_w_mask_o[57] = dma_way_mask_expanded[57] & data_mem_w_mask_way_picked[9];
  assign data_mem_w_mask_o[56] = dma_way_mask_expanded[56] & data_mem_w_mask_way_picked[8];
  assign data_mem_w_mask_o[55] = dma_way_mask_expanded[55] & data_mem_w_mask_way_picked[7];
  assign data_mem_w_mask_o[54] = dma_way_mask_expanded[54] & data_mem_w_mask_way_picked[6];
  assign data_mem_w_mask_o[53] = dma_way_mask_expanded[53] & data_mem_w_mask_way_picked[5];
  assign data_mem_w_mask_o[52] = dma_way_mask_expanded[52] & data_mem_w_mask_way_picked[4];
  assign data_mem_w_mask_o[51] = dma_way_mask_expanded[51] & data_mem_w_mask_way_picked[3];
  assign data_mem_w_mask_o[50] = dma_way_mask_expanded[50] & data_mem_w_mask_way_picked[2];
  assign data_mem_w_mask_o[49] = dma_way_mask_expanded[49] & data_mem_w_mask_way_picked[1];
  assign data_mem_w_mask_o[48] = dma_way_mask_expanded[48] & data_mem_w_mask_way_picked[0];
  assign data_mem_w_mask_o[47] = dma_way_mask_expanded[47] & data_mem_w_mask_way_picked[15];
  assign data_mem_w_mask_o[46] = dma_way_mask_expanded[46] & data_mem_w_mask_way_picked[14];
  assign data_mem_w_mask_o[45] = dma_way_mask_expanded[45] & data_mem_w_mask_way_picked[13];
  assign data_mem_w_mask_o[44] = dma_way_mask_expanded[44] & data_mem_w_mask_way_picked[12];
  assign data_mem_w_mask_o[43] = dma_way_mask_expanded[43] & data_mem_w_mask_way_picked[11];
  assign data_mem_w_mask_o[42] = dma_way_mask_expanded[42] & data_mem_w_mask_way_picked[10];
  assign data_mem_w_mask_o[41] = dma_way_mask_expanded[41] & data_mem_w_mask_way_picked[9];
  assign data_mem_w_mask_o[40] = dma_way_mask_expanded[40] & data_mem_w_mask_way_picked[8];
  assign data_mem_w_mask_o[39] = dma_way_mask_expanded[39] & data_mem_w_mask_way_picked[7];
  assign data_mem_w_mask_o[38] = dma_way_mask_expanded[38] & data_mem_w_mask_way_picked[6];
  assign data_mem_w_mask_o[37] = dma_way_mask_expanded[37] & data_mem_w_mask_way_picked[5];
  assign data_mem_w_mask_o[36] = dma_way_mask_expanded[36] & data_mem_w_mask_way_picked[4];
  assign data_mem_w_mask_o[35] = dma_way_mask_expanded[35] & data_mem_w_mask_way_picked[3];
  assign data_mem_w_mask_o[34] = dma_way_mask_expanded[34] & data_mem_w_mask_way_picked[2];
  assign data_mem_w_mask_o[33] = dma_way_mask_expanded[33] & data_mem_w_mask_way_picked[1];
  assign data_mem_w_mask_o[32] = dma_way_mask_expanded[32] & data_mem_w_mask_way_picked[0];
  assign data_mem_w_mask_o[31] = dma_way_mask_expanded[31] & data_mem_w_mask_way_picked[15];
  assign data_mem_w_mask_o[30] = dma_way_mask_expanded[30] & data_mem_w_mask_way_picked[14];
  assign data_mem_w_mask_o[29] = dma_way_mask_expanded[29] & data_mem_w_mask_way_picked[13];
  assign data_mem_w_mask_o[28] = dma_way_mask_expanded[28] & data_mem_w_mask_way_picked[12];
  assign data_mem_w_mask_o[27] = dma_way_mask_expanded[27] & data_mem_w_mask_way_picked[11];
  assign data_mem_w_mask_o[26] = dma_way_mask_expanded[26] & data_mem_w_mask_way_picked[10];
  assign data_mem_w_mask_o[25] = dma_way_mask_expanded[25] & data_mem_w_mask_way_picked[9];
  assign data_mem_w_mask_o[24] = dma_way_mask_expanded[24] & data_mem_w_mask_way_picked[8];
  assign data_mem_w_mask_o[23] = dma_way_mask_expanded[23] & data_mem_w_mask_way_picked[7];
  assign data_mem_w_mask_o[22] = dma_way_mask_expanded[22] & data_mem_w_mask_way_picked[6];
  assign data_mem_w_mask_o[21] = dma_way_mask_expanded[21] & data_mem_w_mask_way_picked[5];
  assign data_mem_w_mask_o[20] = dma_way_mask_expanded[20] & data_mem_w_mask_way_picked[4];
  assign data_mem_w_mask_o[19] = dma_way_mask_expanded[19] & data_mem_w_mask_way_picked[3];
  assign data_mem_w_mask_o[18] = dma_way_mask_expanded[18] & data_mem_w_mask_way_picked[2];
  assign data_mem_w_mask_o[17] = dma_way_mask_expanded[17] & data_mem_w_mask_way_picked[1];
  assign data_mem_w_mask_o[16] = dma_way_mask_expanded[16] & data_mem_w_mask_way_picked[0];
  assign data_mem_w_mask_o[15] = dma_way_mask_expanded[15] & data_mem_w_mask_way_picked[15];
  assign data_mem_w_mask_o[14] = dma_way_mask_expanded[14] & data_mem_w_mask_way_picked[14];
  assign data_mem_w_mask_o[13] = dma_way_mask_expanded[13] & data_mem_w_mask_way_picked[13];
  assign data_mem_w_mask_o[12] = dma_way_mask_expanded[12] & data_mem_w_mask_way_picked[12];
  assign data_mem_w_mask_o[11] = dma_way_mask_expanded[11] & data_mem_w_mask_way_picked[11];
  assign data_mem_w_mask_o[10] = dma_way_mask_expanded[10] & data_mem_w_mask_way_picked[10];
  assign data_mem_w_mask_o[9] = dma_way_mask_expanded[9] & data_mem_w_mask_way_picked[9];
  assign data_mem_w_mask_o[8] = dma_way_mask_expanded[8] & data_mem_w_mask_way_picked[8];
  assign data_mem_w_mask_o[7] = dma_way_mask_expanded[7] & data_mem_w_mask_way_picked[7];
  assign data_mem_w_mask_o[6] = dma_way_mask_expanded[6] & data_mem_w_mask_way_picked[6];
  assign data_mem_w_mask_o[5] = dma_way_mask_expanded[5] & data_mem_w_mask_way_picked[5];
  assign data_mem_w_mask_o[4] = dma_way_mask_expanded[4] & data_mem_w_mask_way_picked[4];
  assign data_mem_w_mask_o[3] = dma_way_mask_expanded[3] & data_mem_w_mask_way_picked[3];
  assign data_mem_w_mask_o[2] = dma_way_mask_expanded[2] & data_mem_w_mask_way_picked[2];
  assign data_mem_w_mask_o[1] = dma_way_mask_expanded[1] & data_mem_w_mask_way_picked[1];
  assign data_mem_w_mask_o[0] = dma_way_mask_expanded[0] & data_mem_w_mask_way_picked[0];
  assign N29 = ~dma_state_r[1];
  assign N32 = ~N31;
  assign N34 = ~N33;
  assign N38 = ~N37;
  assign N42 = ~N41;
  assign N45 = ~N44;
  assign N49 = ~N48;
  assign N50 = ~dma_cmd_i[3];
  assign N51 = ~dma_cmd_i[2];
  assign N52 = ~dma_cmd_i[1];
  assign N53 = ~dma_cmd_i[0];
  assign N57 = N42 | N38;
  assign N58 = N45 | N57;
  assign N59 = N49 | N58;
  assign N60 = N56 | N59;
  assign N61 = ~N60;
  assign N72 = N97 & in_fifo_v_lo;
  assign N74 = in_fifo_v_lo & N96;
  assign N75 = in_fifo_v_lo & N97;
  assign N76 = N97 & in_fifo_v_lo;
  assign N77 = N92 & out_fifo_ready_lo;
  assign N79 = out_fifo_ready_lo & N91;
  assign N80 = out_fifo_ready_lo & N92;
  assign N81 = N101 & track_bits_offset_picked[0];
  assign N101 = out_fifo_ready_lo & N91;
  assign N82 = N92 & out_fifo_ready_lo;
  assign snoop_word_we = N102 & N83;
  assign N102 = N100 & in_fifo_v_lo;
  assign N84 = ~reset_i;
  assign N85 = reset_i;

  always @(posedge clk_i) begin
    if(N88) begin
      track_mem_data_r_31_sv2v_reg <= track_mem_data_i[31];
      track_mem_data_r_30_sv2v_reg <= track_mem_data_i[30];
      track_mem_data_r_29_sv2v_reg <= track_mem_data_i[29];
      track_mem_data_r_28_sv2v_reg <= track_mem_data_i[28];
      track_mem_data_r_27_sv2v_reg <= track_mem_data_i[27];
      track_mem_data_r_26_sv2v_reg <= track_mem_data_i[26];
      track_mem_data_r_25_sv2v_reg <= track_mem_data_i[25];
      track_mem_data_r_24_sv2v_reg <= track_mem_data_i[24];
      track_mem_data_r_23_sv2v_reg <= track_mem_data_i[23];
      track_mem_data_r_22_sv2v_reg <= track_mem_data_i[22];
      track_mem_data_r_21_sv2v_reg <= track_mem_data_i[21];
      track_mem_data_r_20_sv2v_reg <= track_mem_data_i[20];
      track_mem_data_r_19_sv2v_reg <= track_mem_data_i[19];
      track_mem_data_r_18_sv2v_reg <= track_mem_data_i[18];
      track_mem_data_r_17_sv2v_reg <= track_mem_data_i[17];
      track_mem_data_r_16_sv2v_reg <= track_mem_data_i[16];
      track_mem_data_r_15_sv2v_reg <= track_mem_data_i[15];
      track_mem_data_r_14_sv2v_reg <= track_mem_data_i[14];
      track_mem_data_r_13_sv2v_reg <= track_mem_data_i[13];
      track_mem_data_r_12_sv2v_reg <= track_mem_data_i[12];
      track_mem_data_r_11_sv2v_reg <= track_mem_data_i[11];
      track_mem_data_r_10_sv2v_reg <= track_mem_data_i[10];
      track_mem_data_r_9_sv2v_reg <= track_mem_data_i[9];
      track_mem_data_r_8_sv2v_reg <= track_mem_data_i[8];
      track_mem_data_r_7_sv2v_reg <= track_mem_data_i[7];
      track_mem_data_r_6_sv2v_reg <= track_mem_data_i[6];
      track_mem_data_r_5_sv2v_reg <= track_mem_data_i[5];
      track_mem_data_r_4_sv2v_reg <= track_mem_data_i[4];
      track_mem_data_r_3_sv2v_reg <= track_mem_data_i[3];
      track_mem_data_r_2_sv2v_reg <= track_mem_data_i[2];
      track_mem_data_r_1_sv2v_reg <= track_mem_data_i[1];
      track_mem_data_r_0_sv2v_reg <= track_mem_data_i[0];
    end 
    if(reset_i) begin
      dma_state_r_1_sv2v_reg <= 1'b0;
      dma_state_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      dma_state_r_1_sv2v_reg <= dma_state_n[1];
      dma_state_r_0_sv2v_reg <= dma_state_n[0];
    end 
    if(N86) begin
      snoop_word_o_127_sv2v_reg <= snoop_word_n[127];
      snoop_word_o_126_sv2v_reg <= snoop_word_n[126];
      snoop_word_o_125_sv2v_reg <= snoop_word_n[125];
      snoop_word_o_124_sv2v_reg <= snoop_word_n[124];
      snoop_word_o_123_sv2v_reg <= snoop_word_n[123];
      snoop_word_o_122_sv2v_reg <= snoop_word_n[122];
      snoop_word_o_121_sv2v_reg <= snoop_word_n[121];
      snoop_word_o_120_sv2v_reg <= snoop_word_n[120];
      snoop_word_o_119_sv2v_reg <= snoop_word_n[119];
      snoop_word_o_118_sv2v_reg <= snoop_word_n[118];
      snoop_word_o_117_sv2v_reg <= snoop_word_n[117];
      snoop_word_o_116_sv2v_reg <= snoop_word_n[116];
      snoop_word_o_115_sv2v_reg <= snoop_word_n[115];
      snoop_word_o_114_sv2v_reg <= snoop_word_n[114];
      snoop_word_o_113_sv2v_reg <= snoop_word_n[113];
      snoop_word_o_112_sv2v_reg <= snoop_word_n[112];
      snoop_word_o_111_sv2v_reg <= snoop_word_n[111];
      snoop_word_o_110_sv2v_reg <= snoop_word_n[110];
      snoop_word_o_109_sv2v_reg <= snoop_word_n[109];
      snoop_word_o_108_sv2v_reg <= snoop_word_n[108];
      snoop_word_o_107_sv2v_reg <= snoop_word_n[107];
      snoop_word_o_106_sv2v_reg <= snoop_word_n[106];
      snoop_word_o_105_sv2v_reg <= snoop_word_n[105];
      snoop_word_o_104_sv2v_reg <= snoop_word_n[104];
      snoop_word_o_103_sv2v_reg <= snoop_word_n[103];
      snoop_word_o_102_sv2v_reg <= snoop_word_n[102];
      snoop_word_o_101_sv2v_reg <= snoop_word_n[101];
      snoop_word_o_100_sv2v_reg <= snoop_word_n[100];
      snoop_word_o_99_sv2v_reg <= snoop_word_n[99];
      snoop_word_o_98_sv2v_reg <= snoop_word_n[98];
      snoop_word_o_97_sv2v_reg <= snoop_word_n[97];
      snoop_word_o_96_sv2v_reg <= snoop_word_n[96];
      snoop_word_o_95_sv2v_reg <= snoop_word_n[95];
      snoop_word_o_94_sv2v_reg <= snoop_word_n[94];
      snoop_word_o_93_sv2v_reg <= snoop_word_n[93];
      snoop_word_o_92_sv2v_reg <= snoop_word_n[92];
      snoop_word_o_91_sv2v_reg <= snoop_word_n[91];
      snoop_word_o_90_sv2v_reg <= snoop_word_n[90];
      snoop_word_o_89_sv2v_reg <= snoop_word_n[89];
      snoop_word_o_88_sv2v_reg <= snoop_word_n[88];
      snoop_word_o_87_sv2v_reg <= snoop_word_n[87];
      snoop_word_o_86_sv2v_reg <= snoop_word_n[86];
      snoop_word_o_85_sv2v_reg <= snoop_word_n[85];
      snoop_word_o_84_sv2v_reg <= snoop_word_n[84];
      snoop_word_o_83_sv2v_reg <= snoop_word_n[83];
      snoop_word_o_82_sv2v_reg <= snoop_word_n[82];
      snoop_word_o_81_sv2v_reg <= snoop_word_n[81];
      snoop_word_o_80_sv2v_reg <= snoop_word_n[80];
      snoop_word_o_79_sv2v_reg <= snoop_word_n[79];
      snoop_word_o_78_sv2v_reg <= snoop_word_n[78];
      snoop_word_o_77_sv2v_reg <= snoop_word_n[77];
      snoop_word_o_76_sv2v_reg <= snoop_word_n[76];
      snoop_word_o_75_sv2v_reg <= snoop_word_n[75];
      snoop_word_o_74_sv2v_reg <= snoop_word_n[74];
      snoop_word_o_73_sv2v_reg <= snoop_word_n[73];
      snoop_word_o_72_sv2v_reg <= snoop_word_n[72];
      snoop_word_o_71_sv2v_reg <= snoop_word_n[71];
      snoop_word_o_70_sv2v_reg <= snoop_word_n[70];
      snoop_word_o_69_sv2v_reg <= snoop_word_n[69];
      snoop_word_o_68_sv2v_reg <= snoop_word_n[68];
      snoop_word_o_67_sv2v_reg <= snoop_word_n[67];
      snoop_word_o_66_sv2v_reg <= snoop_word_n[66];
      snoop_word_o_65_sv2v_reg <= snoop_word_n[65];
      snoop_word_o_64_sv2v_reg <= snoop_word_n[64];
      snoop_word_o_63_sv2v_reg <= snoop_word_n[63];
      snoop_word_o_62_sv2v_reg <= snoop_word_n[62];
      snoop_word_o_61_sv2v_reg <= snoop_word_n[61];
      snoop_word_o_60_sv2v_reg <= snoop_word_n[60];
      snoop_word_o_59_sv2v_reg <= snoop_word_n[59];
      snoop_word_o_58_sv2v_reg <= snoop_word_n[58];
      snoop_word_o_57_sv2v_reg <= snoop_word_n[57];
      snoop_word_o_56_sv2v_reg <= snoop_word_n[56];
      snoop_word_o_55_sv2v_reg <= snoop_word_n[55];
      snoop_word_o_54_sv2v_reg <= snoop_word_n[54];
      snoop_word_o_53_sv2v_reg <= snoop_word_n[53];
      snoop_word_o_52_sv2v_reg <= snoop_word_n[52];
      snoop_word_o_51_sv2v_reg <= snoop_word_n[51];
      snoop_word_o_50_sv2v_reg <= snoop_word_n[50];
      snoop_word_o_49_sv2v_reg <= snoop_word_n[49];
      snoop_word_o_48_sv2v_reg <= snoop_word_n[48];
      snoop_word_o_47_sv2v_reg <= snoop_word_n[47];
      snoop_word_o_46_sv2v_reg <= snoop_word_n[46];
      snoop_word_o_45_sv2v_reg <= snoop_word_n[45];
      snoop_word_o_44_sv2v_reg <= snoop_word_n[44];
      snoop_word_o_43_sv2v_reg <= snoop_word_n[43];
      snoop_word_o_42_sv2v_reg <= snoop_word_n[42];
      snoop_word_o_41_sv2v_reg <= snoop_word_n[41];
      snoop_word_o_40_sv2v_reg <= snoop_word_n[40];
      snoop_word_o_39_sv2v_reg <= snoop_word_n[39];
      snoop_word_o_38_sv2v_reg <= snoop_word_n[38];
      snoop_word_o_37_sv2v_reg <= snoop_word_n[37];
      snoop_word_o_36_sv2v_reg <= snoop_word_n[36];
      snoop_word_o_35_sv2v_reg <= snoop_word_n[35];
      snoop_word_o_34_sv2v_reg <= snoop_word_n[34];
      snoop_word_o_33_sv2v_reg <= snoop_word_n[33];
      snoop_word_o_32_sv2v_reg <= snoop_word_n[32];
      snoop_word_o_31_sv2v_reg <= snoop_word_n[31];
      snoop_word_o_30_sv2v_reg <= snoop_word_n[30];
      snoop_word_o_29_sv2v_reg <= snoop_word_n[29];
      snoop_word_o_0_sv2v_reg <= snoop_word_n[0];
    end 
    if(N87) begin
      snoop_word_o_28_sv2v_reg <= snoop_word_n[28];
      snoop_word_o_27_sv2v_reg <= snoop_word_n[27];
      snoop_word_o_26_sv2v_reg <= snoop_word_n[26];
      snoop_word_o_25_sv2v_reg <= snoop_word_n[25];
      snoop_word_o_24_sv2v_reg <= snoop_word_n[24];
      snoop_word_o_23_sv2v_reg <= snoop_word_n[23];
      snoop_word_o_22_sv2v_reg <= snoop_word_n[22];
      snoop_word_o_21_sv2v_reg <= snoop_word_n[21];
      snoop_word_o_20_sv2v_reg <= snoop_word_n[20];
      snoop_word_o_19_sv2v_reg <= snoop_word_n[19];
      snoop_word_o_18_sv2v_reg <= snoop_word_n[18];
      snoop_word_o_17_sv2v_reg <= snoop_word_n[17];
      snoop_word_o_16_sv2v_reg <= snoop_word_n[16];
      snoop_word_o_15_sv2v_reg <= snoop_word_n[15];
      snoop_word_o_14_sv2v_reg <= snoop_word_n[14];
      snoop_word_o_13_sv2v_reg <= snoop_word_n[13];
      snoop_word_o_12_sv2v_reg <= snoop_word_n[12];
      snoop_word_o_11_sv2v_reg <= snoop_word_n[11];
      snoop_word_o_10_sv2v_reg <= snoop_word_n[10];
      snoop_word_o_9_sv2v_reg <= snoop_word_n[9];
      snoop_word_o_8_sv2v_reg <= snoop_word_n[8];
      snoop_word_o_7_sv2v_reg <= snoop_word_n[7];
      snoop_word_o_6_sv2v_reg <= snoop_word_n[6];
      snoop_word_o_5_sv2v_reg <= snoop_word_n[5];
      snoop_word_o_4_sv2v_reg <= snoop_word_n[4];
      snoop_word_o_3_sv2v_reg <= snoop_word_n[3];
      snoop_word_o_2_sv2v_reg <= snoop_word_n[2];
      snoop_word_o_1_sv2v_reg <= snoop_word_n[1];
    end 
  end


endmodule



module bsg_cache_buffer_queue_000000b4
(
  clk_i,
  reset_i,
  v_i,
  data_i,
  v_o,
  data_o,
  yumi_i,
  el0_valid_o,
  el1_valid_o,
  el0_snoop_o,
  el1_snoop_o,
  empty_o,
  full_o
);

  input [179:0] data_i;
  output [179:0] data_o;
  output [179:0] el0_snoop_o;
  output [179:0] el1_snoop_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output v_o;
  output el0_valid_o;
  output el1_valid_o;
  output empty_o;
  output full_o;
  wire [179:0] data_o,el0_snoop_o,el1_snoop_o;
  wire v_o,el0_valid_o,el1_valid_o,empty_o,full_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,
  N11,N12,N13,N14,N15,el0_enable,el1_enable,mux0_sel,mux1_sel,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,
  N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,
  N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,
  N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,
  N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,
  N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,
  N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
  N197,N198,N199,N200,N201,N202,N203,N204,N205,N206;
  wire [1:0] num_els_r;
  reg num_els_r_1_sv2v_reg,num_els_r_0_sv2v_reg,el0_snoop_o_179_sv2v_reg,
  el0_snoop_o_178_sv2v_reg,el0_snoop_o_177_sv2v_reg,el0_snoop_o_176_sv2v_reg,
  el0_snoop_o_175_sv2v_reg,el0_snoop_o_174_sv2v_reg,el0_snoop_o_173_sv2v_reg,
  el0_snoop_o_172_sv2v_reg,el0_snoop_o_171_sv2v_reg,el0_snoop_o_170_sv2v_reg,el0_snoop_o_169_sv2v_reg,
  el0_snoop_o_168_sv2v_reg,el0_snoop_o_167_sv2v_reg,el0_snoop_o_166_sv2v_reg,
  el0_snoop_o_165_sv2v_reg,el0_snoop_o_164_sv2v_reg,el0_snoop_o_163_sv2v_reg,
  el0_snoop_o_162_sv2v_reg,el0_snoop_o_161_sv2v_reg,el0_snoop_o_160_sv2v_reg,
  el0_snoop_o_159_sv2v_reg,el0_snoop_o_158_sv2v_reg,el0_snoop_o_157_sv2v_reg,
  el0_snoop_o_156_sv2v_reg,el0_snoop_o_155_sv2v_reg,el0_snoop_o_154_sv2v_reg,el0_snoop_o_153_sv2v_reg,
  el0_snoop_o_152_sv2v_reg,el0_snoop_o_151_sv2v_reg,el0_snoop_o_150_sv2v_reg,
  el0_snoop_o_149_sv2v_reg,el0_snoop_o_148_sv2v_reg,el0_snoop_o_147_sv2v_reg,
  el0_snoop_o_146_sv2v_reg,el0_snoop_o_145_sv2v_reg,el0_snoop_o_144_sv2v_reg,
  el0_snoop_o_143_sv2v_reg,el0_snoop_o_142_sv2v_reg,el0_snoop_o_141_sv2v_reg,
  el0_snoop_o_140_sv2v_reg,el0_snoop_o_139_sv2v_reg,el0_snoop_o_138_sv2v_reg,el0_snoop_o_137_sv2v_reg,
  el0_snoop_o_136_sv2v_reg,el0_snoop_o_135_sv2v_reg,el0_snoop_o_134_sv2v_reg,
  el0_snoop_o_133_sv2v_reg,el0_snoop_o_132_sv2v_reg,el0_snoop_o_131_sv2v_reg,
  el0_snoop_o_130_sv2v_reg,el0_snoop_o_129_sv2v_reg,el0_snoop_o_128_sv2v_reg,
  el0_snoop_o_127_sv2v_reg,el0_snoop_o_126_sv2v_reg,el0_snoop_o_125_sv2v_reg,
  el0_snoop_o_124_sv2v_reg,el0_snoop_o_123_sv2v_reg,el0_snoop_o_122_sv2v_reg,el0_snoop_o_121_sv2v_reg,
  el0_snoop_o_120_sv2v_reg,el0_snoop_o_119_sv2v_reg,el0_snoop_o_118_sv2v_reg,
  el0_snoop_o_117_sv2v_reg,el0_snoop_o_116_sv2v_reg,el0_snoop_o_115_sv2v_reg,
  el0_snoop_o_114_sv2v_reg,el0_snoop_o_113_sv2v_reg,el0_snoop_o_112_sv2v_reg,
  el0_snoop_o_111_sv2v_reg,el0_snoop_o_110_sv2v_reg,el0_snoop_o_109_sv2v_reg,
  el0_snoop_o_108_sv2v_reg,el0_snoop_o_107_sv2v_reg,el0_snoop_o_106_sv2v_reg,el0_snoop_o_105_sv2v_reg,
  el0_snoop_o_104_sv2v_reg,el0_snoop_o_103_sv2v_reg,el0_snoop_o_102_sv2v_reg,
  el0_snoop_o_101_sv2v_reg,el0_snoop_o_100_sv2v_reg,el0_snoop_o_99_sv2v_reg,
  el0_snoop_o_98_sv2v_reg,el0_snoop_o_97_sv2v_reg,el0_snoop_o_96_sv2v_reg,
  el0_snoop_o_95_sv2v_reg,el0_snoop_o_94_sv2v_reg,el0_snoop_o_93_sv2v_reg,el0_snoop_o_92_sv2v_reg,
  el0_snoop_o_91_sv2v_reg,el0_snoop_o_90_sv2v_reg,el0_snoop_o_89_sv2v_reg,
  el0_snoop_o_88_sv2v_reg,el0_snoop_o_87_sv2v_reg,el0_snoop_o_86_sv2v_reg,
  el0_snoop_o_85_sv2v_reg,el0_snoop_o_84_sv2v_reg,el0_snoop_o_83_sv2v_reg,el0_snoop_o_82_sv2v_reg,
  el0_snoop_o_81_sv2v_reg,el0_snoop_o_80_sv2v_reg,el0_snoop_o_79_sv2v_reg,
  el0_snoop_o_78_sv2v_reg,el0_snoop_o_77_sv2v_reg,el0_snoop_o_76_sv2v_reg,
  el0_snoop_o_75_sv2v_reg,el0_snoop_o_74_sv2v_reg,el0_snoop_o_73_sv2v_reg,el0_snoop_o_72_sv2v_reg,
  el0_snoop_o_71_sv2v_reg,el0_snoop_o_70_sv2v_reg,el0_snoop_o_69_sv2v_reg,
  el0_snoop_o_68_sv2v_reg,el0_snoop_o_67_sv2v_reg,el0_snoop_o_66_sv2v_reg,
  el0_snoop_o_65_sv2v_reg,el0_snoop_o_64_sv2v_reg,el0_snoop_o_63_sv2v_reg,el0_snoop_o_62_sv2v_reg,
  el0_snoop_o_61_sv2v_reg,el0_snoop_o_60_sv2v_reg,el0_snoop_o_59_sv2v_reg,
  el0_snoop_o_58_sv2v_reg,el0_snoop_o_57_sv2v_reg,el0_snoop_o_56_sv2v_reg,
  el0_snoop_o_55_sv2v_reg,el0_snoop_o_54_sv2v_reg,el0_snoop_o_53_sv2v_reg,el0_snoop_o_52_sv2v_reg,
  el0_snoop_o_51_sv2v_reg,el0_snoop_o_50_sv2v_reg,el0_snoop_o_49_sv2v_reg,
  el0_snoop_o_48_sv2v_reg,el0_snoop_o_47_sv2v_reg,el0_snoop_o_46_sv2v_reg,
  el0_snoop_o_45_sv2v_reg,el0_snoop_o_44_sv2v_reg,el0_snoop_o_43_sv2v_reg,el0_snoop_o_42_sv2v_reg,
  el0_snoop_o_41_sv2v_reg,el0_snoop_o_40_sv2v_reg,el0_snoop_o_39_sv2v_reg,
  el0_snoop_o_38_sv2v_reg,el0_snoop_o_37_sv2v_reg,el0_snoop_o_36_sv2v_reg,
  el0_snoop_o_35_sv2v_reg,el0_snoop_o_34_sv2v_reg,el0_snoop_o_33_sv2v_reg,el0_snoop_o_32_sv2v_reg,
  el0_snoop_o_31_sv2v_reg,el0_snoop_o_30_sv2v_reg,el0_snoop_o_29_sv2v_reg,
  el0_snoop_o_28_sv2v_reg,el0_snoop_o_27_sv2v_reg,el0_snoop_o_26_sv2v_reg,
  el0_snoop_o_25_sv2v_reg,el0_snoop_o_24_sv2v_reg,el0_snoop_o_23_sv2v_reg,el0_snoop_o_22_sv2v_reg,
  el0_snoop_o_21_sv2v_reg,el0_snoop_o_20_sv2v_reg,el0_snoop_o_19_sv2v_reg,
  el0_snoop_o_18_sv2v_reg,el0_snoop_o_17_sv2v_reg,el0_snoop_o_16_sv2v_reg,
  el0_snoop_o_15_sv2v_reg,el0_snoop_o_14_sv2v_reg,el0_snoop_o_13_sv2v_reg,el0_snoop_o_12_sv2v_reg,
  el0_snoop_o_11_sv2v_reg,el0_snoop_o_10_sv2v_reg,el0_snoop_o_9_sv2v_reg,
  el0_snoop_o_8_sv2v_reg,el0_snoop_o_7_sv2v_reg,el0_snoop_o_6_sv2v_reg,el0_snoop_o_5_sv2v_reg,
  el0_snoop_o_4_sv2v_reg,el0_snoop_o_3_sv2v_reg,el0_snoop_o_2_sv2v_reg,
  el0_snoop_o_1_sv2v_reg,el0_snoop_o_0_sv2v_reg,el1_snoop_o_179_sv2v_reg,
  el1_snoop_o_178_sv2v_reg,el1_snoop_o_177_sv2v_reg,el1_snoop_o_176_sv2v_reg,el1_snoop_o_175_sv2v_reg,
  el1_snoop_o_174_sv2v_reg,el1_snoop_o_173_sv2v_reg,el1_snoop_o_172_sv2v_reg,
  el1_snoop_o_171_sv2v_reg,el1_snoop_o_170_sv2v_reg,el1_snoop_o_169_sv2v_reg,
  el1_snoop_o_168_sv2v_reg,el1_snoop_o_167_sv2v_reg,el1_snoop_o_166_sv2v_reg,
  el1_snoop_o_165_sv2v_reg,el1_snoop_o_164_sv2v_reg,el1_snoop_o_163_sv2v_reg,
  el1_snoop_o_162_sv2v_reg,el1_snoop_o_161_sv2v_reg,el1_snoop_o_160_sv2v_reg,el1_snoop_o_159_sv2v_reg,
  el1_snoop_o_158_sv2v_reg,el1_snoop_o_157_sv2v_reg,el1_snoop_o_156_sv2v_reg,
  el1_snoop_o_155_sv2v_reg,el1_snoop_o_154_sv2v_reg,el1_snoop_o_153_sv2v_reg,
  el1_snoop_o_152_sv2v_reg,el1_snoop_o_151_sv2v_reg,el1_snoop_o_150_sv2v_reg,
  el1_snoop_o_149_sv2v_reg,el1_snoop_o_148_sv2v_reg,el1_snoop_o_147_sv2v_reg,
  el1_snoop_o_146_sv2v_reg,el1_snoop_o_145_sv2v_reg,el1_snoop_o_144_sv2v_reg,el1_snoop_o_143_sv2v_reg,
  el1_snoop_o_142_sv2v_reg,el1_snoop_o_141_sv2v_reg,el1_snoop_o_140_sv2v_reg,
  el1_snoop_o_139_sv2v_reg,el1_snoop_o_138_sv2v_reg,el1_snoop_o_137_sv2v_reg,
  el1_snoop_o_136_sv2v_reg,el1_snoop_o_135_sv2v_reg,el1_snoop_o_134_sv2v_reg,
  el1_snoop_o_133_sv2v_reg,el1_snoop_o_132_sv2v_reg,el1_snoop_o_131_sv2v_reg,
  el1_snoop_o_130_sv2v_reg,el1_snoop_o_129_sv2v_reg,el1_snoop_o_128_sv2v_reg,el1_snoop_o_127_sv2v_reg,
  el1_snoop_o_126_sv2v_reg,el1_snoop_o_125_sv2v_reg,el1_snoop_o_124_sv2v_reg,
  el1_snoop_o_123_sv2v_reg,el1_snoop_o_122_sv2v_reg,el1_snoop_o_121_sv2v_reg,
  el1_snoop_o_120_sv2v_reg,el1_snoop_o_119_sv2v_reg,el1_snoop_o_118_sv2v_reg,
  el1_snoop_o_117_sv2v_reg,el1_snoop_o_116_sv2v_reg,el1_snoop_o_115_sv2v_reg,
  el1_snoop_o_114_sv2v_reg,el1_snoop_o_113_sv2v_reg,el1_snoop_o_112_sv2v_reg,el1_snoop_o_111_sv2v_reg,
  el1_snoop_o_110_sv2v_reg,el1_snoop_o_109_sv2v_reg,el1_snoop_o_108_sv2v_reg,
  el1_snoop_o_107_sv2v_reg,el1_snoop_o_106_sv2v_reg,el1_snoop_o_105_sv2v_reg,
  el1_snoop_o_104_sv2v_reg,el1_snoop_o_103_sv2v_reg,el1_snoop_o_102_sv2v_reg,
  el1_snoop_o_101_sv2v_reg,el1_snoop_o_100_sv2v_reg,el1_snoop_o_99_sv2v_reg,el1_snoop_o_98_sv2v_reg,
  el1_snoop_o_97_sv2v_reg,el1_snoop_o_96_sv2v_reg,el1_snoop_o_95_sv2v_reg,
  el1_snoop_o_94_sv2v_reg,el1_snoop_o_93_sv2v_reg,el1_snoop_o_92_sv2v_reg,
  el1_snoop_o_91_sv2v_reg,el1_snoop_o_90_sv2v_reg,el1_snoop_o_89_sv2v_reg,el1_snoop_o_88_sv2v_reg,
  el1_snoop_o_87_sv2v_reg,el1_snoop_o_86_sv2v_reg,el1_snoop_o_85_sv2v_reg,
  el1_snoop_o_84_sv2v_reg,el1_snoop_o_83_sv2v_reg,el1_snoop_o_82_sv2v_reg,
  el1_snoop_o_81_sv2v_reg,el1_snoop_o_80_sv2v_reg,el1_snoop_o_79_sv2v_reg,el1_snoop_o_78_sv2v_reg,
  el1_snoop_o_77_sv2v_reg,el1_snoop_o_76_sv2v_reg,el1_snoop_o_75_sv2v_reg,
  el1_snoop_o_74_sv2v_reg,el1_snoop_o_73_sv2v_reg,el1_snoop_o_72_sv2v_reg,
  el1_snoop_o_71_sv2v_reg,el1_snoop_o_70_sv2v_reg,el1_snoop_o_69_sv2v_reg,el1_snoop_o_68_sv2v_reg,
  el1_snoop_o_67_sv2v_reg,el1_snoop_o_66_sv2v_reg,el1_snoop_o_65_sv2v_reg,
  el1_snoop_o_64_sv2v_reg,el1_snoop_o_63_sv2v_reg,el1_snoop_o_62_sv2v_reg,
  el1_snoop_o_61_sv2v_reg,el1_snoop_o_60_sv2v_reg,el1_snoop_o_59_sv2v_reg,el1_snoop_o_58_sv2v_reg,
  el1_snoop_o_57_sv2v_reg,el1_snoop_o_56_sv2v_reg,el1_snoop_o_55_sv2v_reg,
  el1_snoop_o_54_sv2v_reg,el1_snoop_o_53_sv2v_reg,el1_snoop_o_52_sv2v_reg,
  el1_snoop_o_51_sv2v_reg,el1_snoop_o_50_sv2v_reg,el1_snoop_o_49_sv2v_reg,el1_snoop_o_48_sv2v_reg,
  el1_snoop_o_47_sv2v_reg,el1_snoop_o_46_sv2v_reg,el1_snoop_o_45_sv2v_reg,
  el1_snoop_o_44_sv2v_reg,el1_snoop_o_43_sv2v_reg,el1_snoop_o_42_sv2v_reg,
  el1_snoop_o_41_sv2v_reg,el1_snoop_o_40_sv2v_reg,el1_snoop_o_39_sv2v_reg,el1_snoop_o_38_sv2v_reg,
  el1_snoop_o_37_sv2v_reg,el1_snoop_o_36_sv2v_reg,el1_snoop_o_35_sv2v_reg,
  el1_snoop_o_34_sv2v_reg,el1_snoop_o_33_sv2v_reg,el1_snoop_o_32_sv2v_reg,
  el1_snoop_o_31_sv2v_reg,el1_snoop_o_30_sv2v_reg,el1_snoop_o_29_sv2v_reg,el1_snoop_o_28_sv2v_reg,
  el1_snoop_o_27_sv2v_reg,el1_snoop_o_26_sv2v_reg,el1_snoop_o_25_sv2v_reg,
  el1_snoop_o_24_sv2v_reg,el1_snoop_o_23_sv2v_reg,el1_snoop_o_22_sv2v_reg,
  el1_snoop_o_21_sv2v_reg,el1_snoop_o_20_sv2v_reg,el1_snoop_o_19_sv2v_reg,el1_snoop_o_18_sv2v_reg,
  el1_snoop_o_17_sv2v_reg,el1_snoop_o_16_sv2v_reg,el1_snoop_o_15_sv2v_reg,
  el1_snoop_o_14_sv2v_reg,el1_snoop_o_13_sv2v_reg,el1_snoop_o_12_sv2v_reg,
  el1_snoop_o_11_sv2v_reg,el1_snoop_o_10_sv2v_reg,el1_snoop_o_9_sv2v_reg,el1_snoop_o_8_sv2v_reg,
  el1_snoop_o_7_sv2v_reg,el1_snoop_o_6_sv2v_reg,el1_snoop_o_5_sv2v_reg,
  el1_snoop_o_4_sv2v_reg,el1_snoop_o_3_sv2v_reg,el1_snoop_o_2_sv2v_reg,el1_snoop_o_1_sv2v_reg,
  el1_snoop_o_0_sv2v_reg;
  assign num_els_r[1] = num_els_r_1_sv2v_reg;
  assign num_els_r[0] = num_els_r_0_sv2v_reg;
  assign el0_snoop_o[179] = el0_snoop_o_179_sv2v_reg;
  assign el0_snoop_o[178] = el0_snoop_o_178_sv2v_reg;
  assign el0_snoop_o[177] = el0_snoop_o_177_sv2v_reg;
  assign el0_snoop_o[176] = el0_snoop_o_176_sv2v_reg;
  assign el0_snoop_o[175] = el0_snoop_o_175_sv2v_reg;
  assign el0_snoop_o[174] = el0_snoop_o_174_sv2v_reg;
  assign el0_snoop_o[173] = el0_snoop_o_173_sv2v_reg;
  assign el0_snoop_o[172] = el0_snoop_o_172_sv2v_reg;
  assign el0_snoop_o[171] = el0_snoop_o_171_sv2v_reg;
  assign el0_snoop_o[170] = el0_snoop_o_170_sv2v_reg;
  assign el0_snoop_o[169] = el0_snoop_o_169_sv2v_reg;
  assign el0_snoop_o[168] = el0_snoop_o_168_sv2v_reg;
  assign el0_snoop_o[167] = el0_snoop_o_167_sv2v_reg;
  assign el0_snoop_o[166] = el0_snoop_o_166_sv2v_reg;
  assign el0_snoop_o[165] = el0_snoop_o_165_sv2v_reg;
  assign el0_snoop_o[164] = el0_snoop_o_164_sv2v_reg;
  assign el0_snoop_o[163] = el0_snoop_o_163_sv2v_reg;
  assign el0_snoop_o[162] = el0_snoop_o_162_sv2v_reg;
  assign el0_snoop_o[161] = el0_snoop_o_161_sv2v_reg;
  assign el0_snoop_o[160] = el0_snoop_o_160_sv2v_reg;
  assign el0_snoop_o[159] = el0_snoop_o_159_sv2v_reg;
  assign el0_snoop_o[158] = el0_snoop_o_158_sv2v_reg;
  assign el0_snoop_o[157] = el0_snoop_o_157_sv2v_reg;
  assign el0_snoop_o[156] = el0_snoop_o_156_sv2v_reg;
  assign el0_snoop_o[155] = el0_snoop_o_155_sv2v_reg;
  assign el0_snoop_o[154] = el0_snoop_o_154_sv2v_reg;
  assign el0_snoop_o[153] = el0_snoop_o_153_sv2v_reg;
  assign el0_snoop_o[152] = el0_snoop_o_152_sv2v_reg;
  assign el0_snoop_o[151] = el0_snoop_o_151_sv2v_reg;
  assign el0_snoop_o[150] = el0_snoop_o_150_sv2v_reg;
  assign el0_snoop_o[149] = el0_snoop_o_149_sv2v_reg;
  assign el0_snoop_o[148] = el0_snoop_o_148_sv2v_reg;
  assign el0_snoop_o[147] = el0_snoop_o_147_sv2v_reg;
  assign el0_snoop_o[146] = el0_snoop_o_146_sv2v_reg;
  assign el0_snoop_o[145] = el0_snoop_o_145_sv2v_reg;
  assign el0_snoop_o[144] = el0_snoop_o_144_sv2v_reg;
  assign el0_snoop_o[143] = el0_snoop_o_143_sv2v_reg;
  assign el0_snoop_o[142] = el0_snoop_o_142_sv2v_reg;
  assign el0_snoop_o[141] = el0_snoop_o_141_sv2v_reg;
  assign el0_snoop_o[140] = el0_snoop_o_140_sv2v_reg;
  assign el0_snoop_o[139] = el0_snoop_o_139_sv2v_reg;
  assign el0_snoop_o[138] = el0_snoop_o_138_sv2v_reg;
  assign el0_snoop_o[137] = el0_snoop_o_137_sv2v_reg;
  assign el0_snoop_o[136] = el0_snoop_o_136_sv2v_reg;
  assign el0_snoop_o[135] = el0_snoop_o_135_sv2v_reg;
  assign el0_snoop_o[134] = el0_snoop_o_134_sv2v_reg;
  assign el0_snoop_o[133] = el0_snoop_o_133_sv2v_reg;
  assign el0_snoop_o[132] = el0_snoop_o_132_sv2v_reg;
  assign el0_snoop_o[131] = el0_snoop_o_131_sv2v_reg;
  assign el0_snoop_o[130] = el0_snoop_o_130_sv2v_reg;
  assign el0_snoop_o[129] = el0_snoop_o_129_sv2v_reg;
  assign el0_snoop_o[128] = el0_snoop_o_128_sv2v_reg;
  assign el0_snoop_o[127] = el0_snoop_o_127_sv2v_reg;
  assign el0_snoop_o[126] = el0_snoop_o_126_sv2v_reg;
  assign el0_snoop_o[125] = el0_snoop_o_125_sv2v_reg;
  assign el0_snoop_o[124] = el0_snoop_o_124_sv2v_reg;
  assign el0_snoop_o[123] = el0_snoop_o_123_sv2v_reg;
  assign el0_snoop_o[122] = el0_snoop_o_122_sv2v_reg;
  assign el0_snoop_o[121] = el0_snoop_o_121_sv2v_reg;
  assign el0_snoop_o[120] = el0_snoop_o_120_sv2v_reg;
  assign el0_snoop_o[119] = el0_snoop_o_119_sv2v_reg;
  assign el0_snoop_o[118] = el0_snoop_o_118_sv2v_reg;
  assign el0_snoop_o[117] = el0_snoop_o_117_sv2v_reg;
  assign el0_snoop_o[116] = el0_snoop_o_116_sv2v_reg;
  assign el0_snoop_o[115] = el0_snoop_o_115_sv2v_reg;
  assign el0_snoop_o[114] = el0_snoop_o_114_sv2v_reg;
  assign el0_snoop_o[113] = el0_snoop_o_113_sv2v_reg;
  assign el0_snoop_o[112] = el0_snoop_o_112_sv2v_reg;
  assign el0_snoop_o[111] = el0_snoop_o_111_sv2v_reg;
  assign el0_snoop_o[110] = el0_snoop_o_110_sv2v_reg;
  assign el0_snoop_o[109] = el0_snoop_o_109_sv2v_reg;
  assign el0_snoop_o[108] = el0_snoop_o_108_sv2v_reg;
  assign el0_snoop_o[107] = el0_snoop_o_107_sv2v_reg;
  assign el0_snoop_o[106] = el0_snoop_o_106_sv2v_reg;
  assign el0_snoop_o[105] = el0_snoop_o_105_sv2v_reg;
  assign el0_snoop_o[104] = el0_snoop_o_104_sv2v_reg;
  assign el0_snoop_o[103] = el0_snoop_o_103_sv2v_reg;
  assign el0_snoop_o[102] = el0_snoop_o_102_sv2v_reg;
  assign el0_snoop_o[101] = el0_snoop_o_101_sv2v_reg;
  assign el0_snoop_o[100] = el0_snoop_o_100_sv2v_reg;
  assign el0_snoop_o[99] = el0_snoop_o_99_sv2v_reg;
  assign el0_snoop_o[98] = el0_snoop_o_98_sv2v_reg;
  assign el0_snoop_o[97] = el0_snoop_o_97_sv2v_reg;
  assign el0_snoop_o[96] = el0_snoop_o_96_sv2v_reg;
  assign el0_snoop_o[95] = el0_snoop_o_95_sv2v_reg;
  assign el0_snoop_o[94] = el0_snoop_o_94_sv2v_reg;
  assign el0_snoop_o[93] = el0_snoop_o_93_sv2v_reg;
  assign el0_snoop_o[92] = el0_snoop_o_92_sv2v_reg;
  assign el0_snoop_o[91] = el0_snoop_o_91_sv2v_reg;
  assign el0_snoop_o[90] = el0_snoop_o_90_sv2v_reg;
  assign el0_snoop_o[89] = el0_snoop_o_89_sv2v_reg;
  assign el0_snoop_o[88] = el0_snoop_o_88_sv2v_reg;
  assign el0_snoop_o[87] = el0_snoop_o_87_sv2v_reg;
  assign el0_snoop_o[86] = el0_snoop_o_86_sv2v_reg;
  assign el0_snoop_o[85] = el0_snoop_o_85_sv2v_reg;
  assign el0_snoop_o[84] = el0_snoop_o_84_sv2v_reg;
  assign el0_snoop_o[83] = el0_snoop_o_83_sv2v_reg;
  assign el0_snoop_o[82] = el0_snoop_o_82_sv2v_reg;
  assign el0_snoop_o[81] = el0_snoop_o_81_sv2v_reg;
  assign el0_snoop_o[80] = el0_snoop_o_80_sv2v_reg;
  assign el0_snoop_o[79] = el0_snoop_o_79_sv2v_reg;
  assign el0_snoop_o[78] = el0_snoop_o_78_sv2v_reg;
  assign el0_snoop_o[77] = el0_snoop_o_77_sv2v_reg;
  assign el0_snoop_o[76] = el0_snoop_o_76_sv2v_reg;
  assign el0_snoop_o[75] = el0_snoop_o_75_sv2v_reg;
  assign el0_snoop_o[74] = el0_snoop_o_74_sv2v_reg;
  assign el0_snoop_o[73] = el0_snoop_o_73_sv2v_reg;
  assign el0_snoop_o[72] = el0_snoop_o_72_sv2v_reg;
  assign el0_snoop_o[71] = el0_snoop_o_71_sv2v_reg;
  assign el0_snoop_o[70] = el0_snoop_o_70_sv2v_reg;
  assign el0_snoop_o[69] = el0_snoop_o_69_sv2v_reg;
  assign el0_snoop_o[68] = el0_snoop_o_68_sv2v_reg;
  assign el0_snoop_o[67] = el0_snoop_o_67_sv2v_reg;
  assign el0_snoop_o[66] = el0_snoop_o_66_sv2v_reg;
  assign el0_snoop_o[65] = el0_snoop_o_65_sv2v_reg;
  assign el0_snoop_o[64] = el0_snoop_o_64_sv2v_reg;
  assign el0_snoop_o[63] = el0_snoop_o_63_sv2v_reg;
  assign el0_snoop_o[62] = el0_snoop_o_62_sv2v_reg;
  assign el0_snoop_o[61] = el0_snoop_o_61_sv2v_reg;
  assign el0_snoop_o[60] = el0_snoop_o_60_sv2v_reg;
  assign el0_snoop_o[59] = el0_snoop_o_59_sv2v_reg;
  assign el0_snoop_o[58] = el0_snoop_o_58_sv2v_reg;
  assign el0_snoop_o[57] = el0_snoop_o_57_sv2v_reg;
  assign el0_snoop_o[56] = el0_snoop_o_56_sv2v_reg;
  assign el0_snoop_o[55] = el0_snoop_o_55_sv2v_reg;
  assign el0_snoop_o[54] = el0_snoop_o_54_sv2v_reg;
  assign el0_snoop_o[53] = el0_snoop_o_53_sv2v_reg;
  assign el0_snoop_o[52] = el0_snoop_o_52_sv2v_reg;
  assign el0_snoop_o[51] = el0_snoop_o_51_sv2v_reg;
  assign el0_snoop_o[50] = el0_snoop_o_50_sv2v_reg;
  assign el0_snoop_o[49] = el0_snoop_o_49_sv2v_reg;
  assign el0_snoop_o[48] = el0_snoop_o_48_sv2v_reg;
  assign el0_snoop_o[47] = el0_snoop_o_47_sv2v_reg;
  assign el0_snoop_o[46] = el0_snoop_o_46_sv2v_reg;
  assign el0_snoop_o[45] = el0_snoop_o_45_sv2v_reg;
  assign el0_snoop_o[44] = el0_snoop_o_44_sv2v_reg;
  assign el0_snoop_o[43] = el0_snoop_o_43_sv2v_reg;
  assign el0_snoop_o[42] = el0_snoop_o_42_sv2v_reg;
  assign el0_snoop_o[41] = el0_snoop_o_41_sv2v_reg;
  assign el0_snoop_o[40] = el0_snoop_o_40_sv2v_reg;
  assign el0_snoop_o[39] = el0_snoop_o_39_sv2v_reg;
  assign el0_snoop_o[38] = el0_snoop_o_38_sv2v_reg;
  assign el0_snoop_o[37] = el0_snoop_o_37_sv2v_reg;
  assign el0_snoop_o[36] = el0_snoop_o_36_sv2v_reg;
  assign el0_snoop_o[35] = el0_snoop_o_35_sv2v_reg;
  assign el0_snoop_o[34] = el0_snoop_o_34_sv2v_reg;
  assign el0_snoop_o[33] = el0_snoop_o_33_sv2v_reg;
  assign el0_snoop_o[32] = el0_snoop_o_32_sv2v_reg;
  assign el0_snoop_o[31] = el0_snoop_o_31_sv2v_reg;
  assign el0_snoop_o[30] = el0_snoop_o_30_sv2v_reg;
  assign el0_snoop_o[29] = el0_snoop_o_29_sv2v_reg;
  assign el0_snoop_o[28] = el0_snoop_o_28_sv2v_reg;
  assign el0_snoop_o[27] = el0_snoop_o_27_sv2v_reg;
  assign el0_snoop_o[26] = el0_snoop_o_26_sv2v_reg;
  assign el0_snoop_o[25] = el0_snoop_o_25_sv2v_reg;
  assign el0_snoop_o[24] = el0_snoop_o_24_sv2v_reg;
  assign el0_snoop_o[23] = el0_snoop_o_23_sv2v_reg;
  assign el0_snoop_o[22] = el0_snoop_o_22_sv2v_reg;
  assign el0_snoop_o[21] = el0_snoop_o_21_sv2v_reg;
  assign el0_snoop_o[20] = el0_snoop_o_20_sv2v_reg;
  assign el0_snoop_o[19] = el0_snoop_o_19_sv2v_reg;
  assign el0_snoop_o[18] = el0_snoop_o_18_sv2v_reg;
  assign el0_snoop_o[17] = el0_snoop_o_17_sv2v_reg;
  assign el0_snoop_o[16] = el0_snoop_o_16_sv2v_reg;
  assign el0_snoop_o[15] = el0_snoop_o_15_sv2v_reg;
  assign el0_snoop_o[14] = el0_snoop_o_14_sv2v_reg;
  assign el0_snoop_o[13] = el0_snoop_o_13_sv2v_reg;
  assign el0_snoop_o[12] = el0_snoop_o_12_sv2v_reg;
  assign el0_snoop_o[11] = el0_snoop_o_11_sv2v_reg;
  assign el0_snoop_o[10] = el0_snoop_o_10_sv2v_reg;
  assign el0_snoop_o[9] = el0_snoop_o_9_sv2v_reg;
  assign el0_snoop_o[8] = el0_snoop_o_8_sv2v_reg;
  assign el0_snoop_o[7] = el0_snoop_o_7_sv2v_reg;
  assign el0_snoop_o[6] = el0_snoop_o_6_sv2v_reg;
  assign el0_snoop_o[5] = el0_snoop_o_5_sv2v_reg;
  assign el0_snoop_o[4] = el0_snoop_o_4_sv2v_reg;
  assign el0_snoop_o[3] = el0_snoop_o_3_sv2v_reg;
  assign el0_snoop_o[2] = el0_snoop_o_2_sv2v_reg;
  assign el0_snoop_o[1] = el0_snoop_o_1_sv2v_reg;
  assign el0_snoop_o[0] = el0_snoop_o_0_sv2v_reg;
  assign el1_snoop_o[179] = el1_snoop_o_179_sv2v_reg;
  assign el1_snoop_o[178] = el1_snoop_o_178_sv2v_reg;
  assign el1_snoop_o[177] = el1_snoop_o_177_sv2v_reg;
  assign el1_snoop_o[176] = el1_snoop_o_176_sv2v_reg;
  assign el1_snoop_o[175] = el1_snoop_o_175_sv2v_reg;
  assign el1_snoop_o[174] = el1_snoop_o_174_sv2v_reg;
  assign el1_snoop_o[173] = el1_snoop_o_173_sv2v_reg;
  assign el1_snoop_o[172] = el1_snoop_o_172_sv2v_reg;
  assign el1_snoop_o[171] = el1_snoop_o_171_sv2v_reg;
  assign el1_snoop_o[170] = el1_snoop_o_170_sv2v_reg;
  assign el1_snoop_o[169] = el1_snoop_o_169_sv2v_reg;
  assign el1_snoop_o[168] = el1_snoop_o_168_sv2v_reg;
  assign el1_snoop_o[167] = el1_snoop_o_167_sv2v_reg;
  assign el1_snoop_o[166] = el1_snoop_o_166_sv2v_reg;
  assign el1_snoop_o[165] = el1_snoop_o_165_sv2v_reg;
  assign el1_snoop_o[164] = el1_snoop_o_164_sv2v_reg;
  assign el1_snoop_o[163] = el1_snoop_o_163_sv2v_reg;
  assign el1_snoop_o[162] = el1_snoop_o_162_sv2v_reg;
  assign el1_snoop_o[161] = el1_snoop_o_161_sv2v_reg;
  assign el1_snoop_o[160] = el1_snoop_o_160_sv2v_reg;
  assign el1_snoop_o[159] = el1_snoop_o_159_sv2v_reg;
  assign el1_snoop_o[158] = el1_snoop_o_158_sv2v_reg;
  assign el1_snoop_o[157] = el1_snoop_o_157_sv2v_reg;
  assign el1_snoop_o[156] = el1_snoop_o_156_sv2v_reg;
  assign el1_snoop_o[155] = el1_snoop_o_155_sv2v_reg;
  assign el1_snoop_o[154] = el1_snoop_o_154_sv2v_reg;
  assign el1_snoop_o[153] = el1_snoop_o_153_sv2v_reg;
  assign el1_snoop_o[152] = el1_snoop_o_152_sv2v_reg;
  assign el1_snoop_o[151] = el1_snoop_o_151_sv2v_reg;
  assign el1_snoop_o[150] = el1_snoop_o_150_sv2v_reg;
  assign el1_snoop_o[149] = el1_snoop_o_149_sv2v_reg;
  assign el1_snoop_o[148] = el1_snoop_o_148_sv2v_reg;
  assign el1_snoop_o[147] = el1_snoop_o_147_sv2v_reg;
  assign el1_snoop_o[146] = el1_snoop_o_146_sv2v_reg;
  assign el1_snoop_o[145] = el1_snoop_o_145_sv2v_reg;
  assign el1_snoop_o[144] = el1_snoop_o_144_sv2v_reg;
  assign el1_snoop_o[143] = el1_snoop_o_143_sv2v_reg;
  assign el1_snoop_o[142] = el1_snoop_o_142_sv2v_reg;
  assign el1_snoop_o[141] = el1_snoop_o_141_sv2v_reg;
  assign el1_snoop_o[140] = el1_snoop_o_140_sv2v_reg;
  assign el1_snoop_o[139] = el1_snoop_o_139_sv2v_reg;
  assign el1_snoop_o[138] = el1_snoop_o_138_sv2v_reg;
  assign el1_snoop_o[137] = el1_snoop_o_137_sv2v_reg;
  assign el1_snoop_o[136] = el1_snoop_o_136_sv2v_reg;
  assign el1_snoop_o[135] = el1_snoop_o_135_sv2v_reg;
  assign el1_snoop_o[134] = el1_snoop_o_134_sv2v_reg;
  assign el1_snoop_o[133] = el1_snoop_o_133_sv2v_reg;
  assign el1_snoop_o[132] = el1_snoop_o_132_sv2v_reg;
  assign el1_snoop_o[131] = el1_snoop_o_131_sv2v_reg;
  assign el1_snoop_o[130] = el1_snoop_o_130_sv2v_reg;
  assign el1_snoop_o[129] = el1_snoop_o_129_sv2v_reg;
  assign el1_snoop_o[128] = el1_snoop_o_128_sv2v_reg;
  assign el1_snoop_o[127] = el1_snoop_o_127_sv2v_reg;
  assign el1_snoop_o[126] = el1_snoop_o_126_sv2v_reg;
  assign el1_snoop_o[125] = el1_snoop_o_125_sv2v_reg;
  assign el1_snoop_o[124] = el1_snoop_o_124_sv2v_reg;
  assign el1_snoop_o[123] = el1_snoop_o_123_sv2v_reg;
  assign el1_snoop_o[122] = el1_snoop_o_122_sv2v_reg;
  assign el1_snoop_o[121] = el1_snoop_o_121_sv2v_reg;
  assign el1_snoop_o[120] = el1_snoop_o_120_sv2v_reg;
  assign el1_snoop_o[119] = el1_snoop_o_119_sv2v_reg;
  assign el1_snoop_o[118] = el1_snoop_o_118_sv2v_reg;
  assign el1_snoop_o[117] = el1_snoop_o_117_sv2v_reg;
  assign el1_snoop_o[116] = el1_snoop_o_116_sv2v_reg;
  assign el1_snoop_o[115] = el1_snoop_o_115_sv2v_reg;
  assign el1_snoop_o[114] = el1_snoop_o_114_sv2v_reg;
  assign el1_snoop_o[113] = el1_snoop_o_113_sv2v_reg;
  assign el1_snoop_o[112] = el1_snoop_o_112_sv2v_reg;
  assign el1_snoop_o[111] = el1_snoop_o_111_sv2v_reg;
  assign el1_snoop_o[110] = el1_snoop_o_110_sv2v_reg;
  assign el1_snoop_o[109] = el1_snoop_o_109_sv2v_reg;
  assign el1_snoop_o[108] = el1_snoop_o_108_sv2v_reg;
  assign el1_snoop_o[107] = el1_snoop_o_107_sv2v_reg;
  assign el1_snoop_o[106] = el1_snoop_o_106_sv2v_reg;
  assign el1_snoop_o[105] = el1_snoop_o_105_sv2v_reg;
  assign el1_snoop_o[104] = el1_snoop_o_104_sv2v_reg;
  assign el1_snoop_o[103] = el1_snoop_o_103_sv2v_reg;
  assign el1_snoop_o[102] = el1_snoop_o_102_sv2v_reg;
  assign el1_snoop_o[101] = el1_snoop_o_101_sv2v_reg;
  assign el1_snoop_o[100] = el1_snoop_o_100_sv2v_reg;
  assign el1_snoop_o[99] = el1_snoop_o_99_sv2v_reg;
  assign el1_snoop_o[98] = el1_snoop_o_98_sv2v_reg;
  assign el1_snoop_o[97] = el1_snoop_o_97_sv2v_reg;
  assign el1_snoop_o[96] = el1_snoop_o_96_sv2v_reg;
  assign el1_snoop_o[95] = el1_snoop_o_95_sv2v_reg;
  assign el1_snoop_o[94] = el1_snoop_o_94_sv2v_reg;
  assign el1_snoop_o[93] = el1_snoop_o_93_sv2v_reg;
  assign el1_snoop_o[92] = el1_snoop_o_92_sv2v_reg;
  assign el1_snoop_o[91] = el1_snoop_o_91_sv2v_reg;
  assign el1_snoop_o[90] = el1_snoop_o_90_sv2v_reg;
  assign el1_snoop_o[89] = el1_snoop_o_89_sv2v_reg;
  assign el1_snoop_o[88] = el1_snoop_o_88_sv2v_reg;
  assign el1_snoop_o[87] = el1_snoop_o_87_sv2v_reg;
  assign el1_snoop_o[86] = el1_snoop_o_86_sv2v_reg;
  assign el1_snoop_o[85] = el1_snoop_o_85_sv2v_reg;
  assign el1_snoop_o[84] = el1_snoop_o_84_sv2v_reg;
  assign el1_snoop_o[83] = el1_snoop_o_83_sv2v_reg;
  assign el1_snoop_o[82] = el1_snoop_o_82_sv2v_reg;
  assign el1_snoop_o[81] = el1_snoop_o_81_sv2v_reg;
  assign el1_snoop_o[80] = el1_snoop_o_80_sv2v_reg;
  assign el1_snoop_o[79] = el1_snoop_o_79_sv2v_reg;
  assign el1_snoop_o[78] = el1_snoop_o_78_sv2v_reg;
  assign el1_snoop_o[77] = el1_snoop_o_77_sv2v_reg;
  assign el1_snoop_o[76] = el1_snoop_o_76_sv2v_reg;
  assign el1_snoop_o[75] = el1_snoop_o_75_sv2v_reg;
  assign el1_snoop_o[74] = el1_snoop_o_74_sv2v_reg;
  assign el1_snoop_o[73] = el1_snoop_o_73_sv2v_reg;
  assign el1_snoop_o[72] = el1_snoop_o_72_sv2v_reg;
  assign el1_snoop_o[71] = el1_snoop_o_71_sv2v_reg;
  assign el1_snoop_o[70] = el1_snoop_o_70_sv2v_reg;
  assign el1_snoop_o[69] = el1_snoop_o_69_sv2v_reg;
  assign el1_snoop_o[68] = el1_snoop_o_68_sv2v_reg;
  assign el1_snoop_o[67] = el1_snoop_o_67_sv2v_reg;
  assign el1_snoop_o[66] = el1_snoop_o_66_sv2v_reg;
  assign el1_snoop_o[65] = el1_snoop_o_65_sv2v_reg;
  assign el1_snoop_o[64] = el1_snoop_o_64_sv2v_reg;
  assign el1_snoop_o[63] = el1_snoop_o_63_sv2v_reg;
  assign el1_snoop_o[62] = el1_snoop_o_62_sv2v_reg;
  assign el1_snoop_o[61] = el1_snoop_o_61_sv2v_reg;
  assign el1_snoop_o[60] = el1_snoop_o_60_sv2v_reg;
  assign el1_snoop_o[59] = el1_snoop_o_59_sv2v_reg;
  assign el1_snoop_o[58] = el1_snoop_o_58_sv2v_reg;
  assign el1_snoop_o[57] = el1_snoop_o_57_sv2v_reg;
  assign el1_snoop_o[56] = el1_snoop_o_56_sv2v_reg;
  assign el1_snoop_o[55] = el1_snoop_o_55_sv2v_reg;
  assign el1_snoop_o[54] = el1_snoop_o_54_sv2v_reg;
  assign el1_snoop_o[53] = el1_snoop_o_53_sv2v_reg;
  assign el1_snoop_o[52] = el1_snoop_o_52_sv2v_reg;
  assign el1_snoop_o[51] = el1_snoop_o_51_sv2v_reg;
  assign el1_snoop_o[50] = el1_snoop_o_50_sv2v_reg;
  assign el1_snoop_o[49] = el1_snoop_o_49_sv2v_reg;
  assign el1_snoop_o[48] = el1_snoop_o_48_sv2v_reg;
  assign el1_snoop_o[47] = el1_snoop_o_47_sv2v_reg;
  assign el1_snoop_o[46] = el1_snoop_o_46_sv2v_reg;
  assign el1_snoop_o[45] = el1_snoop_o_45_sv2v_reg;
  assign el1_snoop_o[44] = el1_snoop_o_44_sv2v_reg;
  assign el1_snoop_o[43] = el1_snoop_o_43_sv2v_reg;
  assign el1_snoop_o[42] = el1_snoop_o_42_sv2v_reg;
  assign el1_snoop_o[41] = el1_snoop_o_41_sv2v_reg;
  assign el1_snoop_o[40] = el1_snoop_o_40_sv2v_reg;
  assign el1_snoop_o[39] = el1_snoop_o_39_sv2v_reg;
  assign el1_snoop_o[38] = el1_snoop_o_38_sv2v_reg;
  assign el1_snoop_o[37] = el1_snoop_o_37_sv2v_reg;
  assign el1_snoop_o[36] = el1_snoop_o_36_sv2v_reg;
  assign el1_snoop_o[35] = el1_snoop_o_35_sv2v_reg;
  assign el1_snoop_o[34] = el1_snoop_o_34_sv2v_reg;
  assign el1_snoop_o[33] = el1_snoop_o_33_sv2v_reg;
  assign el1_snoop_o[32] = el1_snoop_o_32_sv2v_reg;
  assign el1_snoop_o[31] = el1_snoop_o_31_sv2v_reg;
  assign el1_snoop_o[30] = el1_snoop_o_30_sv2v_reg;
  assign el1_snoop_o[29] = el1_snoop_o_29_sv2v_reg;
  assign el1_snoop_o[28] = el1_snoop_o_28_sv2v_reg;
  assign el1_snoop_o[27] = el1_snoop_o_27_sv2v_reg;
  assign el1_snoop_o[26] = el1_snoop_o_26_sv2v_reg;
  assign el1_snoop_o[25] = el1_snoop_o_25_sv2v_reg;
  assign el1_snoop_o[24] = el1_snoop_o_24_sv2v_reg;
  assign el1_snoop_o[23] = el1_snoop_o_23_sv2v_reg;
  assign el1_snoop_o[22] = el1_snoop_o_22_sv2v_reg;
  assign el1_snoop_o[21] = el1_snoop_o_21_sv2v_reg;
  assign el1_snoop_o[20] = el1_snoop_o_20_sv2v_reg;
  assign el1_snoop_o[19] = el1_snoop_o_19_sv2v_reg;
  assign el1_snoop_o[18] = el1_snoop_o_18_sv2v_reg;
  assign el1_snoop_o[17] = el1_snoop_o_17_sv2v_reg;
  assign el1_snoop_o[16] = el1_snoop_o_16_sv2v_reg;
  assign el1_snoop_o[15] = el1_snoop_o_15_sv2v_reg;
  assign el1_snoop_o[14] = el1_snoop_o_14_sv2v_reg;
  assign el1_snoop_o[13] = el1_snoop_o_13_sv2v_reg;
  assign el1_snoop_o[12] = el1_snoop_o_12_sv2v_reg;
  assign el1_snoop_o[11] = el1_snoop_o_11_sv2v_reg;
  assign el1_snoop_o[10] = el1_snoop_o_10_sv2v_reg;
  assign el1_snoop_o[9] = el1_snoop_o_9_sv2v_reg;
  assign el1_snoop_o[8] = el1_snoop_o_8_sv2v_reg;
  assign el1_snoop_o[7] = el1_snoop_o_7_sv2v_reg;
  assign el1_snoop_o[6] = el1_snoop_o_6_sv2v_reg;
  assign el1_snoop_o[5] = el1_snoop_o_5_sv2v_reg;
  assign el1_snoop_o[4] = el1_snoop_o_4_sv2v_reg;
  assign el1_snoop_o[3] = el1_snoop_o_3_sv2v_reg;
  assign el1_snoop_o[2] = el1_snoop_o_2_sv2v_reg;
  assign el1_snoop_o[1] = el1_snoop_o_1_sv2v_reg;
  assign el1_snoop_o[0] = el1_snoop_o_0_sv2v_reg;
  assign N10 = N8 & N9;
  assign N11 = num_els_r[1] | N9;
  assign N13 = N8 | num_els_r[0];
  assign N15 = num_els_r[1] & num_els_r[0];
  assign { N20, N19 } = num_els_r + v_i;
  assign { N23, N22 } = { N20, N19 } - N21;
  assign v_o = (N0)? v_i : 
               (N1)? 1'b1 : 
               (N2)? 1'b1 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = N10;
  assign N1 = N12;
  assign N2 = N14;
  assign N3 = N15;
  assign empty_o = (N0)? 1'b1 : 
                   (N1)? 1'b0 : 
                   (N2)? 1'b0 : 
                   (N3)? 1'b0 : 1'b0;
  assign full_o = (N0)? 1'b0 : 
                  (N1)? 1'b0 : 
                  (N2)? 1'b1 : 
                  (N3)? 1'b0 : 1'b0;
  assign el0_valid_o = (N0)? 1'b0 : 
                       (N1)? 1'b0 : 
                       (N2)? 1'b1 : 
                       (N3)? 1'b0 : 1'b0;
  assign el1_valid_o = (N0)? 1'b0 : 
                       (N1)? 1'b1 : 
                       (N2)? 1'b1 : 
                       (N3)? 1'b0 : 1'b0;
  assign el0_enable = (N0)? 1'b0 : 
                      (N1)? N16 : 
                      (N2)? N17 : 
                      (N3)? 1'b0 : 1'b0;
  assign el1_enable = (N0)? N16 : 
                      (N1)? N17 : 
                      (N2)? yumi_i : 
                      (N3)? 1'b0 : 1'b0;
  assign mux0_sel = (N0)? 1'b0 : 
                    (N1)? 1'b0 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b0 : 1'b0;
  assign mux1_sel = (N0)? 1'b0 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b0 : 1'b0;
  assign { N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25 } = (N4)? el0_snoop_o : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           (N5)? data_i : 1'b0;
  assign N4 = mux0_sel;
  assign N5 = N24;
  assign data_o = (N6)? el1_snoop_o : 
                  (N7)? data_i : 1'b0;
  assign N6 = mux1_sel;
  assign N7 = N205;
  assign N8 = ~num_els_r[1];
  assign N9 = ~num_els_r[0];
  assign N12 = ~N11;
  assign N14 = ~N13;
  assign N16 = v_i & N206;
  assign N206 = ~yumi_i;
  assign N17 = v_i & yumi_i;
  assign N18 = ~reset_i;
  assign N21 = v_o & yumi_i;
  assign N24 = ~mux0_sel;
  assign N205 = ~mux1_sel;

  always @(posedge clk_i) begin
    if(reset_i) begin
      num_els_r_1_sv2v_reg <= 1'b0;
      num_els_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      num_els_r_1_sv2v_reg <= N23;
      num_els_r_0_sv2v_reg <= N22;
    end 
    if(el0_enable) begin
      el0_snoop_o_179_sv2v_reg <= data_i[179];
      el0_snoop_o_178_sv2v_reg <= data_i[178];
      el0_snoop_o_177_sv2v_reg <= data_i[177];
      el0_snoop_o_176_sv2v_reg <= data_i[176];
      el0_snoop_o_175_sv2v_reg <= data_i[175];
      el0_snoop_o_174_sv2v_reg <= data_i[174];
      el0_snoop_o_173_sv2v_reg <= data_i[173];
      el0_snoop_o_172_sv2v_reg <= data_i[172];
      el0_snoop_o_171_sv2v_reg <= data_i[171];
      el0_snoop_o_170_sv2v_reg <= data_i[170];
      el0_snoop_o_169_sv2v_reg <= data_i[169];
      el0_snoop_o_168_sv2v_reg <= data_i[168];
      el0_snoop_o_167_sv2v_reg <= data_i[167];
      el0_snoop_o_166_sv2v_reg <= data_i[166];
      el0_snoop_o_165_sv2v_reg <= data_i[165];
      el0_snoop_o_164_sv2v_reg <= data_i[164];
      el0_snoop_o_163_sv2v_reg <= data_i[163];
      el0_snoop_o_162_sv2v_reg <= data_i[162];
      el0_snoop_o_161_sv2v_reg <= data_i[161];
      el0_snoop_o_160_sv2v_reg <= data_i[160];
      el0_snoop_o_159_sv2v_reg <= data_i[159];
      el0_snoop_o_158_sv2v_reg <= data_i[158];
      el0_snoop_o_157_sv2v_reg <= data_i[157];
      el0_snoop_o_156_sv2v_reg <= data_i[156];
      el0_snoop_o_155_sv2v_reg <= data_i[155];
      el0_snoop_o_154_sv2v_reg <= data_i[154];
      el0_snoop_o_153_sv2v_reg <= data_i[153];
      el0_snoop_o_152_sv2v_reg <= data_i[152];
      el0_snoop_o_151_sv2v_reg <= data_i[151];
      el0_snoop_o_150_sv2v_reg <= data_i[150];
      el0_snoop_o_149_sv2v_reg <= data_i[149];
      el0_snoop_o_148_sv2v_reg <= data_i[148];
      el0_snoop_o_147_sv2v_reg <= data_i[147];
      el0_snoop_o_146_sv2v_reg <= data_i[146];
      el0_snoop_o_145_sv2v_reg <= data_i[145];
      el0_snoop_o_144_sv2v_reg <= data_i[144];
      el0_snoop_o_143_sv2v_reg <= data_i[143];
      el0_snoop_o_142_sv2v_reg <= data_i[142];
      el0_snoop_o_141_sv2v_reg <= data_i[141];
      el0_snoop_o_140_sv2v_reg <= data_i[140];
      el0_snoop_o_139_sv2v_reg <= data_i[139];
      el0_snoop_o_138_sv2v_reg <= data_i[138];
      el0_snoop_o_137_sv2v_reg <= data_i[137];
      el0_snoop_o_136_sv2v_reg <= data_i[136];
      el0_snoop_o_135_sv2v_reg <= data_i[135];
      el0_snoop_o_134_sv2v_reg <= data_i[134];
      el0_snoop_o_133_sv2v_reg <= data_i[133];
      el0_snoop_o_132_sv2v_reg <= data_i[132];
      el0_snoop_o_131_sv2v_reg <= data_i[131];
      el0_snoop_o_130_sv2v_reg <= data_i[130];
      el0_snoop_o_129_sv2v_reg <= data_i[129];
      el0_snoop_o_128_sv2v_reg <= data_i[128];
      el0_snoop_o_127_sv2v_reg <= data_i[127];
      el0_snoop_o_126_sv2v_reg <= data_i[126];
      el0_snoop_o_125_sv2v_reg <= data_i[125];
      el0_snoop_o_124_sv2v_reg <= data_i[124];
      el0_snoop_o_123_sv2v_reg <= data_i[123];
      el0_snoop_o_122_sv2v_reg <= data_i[122];
      el0_snoop_o_121_sv2v_reg <= data_i[121];
      el0_snoop_o_120_sv2v_reg <= data_i[120];
      el0_snoop_o_119_sv2v_reg <= data_i[119];
      el0_snoop_o_118_sv2v_reg <= data_i[118];
      el0_snoop_o_117_sv2v_reg <= data_i[117];
      el0_snoop_o_116_sv2v_reg <= data_i[116];
      el0_snoop_o_115_sv2v_reg <= data_i[115];
      el0_snoop_o_114_sv2v_reg <= data_i[114];
      el0_snoop_o_113_sv2v_reg <= data_i[113];
      el0_snoop_o_112_sv2v_reg <= data_i[112];
      el0_snoop_o_111_sv2v_reg <= data_i[111];
      el0_snoop_o_110_sv2v_reg <= data_i[110];
      el0_snoop_o_109_sv2v_reg <= data_i[109];
      el0_snoop_o_108_sv2v_reg <= data_i[108];
      el0_snoop_o_107_sv2v_reg <= data_i[107];
      el0_snoop_o_106_sv2v_reg <= data_i[106];
      el0_snoop_o_105_sv2v_reg <= data_i[105];
      el0_snoop_o_104_sv2v_reg <= data_i[104];
      el0_snoop_o_103_sv2v_reg <= data_i[103];
      el0_snoop_o_102_sv2v_reg <= data_i[102];
      el0_snoop_o_101_sv2v_reg <= data_i[101];
      el0_snoop_o_100_sv2v_reg <= data_i[100];
      el0_snoop_o_99_sv2v_reg <= data_i[99];
      el0_snoop_o_98_sv2v_reg <= data_i[98];
      el0_snoop_o_97_sv2v_reg <= data_i[97];
      el0_snoop_o_96_sv2v_reg <= data_i[96];
      el0_snoop_o_95_sv2v_reg <= data_i[95];
      el0_snoop_o_94_sv2v_reg <= data_i[94];
      el0_snoop_o_93_sv2v_reg <= data_i[93];
      el0_snoop_o_92_sv2v_reg <= data_i[92];
      el0_snoop_o_91_sv2v_reg <= data_i[91];
      el0_snoop_o_90_sv2v_reg <= data_i[90];
      el0_snoop_o_89_sv2v_reg <= data_i[89];
      el0_snoop_o_88_sv2v_reg <= data_i[88];
      el0_snoop_o_87_sv2v_reg <= data_i[87];
      el0_snoop_o_86_sv2v_reg <= data_i[86];
      el0_snoop_o_85_sv2v_reg <= data_i[85];
      el0_snoop_o_84_sv2v_reg <= data_i[84];
      el0_snoop_o_83_sv2v_reg <= data_i[83];
      el0_snoop_o_82_sv2v_reg <= data_i[82];
      el0_snoop_o_81_sv2v_reg <= data_i[81];
      el0_snoop_o_80_sv2v_reg <= data_i[80];
      el0_snoop_o_79_sv2v_reg <= data_i[79];
      el0_snoop_o_78_sv2v_reg <= data_i[78];
      el0_snoop_o_77_sv2v_reg <= data_i[77];
      el0_snoop_o_76_sv2v_reg <= data_i[76];
      el0_snoop_o_75_sv2v_reg <= data_i[75];
      el0_snoop_o_74_sv2v_reg <= data_i[74];
      el0_snoop_o_73_sv2v_reg <= data_i[73];
      el0_snoop_o_72_sv2v_reg <= data_i[72];
      el0_snoop_o_71_sv2v_reg <= data_i[71];
      el0_snoop_o_70_sv2v_reg <= data_i[70];
      el0_snoop_o_69_sv2v_reg <= data_i[69];
      el0_snoop_o_68_sv2v_reg <= data_i[68];
      el0_snoop_o_67_sv2v_reg <= data_i[67];
      el0_snoop_o_66_sv2v_reg <= data_i[66];
      el0_snoop_o_65_sv2v_reg <= data_i[65];
      el0_snoop_o_64_sv2v_reg <= data_i[64];
      el0_snoop_o_63_sv2v_reg <= data_i[63];
      el0_snoop_o_62_sv2v_reg <= data_i[62];
      el0_snoop_o_61_sv2v_reg <= data_i[61];
      el0_snoop_o_60_sv2v_reg <= data_i[60];
      el0_snoop_o_59_sv2v_reg <= data_i[59];
      el0_snoop_o_58_sv2v_reg <= data_i[58];
      el0_snoop_o_57_sv2v_reg <= data_i[57];
      el0_snoop_o_56_sv2v_reg <= data_i[56];
      el0_snoop_o_55_sv2v_reg <= data_i[55];
      el0_snoop_o_54_sv2v_reg <= data_i[54];
      el0_snoop_o_53_sv2v_reg <= data_i[53];
      el0_snoop_o_52_sv2v_reg <= data_i[52];
      el0_snoop_o_51_sv2v_reg <= data_i[51];
      el0_snoop_o_50_sv2v_reg <= data_i[50];
      el0_snoop_o_49_sv2v_reg <= data_i[49];
      el0_snoop_o_48_sv2v_reg <= data_i[48];
      el0_snoop_o_47_sv2v_reg <= data_i[47];
      el0_snoop_o_46_sv2v_reg <= data_i[46];
      el0_snoop_o_45_sv2v_reg <= data_i[45];
      el0_snoop_o_44_sv2v_reg <= data_i[44];
      el0_snoop_o_43_sv2v_reg <= data_i[43];
      el0_snoop_o_42_sv2v_reg <= data_i[42];
      el0_snoop_o_41_sv2v_reg <= data_i[41];
      el0_snoop_o_40_sv2v_reg <= data_i[40];
      el0_snoop_o_39_sv2v_reg <= data_i[39];
      el0_snoop_o_38_sv2v_reg <= data_i[38];
      el0_snoop_o_37_sv2v_reg <= data_i[37];
      el0_snoop_o_36_sv2v_reg <= data_i[36];
      el0_snoop_o_35_sv2v_reg <= data_i[35];
      el0_snoop_o_34_sv2v_reg <= data_i[34];
      el0_snoop_o_33_sv2v_reg <= data_i[33];
      el0_snoop_o_32_sv2v_reg <= data_i[32];
      el0_snoop_o_31_sv2v_reg <= data_i[31];
      el0_snoop_o_30_sv2v_reg <= data_i[30];
      el0_snoop_o_29_sv2v_reg <= data_i[29];
      el0_snoop_o_28_sv2v_reg <= data_i[28];
      el0_snoop_o_27_sv2v_reg <= data_i[27];
      el0_snoop_o_26_sv2v_reg <= data_i[26];
      el0_snoop_o_25_sv2v_reg <= data_i[25];
      el0_snoop_o_24_sv2v_reg <= data_i[24];
      el0_snoop_o_23_sv2v_reg <= data_i[23];
      el0_snoop_o_22_sv2v_reg <= data_i[22];
      el0_snoop_o_21_sv2v_reg <= data_i[21];
      el0_snoop_o_20_sv2v_reg <= data_i[20];
      el0_snoop_o_19_sv2v_reg <= data_i[19];
      el0_snoop_o_18_sv2v_reg <= data_i[18];
      el0_snoop_o_17_sv2v_reg <= data_i[17];
      el0_snoop_o_16_sv2v_reg <= data_i[16];
      el0_snoop_o_15_sv2v_reg <= data_i[15];
      el0_snoop_o_14_sv2v_reg <= data_i[14];
      el0_snoop_o_13_sv2v_reg <= data_i[13];
      el0_snoop_o_12_sv2v_reg <= data_i[12];
      el0_snoop_o_11_sv2v_reg <= data_i[11];
      el0_snoop_o_10_sv2v_reg <= data_i[10];
      el0_snoop_o_9_sv2v_reg <= data_i[9];
      el0_snoop_o_8_sv2v_reg <= data_i[8];
      el0_snoop_o_7_sv2v_reg <= data_i[7];
      el0_snoop_o_6_sv2v_reg <= data_i[6];
      el0_snoop_o_5_sv2v_reg <= data_i[5];
      el0_snoop_o_4_sv2v_reg <= data_i[4];
      el0_snoop_o_3_sv2v_reg <= data_i[3];
      el0_snoop_o_2_sv2v_reg <= data_i[2];
      el0_snoop_o_1_sv2v_reg <= data_i[1];
      el0_snoop_o_0_sv2v_reg <= data_i[0];
    end 
    if(el1_enable) begin
      el1_snoop_o_179_sv2v_reg <= N204;
      el1_snoop_o_178_sv2v_reg <= N203;
      el1_snoop_o_177_sv2v_reg <= N202;
      el1_snoop_o_176_sv2v_reg <= N201;
      el1_snoop_o_175_sv2v_reg <= N200;
      el1_snoop_o_174_sv2v_reg <= N199;
      el1_snoop_o_173_sv2v_reg <= N198;
      el1_snoop_o_172_sv2v_reg <= N197;
      el1_snoop_o_171_sv2v_reg <= N196;
      el1_snoop_o_170_sv2v_reg <= N195;
      el1_snoop_o_169_sv2v_reg <= N194;
      el1_snoop_o_168_sv2v_reg <= N193;
      el1_snoop_o_167_sv2v_reg <= N192;
      el1_snoop_o_166_sv2v_reg <= N191;
      el1_snoop_o_165_sv2v_reg <= N190;
      el1_snoop_o_164_sv2v_reg <= N189;
      el1_snoop_o_163_sv2v_reg <= N188;
      el1_snoop_o_162_sv2v_reg <= N187;
      el1_snoop_o_161_sv2v_reg <= N186;
      el1_snoop_o_160_sv2v_reg <= N185;
      el1_snoop_o_159_sv2v_reg <= N184;
      el1_snoop_o_158_sv2v_reg <= N183;
      el1_snoop_o_157_sv2v_reg <= N182;
      el1_snoop_o_156_sv2v_reg <= N181;
      el1_snoop_o_155_sv2v_reg <= N180;
      el1_snoop_o_154_sv2v_reg <= N179;
      el1_snoop_o_153_sv2v_reg <= N178;
      el1_snoop_o_152_sv2v_reg <= N177;
      el1_snoop_o_151_sv2v_reg <= N176;
      el1_snoop_o_150_sv2v_reg <= N175;
      el1_snoop_o_149_sv2v_reg <= N174;
      el1_snoop_o_148_sv2v_reg <= N173;
      el1_snoop_o_147_sv2v_reg <= N172;
      el1_snoop_o_146_sv2v_reg <= N171;
      el1_snoop_o_145_sv2v_reg <= N170;
      el1_snoop_o_144_sv2v_reg <= N169;
      el1_snoop_o_143_sv2v_reg <= N168;
      el1_snoop_o_142_sv2v_reg <= N167;
      el1_snoop_o_141_sv2v_reg <= N166;
      el1_snoop_o_140_sv2v_reg <= N165;
      el1_snoop_o_139_sv2v_reg <= N164;
      el1_snoop_o_138_sv2v_reg <= N163;
      el1_snoop_o_137_sv2v_reg <= N162;
      el1_snoop_o_136_sv2v_reg <= N161;
      el1_snoop_o_135_sv2v_reg <= N160;
      el1_snoop_o_134_sv2v_reg <= N159;
      el1_snoop_o_133_sv2v_reg <= N158;
      el1_snoop_o_132_sv2v_reg <= N157;
      el1_snoop_o_131_sv2v_reg <= N156;
      el1_snoop_o_130_sv2v_reg <= N155;
      el1_snoop_o_129_sv2v_reg <= N154;
      el1_snoop_o_128_sv2v_reg <= N153;
      el1_snoop_o_127_sv2v_reg <= N152;
      el1_snoop_o_126_sv2v_reg <= N151;
      el1_snoop_o_125_sv2v_reg <= N150;
      el1_snoop_o_124_sv2v_reg <= N149;
      el1_snoop_o_123_sv2v_reg <= N148;
      el1_snoop_o_122_sv2v_reg <= N147;
      el1_snoop_o_121_sv2v_reg <= N146;
      el1_snoop_o_120_sv2v_reg <= N145;
      el1_snoop_o_119_sv2v_reg <= N144;
      el1_snoop_o_118_sv2v_reg <= N143;
      el1_snoop_o_117_sv2v_reg <= N142;
      el1_snoop_o_116_sv2v_reg <= N141;
      el1_snoop_o_115_sv2v_reg <= N140;
      el1_snoop_o_114_sv2v_reg <= N139;
      el1_snoop_o_113_sv2v_reg <= N138;
      el1_snoop_o_112_sv2v_reg <= N137;
      el1_snoop_o_111_sv2v_reg <= N136;
      el1_snoop_o_110_sv2v_reg <= N135;
      el1_snoop_o_109_sv2v_reg <= N134;
      el1_snoop_o_108_sv2v_reg <= N133;
      el1_snoop_o_107_sv2v_reg <= N132;
      el1_snoop_o_106_sv2v_reg <= N131;
      el1_snoop_o_105_sv2v_reg <= N130;
      el1_snoop_o_104_sv2v_reg <= N129;
      el1_snoop_o_103_sv2v_reg <= N128;
      el1_snoop_o_102_sv2v_reg <= N127;
      el1_snoop_o_101_sv2v_reg <= N126;
      el1_snoop_o_100_sv2v_reg <= N125;
      el1_snoop_o_99_sv2v_reg <= N124;
      el1_snoop_o_98_sv2v_reg <= N123;
      el1_snoop_o_97_sv2v_reg <= N122;
      el1_snoop_o_96_sv2v_reg <= N121;
      el1_snoop_o_95_sv2v_reg <= N120;
      el1_snoop_o_94_sv2v_reg <= N119;
      el1_snoop_o_93_sv2v_reg <= N118;
      el1_snoop_o_92_sv2v_reg <= N117;
      el1_snoop_o_91_sv2v_reg <= N116;
      el1_snoop_o_90_sv2v_reg <= N115;
      el1_snoop_o_89_sv2v_reg <= N114;
      el1_snoop_o_88_sv2v_reg <= N113;
      el1_snoop_o_87_sv2v_reg <= N112;
      el1_snoop_o_86_sv2v_reg <= N111;
      el1_snoop_o_85_sv2v_reg <= N110;
      el1_snoop_o_84_sv2v_reg <= N109;
      el1_snoop_o_83_sv2v_reg <= N108;
      el1_snoop_o_82_sv2v_reg <= N107;
      el1_snoop_o_81_sv2v_reg <= N106;
      el1_snoop_o_80_sv2v_reg <= N105;
      el1_snoop_o_79_sv2v_reg <= N104;
      el1_snoop_o_78_sv2v_reg <= N103;
      el1_snoop_o_77_sv2v_reg <= N102;
      el1_snoop_o_76_sv2v_reg <= N101;
      el1_snoop_o_75_sv2v_reg <= N100;
      el1_snoop_o_74_sv2v_reg <= N99;
      el1_snoop_o_73_sv2v_reg <= N98;
      el1_snoop_o_72_sv2v_reg <= N97;
      el1_snoop_o_71_sv2v_reg <= N96;
      el1_snoop_o_70_sv2v_reg <= N95;
      el1_snoop_o_69_sv2v_reg <= N94;
      el1_snoop_o_68_sv2v_reg <= N93;
      el1_snoop_o_67_sv2v_reg <= N92;
      el1_snoop_o_66_sv2v_reg <= N91;
      el1_snoop_o_65_sv2v_reg <= N90;
      el1_snoop_o_64_sv2v_reg <= N89;
      el1_snoop_o_63_sv2v_reg <= N88;
      el1_snoop_o_62_sv2v_reg <= N87;
      el1_snoop_o_61_sv2v_reg <= N86;
      el1_snoop_o_60_sv2v_reg <= N85;
      el1_snoop_o_59_sv2v_reg <= N84;
      el1_snoop_o_58_sv2v_reg <= N83;
      el1_snoop_o_57_sv2v_reg <= N82;
      el1_snoop_o_56_sv2v_reg <= N81;
      el1_snoop_o_55_sv2v_reg <= N80;
      el1_snoop_o_54_sv2v_reg <= N79;
      el1_snoop_o_53_sv2v_reg <= N78;
      el1_snoop_o_52_sv2v_reg <= N77;
      el1_snoop_o_51_sv2v_reg <= N76;
      el1_snoop_o_50_sv2v_reg <= N75;
      el1_snoop_o_49_sv2v_reg <= N74;
      el1_snoop_o_48_sv2v_reg <= N73;
      el1_snoop_o_47_sv2v_reg <= N72;
      el1_snoop_o_46_sv2v_reg <= N71;
      el1_snoop_o_45_sv2v_reg <= N70;
      el1_snoop_o_44_sv2v_reg <= N69;
      el1_snoop_o_43_sv2v_reg <= N68;
      el1_snoop_o_42_sv2v_reg <= N67;
      el1_snoop_o_41_sv2v_reg <= N66;
      el1_snoop_o_40_sv2v_reg <= N65;
      el1_snoop_o_39_sv2v_reg <= N64;
      el1_snoop_o_38_sv2v_reg <= N63;
      el1_snoop_o_37_sv2v_reg <= N62;
      el1_snoop_o_36_sv2v_reg <= N61;
      el1_snoop_o_35_sv2v_reg <= N60;
      el1_snoop_o_34_sv2v_reg <= N59;
      el1_snoop_o_33_sv2v_reg <= N58;
      el1_snoop_o_32_sv2v_reg <= N57;
      el1_snoop_o_31_sv2v_reg <= N56;
      el1_snoop_o_30_sv2v_reg <= N55;
      el1_snoop_o_29_sv2v_reg <= N54;
      el1_snoop_o_28_sv2v_reg <= N53;
      el1_snoop_o_27_sv2v_reg <= N52;
      el1_snoop_o_26_sv2v_reg <= N51;
      el1_snoop_o_25_sv2v_reg <= N50;
      el1_snoop_o_24_sv2v_reg <= N49;
      el1_snoop_o_23_sv2v_reg <= N48;
      el1_snoop_o_22_sv2v_reg <= N47;
      el1_snoop_o_21_sv2v_reg <= N46;
      el1_snoop_o_20_sv2v_reg <= N45;
      el1_snoop_o_19_sv2v_reg <= N44;
      el1_snoop_o_18_sv2v_reg <= N43;
      el1_snoop_o_17_sv2v_reg <= N42;
      el1_snoop_o_16_sv2v_reg <= N41;
      el1_snoop_o_15_sv2v_reg <= N40;
      el1_snoop_o_14_sv2v_reg <= N39;
      el1_snoop_o_13_sv2v_reg <= N38;
      el1_snoop_o_12_sv2v_reg <= N37;
      el1_snoop_o_11_sv2v_reg <= N36;
      el1_snoop_o_10_sv2v_reg <= N35;
      el1_snoop_o_9_sv2v_reg <= N34;
      el1_snoop_o_8_sv2v_reg <= N33;
      el1_snoop_o_7_sv2v_reg <= N32;
      el1_snoop_o_6_sv2v_reg <= N31;
      el1_snoop_o_5_sv2v_reg <= N30;
      el1_snoop_o_4_sv2v_reg <= N29;
      el1_snoop_o_3_sv2v_reg <= N28;
      el1_snoop_o_2_sv2v_reg <= N27;
      el1_snoop_o_1_sv2v_reg <= N26;
      el1_snoop_o_0_sv2v_reg <= N25;
    end 
  end


endmodule



module bsg_mux_segmented_00000010_8
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [127:0] data0_i;
  input [127:0] data1_i;
  input [15:0] sel_i;
  output [127:0] data_o;
  wire [127:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31;
  assign data_o[7:0] = (N0)? data1_i[7:0] : 
                       (N16)? data0_i[7:0] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[15:8] = (N1)? data1_i[15:8] : 
                        (N17)? data0_i[15:8] : 1'b0;
  assign N1 = sel_i[1];
  assign data_o[23:16] = (N2)? data1_i[23:16] : 
                         (N18)? data0_i[23:16] : 1'b0;
  assign N2 = sel_i[2];
  assign data_o[31:24] = (N3)? data1_i[31:24] : 
                         (N19)? data0_i[31:24] : 1'b0;
  assign N3 = sel_i[3];
  assign data_o[39:32] = (N4)? data1_i[39:32] : 
                         (N20)? data0_i[39:32] : 1'b0;
  assign N4 = sel_i[4];
  assign data_o[47:40] = (N5)? data1_i[47:40] : 
                         (N21)? data0_i[47:40] : 1'b0;
  assign N5 = sel_i[5];
  assign data_o[55:48] = (N6)? data1_i[55:48] : 
                         (N22)? data0_i[55:48] : 1'b0;
  assign N6 = sel_i[6];
  assign data_o[63:56] = (N7)? data1_i[63:56] : 
                         (N23)? data0_i[63:56] : 1'b0;
  assign N7 = sel_i[7];
  assign data_o[71:64] = (N8)? data1_i[71:64] : 
                         (N24)? data0_i[71:64] : 1'b0;
  assign N8 = sel_i[8];
  assign data_o[79:72] = (N9)? data1_i[79:72] : 
                         (N25)? data0_i[79:72] : 1'b0;
  assign N9 = sel_i[9];
  assign data_o[87:80] = (N10)? data1_i[87:80] : 
                         (N26)? data0_i[87:80] : 1'b0;
  assign N10 = sel_i[10];
  assign data_o[95:88] = (N11)? data1_i[95:88] : 
                         (N27)? data0_i[95:88] : 1'b0;
  assign N11 = sel_i[11];
  assign data_o[103:96] = (N12)? data1_i[103:96] : 
                          (N28)? data0_i[103:96] : 1'b0;
  assign N12 = sel_i[12];
  assign data_o[111:104] = (N13)? data1_i[111:104] : 
                           (N29)? data0_i[111:104] : 1'b0;
  assign N13 = sel_i[13];
  assign data_o[119:112] = (N14)? data1_i[119:112] : 
                           (N30)? data0_i[119:112] : 1'b0;
  assign N14 = sel_i[14];
  assign data_o[127:120] = (N15)? data1_i[127:120] : 
                           (N31)? data0_i[127:120] : 1'b0;
  assign N15 = sel_i[15];
  assign N16 = ~sel_i[0];
  assign N17 = ~sel_i[1];
  assign N18 = ~sel_i[2];
  assign N19 = ~sel_i[3];
  assign N20 = ~sel_i[4];
  assign N21 = ~sel_i[5];
  assign N22 = ~sel_i[6];
  assign N23 = ~sel_i[7];
  assign N24 = ~sel_i[8];
  assign N25 = ~sel_i[9];
  assign N26 = ~sel_i[10];
  assign N27 = ~sel_i[11];
  assign N28 = ~sel_i[12];
  assign N29 = ~sel_i[13];
  assign N30 = ~sel_i[14];
  assign N31 = ~sel_i[15];

endmodule



module bsg_cache_sbuf_00000080_00000021_00000008
(
  clk_i,
  reset_i,
  sbuf_entry_i,
  v_i,
  sbuf_entry_o,
  v_o,
  yumi_i,
  empty_o,
  full_o,
  bypass_addr_i,
  bypass_v_i,
  bypass_data_o,
  bypass_mask_o
);

  input [179:0] sbuf_entry_i;
  output [179:0] sbuf_entry_o;
  input [32:0] bypass_addr_i;
  output [127:0] bypass_data_o;
  output [15:0] bypass_mask_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input bypass_v_i;
  output v_o;
  output empty_o;
  output full_o;
  wire [179:0] sbuf_entry_o,el0,el1;
  wire [127:0] bypass_data_o,el0or1_data,bypass_data_n;
  wire [15:0] bypass_mask_o,bypass_mask_n;
  wire v_o,empty_o,full_o,N0,el0_valid,el1_valid,tag_hit0_n,tag_hit1_n,tag_hit2_n,
  _2_net__15_,_2_net__14_,_2_net__13_,_2_net__12_,_2_net__11_,_2_net__10_,_2_net__9_,
  _2_net__8_,_2_net__7_,_2_net__6_,_2_net__5_,_2_net__4_,_2_net__3_,_2_net__2_,
  _2_net__1_,_2_net__0_,_4_net__15_,_4_net__14_,_4_net__13_,_4_net__12_,_4_net__11_,
  _4_net__10_,_4_net__9_,_4_net__8_,_4_net__7_,_4_net__6_,_4_net__5_,_4_net__4_,
  _4_net__3_,_4_net__2_,_4_net__1_,_4_net__0_,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,
  N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,
  N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,
  N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67;
  wire [15:15] tag_hit0x4,tag_hit1x4,tag_hit2x4;
  reg bypass_data_o_127_sv2v_reg,bypass_data_o_126_sv2v_reg,
  bypass_data_o_125_sv2v_reg,bypass_data_o_124_sv2v_reg,bypass_data_o_123_sv2v_reg,
  bypass_data_o_122_sv2v_reg,bypass_data_o_121_sv2v_reg,bypass_data_o_120_sv2v_reg,
  bypass_data_o_119_sv2v_reg,bypass_data_o_118_sv2v_reg,bypass_data_o_117_sv2v_reg,
  bypass_data_o_116_sv2v_reg,bypass_data_o_115_sv2v_reg,bypass_data_o_114_sv2v_reg,
  bypass_data_o_113_sv2v_reg,bypass_data_o_112_sv2v_reg,bypass_data_o_111_sv2v_reg,
  bypass_data_o_110_sv2v_reg,bypass_data_o_109_sv2v_reg,bypass_data_o_108_sv2v_reg,
  bypass_data_o_107_sv2v_reg,bypass_data_o_106_sv2v_reg,bypass_data_o_105_sv2v_reg,
  bypass_data_o_104_sv2v_reg,bypass_data_o_103_sv2v_reg,bypass_data_o_102_sv2v_reg,
  bypass_data_o_101_sv2v_reg,bypass_data_o_100_sv2v_reg,bypass_data_o_99_sv2v_reg,
  bypass_data_o_98_sv2v_reg,bypass_data_o_97_sv2v_reg,bypass_data_o_96_sv2v_reg,
  bypass_data_o_95_sv2v_reg,bypass_data_o_94_sv2v_reg,bypass_data_o_93_sv2v_reg,
  bypass_data_o_92_sv2v_reg,bypass_data_o_91_sv2v_reg,bypass_data_o_90_sv2v_reg,
  bypass_data_o_89_sv2v_reg,bypass_data_o_88_sv2v_reg,bypass_data_o_87_sv2v_reg,bypass_data_o_86_sv2v_reg,
  bypass_data_o_85_sv2v_reg,bypass_data_o_84_sv2v_reg,bypass_data_o_83_sv2v_reg,
  bypass_data_o_82_sv2v_reg,bypass_data_o_81_sv2v_reg,bypass_data_o_80_sv2v_reg,
  bypass_data_o_79_sv2v_reg,bypass_data_o_78_sv2v_reg,bypass_data_o_77_sv2v_reg,
  bypass_data_o_76_sv2v_reg,bypass_data_o_75_sv2v_reg,bypass_data_o_74_sv2v_reg,
  bypass_data_o_73_sv2v_reg,bypass_data_o_72_sv2v_reg,bypass_data_o_71_sv2v_reg,
  bypass_data_o_70_sv2v_reg,bypass_data_o_69_sv2v_reg,bypass_data_o_68_sv2v_reg,
  bypass_data_o_67_sv2v_reg,bypass_data_o_66_sv2v_reg,bypass_data_o_65_sv2v_reg,
  bypass_data_o_64_sv2v_reg,bypass_data_o_63_sv2v_reg,bypass_data_o_62_sv2v_reg,
  bypass_data_o_61_sv2v_reg,bypass_data_o_60_sv2v_reg,bypass_data_o_59_sv2v_reg,
  bypass_data_o_58_sv2v_reg,bypass_data_o_57_sv2v_reg,bypass_data_o_56_sv2v_reg,
  bypass_data_o_55_sv2v_reg,bypass_data_o_54_sv2v_reg,bypass_data_o_53_sv2v_reg,
  bypass_data_o_52_sv2v_reg,bypass_data_o_51_sv2v_reg,bypass_data_o_50_sv2v_reg,
  bypass_data_o_49_sv2v_reg,bypass_data_o_48_sv2v_reg,bypass_data_o_47_sv2v_reg,bypass_data_o_46_sv2v_reg,
  bypass_data_o_45_sv2v_reg,bypass_data_o_44_sv2v_reg,bypass_data_o_43_sv2v_reg,
  bypass_data_o_42_sv2v_reg,bypass_data_o_41_sv2v_reg,bypass_data_o_40_sv2v_reg,
  bypass_data_o_39_sv2v_reg,bypass_data_o_38_sv2v_reg,bypass_data_o_37_sv2v_reg,
  bypass_data_o_36_sv2v_reg,bypass_data_o_35_sv2v_reg,bypass_data_o_34_sv2v_reg,
  bypass_data_o_33_sv2v_reg,bypass_data_o_32_sv2v_reg,bypass_data_o_31_sv2v_reg,
  bypass_data_o_30_sv2v_reg,bypass_data_o_29_sv2v_reg,bypass_data_o_28_sv2v_reg,
  bypass_data_o_27_sv2v_reg,bypass_data_o_26_sv2v_reg,bypass_data_o_25_sv2v_reg,
  bypass_data_o_24_sv2v_reg,bypass_data_o_23_sv2v_reg,bypass_data_o_22_sv2v_reg,
  bypass_data_o_21_sv2v_reg,bypass_data_o_20_sv2v_reg,bypass_data_o_19_sv2v_reg,
  bypass_data_o_18_sv2v_reg,bypass_data_o_17_sv2v_reg,bypass_data_o_16_sv2v_reg,
  bypass_data_o_15_sv2v_reg,bypass_data_o_14_sv2v_reg,bypass_data_o_13_sv2v_reg,
  bypass_data_o_12_sv2v_reg,bypass_data_o_11_sv2v_reg,bypass_data_o_10_sv2v_reg,
  bypass_data_o_9_sv2v_reg,bypass_data_o_8_sv2v_reg,bypass_data_o_7_sv2v_reg,bypass_data_o_6_sv2v_reg,
  bypass_data_o_5_sv2v_reg,bypass_data_o_4_sv2v_reg,bypass_data_o_3_sv2v_reg,
  bypass_data_o_2_sv2v_reg,bypass_data_o_1_sv2v_reg,bypass_data_o_0_sv2v_reg,
  bypass_mask_o_15_sv2v_reg,bypass_mask_o_14_sv2v_reg,bypass_mask_o_13_sv2v_reg,
  bypass_mask_o_12_sv2v_reg,bypass_mask_o_11_sv2v_reg,bypass_mask_o_10_sv2v_reg,
  bypass_mask_o_9_sv2v_reg,bypass_mask_o_8_sv2v_reg,bypass_mask_o_7_sv2v_reg,
  bypass_mask_o_6_sv2v_reg,bypass_mask_o_5_sv2v_reg,bypass_mask_o_4_sv2v_reg,bypass_mask_o_3_sv2v_reg,
  bypass_mask_o_2_sv2v_reg,bypass_mask_o_1_sv2v_reg,bypass_mask_o_0_sv2v_reg;
  assign bypass_data_o[127] = bypass_data_o_127_sv2v_reg;
  assign bypass_data_o[126] = bypass_data_o_126_sv2v_reg;
  assign bypass_data_o[125] = bypass_data_o_125_sv2v_reg;
  assign bypass_data_o[124] = bypass_data_o_124_sv2v_reg;
  assign bypass_data_o[123] = bypass_data_o_123_sv2v_reg;
  assign bypass_data_o[122] = bypass_data_o_122_sv2v_reg;
  assign bypass_data_o[121] = bypass_data_o_121_sv2v_reg;
  assign bypass_data_o[120] = bypass_data_o_120_sv2v_reg;
  assign bypass_data_o[119] = bypass_data_o_119_sv2v_reg;
  assign bypass_data_o[118] = bypass_data_o_118_sv2v_reg;
  assign bypass_data_o[117] = bypass_data_o_117_sv2v_reg;
  assign bypass_data_o[116] = bypass_data_o_116_sv2v_reg;
  assign bypass_data_o[115] = bypass_data_o_115_sv2v_reg;
  assign bypass_data_o[114] = bypass_data_o_114_sv2v_reg;
  assign bypass_data_o[113] = bypass_data_o_113_sv2v_reg;
  assign bypass_data_o[112] = bypass_data_o_112_sv2v_reg;
  assign bypass_data_o[111] = bypass_data_o_111_sv2v_reg;
  assign bypass_data_o[110] = bypass_data_o_110_sv2v_reg;
  assign bypass_data_o[109] = bypass_data_o_109_sv2v_reg;
  assign bypass_data_o[108] = bypass_data_o_108_sv2v_reg;
  assign bypass_data_o[107] = bypass_data_o_107_sv2v_reg;
  assign bypass_data_o[106] = bypass_data_o_106_sv2v_reg;
  assign bypass_data_o[105] = bypass_data_o_105_sv2v_reg;
  assign bypass_data_o[104] = bypass_data_o_104_sv2v_reg;
  assign bypass_data_o[103] = bypass_data_o_103_sv2v_reg;
  assign bypass_data_o[102] = bypass_data_o_102_sv2v_reg;
  assign bypass_data_o[101] = bypass_data_o_101_sv2v_reg;
  assign bypass_data_o[100] = bypass_data_o_100_sv2v_reg;
  assign bypass_data_o[99] = bypass_data_o_99_sv2v_reg;
  assign bypass_data_o[98] = bypass_data_o_98_sv2v_reg;
  assign bypass_data_o[97] = bypass_data_o_97_sv2v_reg;
  assign bypass_data_o[96] = bypass_data_o_96_sv2v_reg;
  assign bypass_data_o[95] = bypass_data_o_95_sv2v_reg;
  assign bypass_data_o[94] = bypass_data_o_94_sv2v_reg;
  assign bypass_data_o[93] = bypass_data_o_93_sv2v_reg;
  assign bypass_data_o[92] = bypass_data_o_92_sv2v_reg;
  assign bypass_data_o[91] = bypass_data_o_91_sv2v_reg;
  assign bypass_data_o[90] = bypass_data_o_90_sv2v_reg;
  assign bypass_data_o[89] = bypass_data_o_89_sv2v_reg;
  assign bypass_data_o[88] = bypass_data_o_88_sv2v_reg;
  assign bypass_data_o[87] = bypass_data_o_87_sv2v_reg;
  assign bypass_data_o[86] = bypass_data_o_86_sv2v_reg;
  assign bypass_data_o[85] = bypass_data_o_85_sv2v_reg;
  assign bypass_data_o[84] = bypass_data_o_84_sv2v_reg;
  assign bypass_data_o[83] = bypass_data_o_83_sv2v_reg;
  assign bypass_data_o[82] = bypass_data_o_82_sv2v_reg;
  assign bypass_data_o[81] = bypass_data_o_81_sv2v_reg;
  assign bypass_data_o[80] = bypass_data_o_80_sv2v_reg;
  assign bypass_data_o[79] = bypass_data_o_79_sv2v_reg;
  assign bypass_data_o[78] = bypass_data_o_78_sv2v_reg;
  assign bypass_data_o[77] = bypass_data_o_77_sv2v_reg;
  assign bypass_data_o[76] = bypass_data_o_76_sv2v_reg;
  assign bypass_data_o[75] = bypass_data_o_75_sv2v_reg;
  assign bypass_data_o[74] = bypass_data_o_74_sv2v_reg;
  assign bypass_data_o[73] = bypass_data_o_73_sv2v_reg;
  assign bypass_data_o[72] = bypass_data_o_72_sv2v_reg;
  assign bypass_data_o[71] = bypass_data_o_71_sv2v_reg;
  assign bypass_data_o[70] = bypass_data_o_70_sv2v_reg;
  assign bypass_data_o[69] = bypass_data_o_69_sv2v_reg;
  assign bypass_data_o[68] = bypass_data_o_68_sv2v_reg;
  assign bypass_data_o[67] = bypass_data_o_67_sv2v_reg;
  assign bypass_data_o[66] = bypass_data_o_66_sv2v_reg;
  assign bypass_data_o[65] = bypass_data_o_65_sv2v_reg;
  assign bypass_data_o[64] = bypass_data_o_64_sv2v_reg;
  assign bypass_data_o[63] = bypass_data_o_63_sv2v_reg;
  assign bypass_data_o[62] = bypass_data_o_62_sv2v_reg;
  assign bypass_data_o[61] = bypass_data_o_61_sv2v_reg;
  assign bypass_data_o[60] = bypass_data_o_60_sv2v_reg;
  assign bypass_data_o[59] = bypass_data_o_59_sv2v_reg;
  assign bypass_data_o[58] = bypass_data_o_58_sv2v_reg;
  assign bypass_data_o[57] = bypass_data_o_57_sv2v_reg;
  assign bypass_data_o[56] = bypass_data_o_56_sv2v_reg;
  assign bypass_data_o[55] = bypass_data_o_55_sv2v_reg;
  assign bypass_data_o[54] = bypass_data_o_54_sv2v_reg;
  assign bypass_data_o[53] = bypass_data_o_53_sv2v_reg;
  assign bypass_data_o[52] = bypass_data_o_52_sv2v_reg;
  assign bypass_data_o[51] = bypass_data_o_51_sv2v_reg;
  assign bypass_data_o[50] = bypass_data_o_50_sv2v_reg;
  assign bypass_data_o[49] = bypass_data_o_49_sv2v_reg;
  assign bypass_data_o[48] = bypass_data_o_48_sv2v_reg;
  assign bypass_data_o[47] = bypass_data_o_47_sv2v_reg;
  assign bypass_data_o[46] = bypass_data_o_46_sv2v_reg;
  assign bypass_data_o[45] = bypass_data_o_45_sv2v_reg;
  assign bypass_data_o[44] = bypass_data_o_44_sv2v_reg;
  assign bypass_data_o[43] = bypass_data_o_43_sv2v_reg;
  assign bypass_data_o[42] = bypass_data_o_42_sv2v_reg;
  assign bypass_data_o[41] = bypass_data_o_41_sv2v_reg;
  assign bypass_data_o[40] = bypass_data_o_40_sv2v_reg;
  assign bypass_data_o[39] = bypass_data_o_39_sv2v_reg;
  assign bypass_data_o[38] = bypass_data_o_38_sv2v_reg;
  assign bypass_data_o[37] = bypass_data_o_37_sv2v_reg;
  assign bypass_data_o[36] = bypass_data_o_36_sv2v_reg;
  assign bypass_data_o[35] = bypass_data_o_35_sv2v_reg;
  assign bypass_data_o[34] = bypass_data_o_34_sv2v_reg;
  assign bypass_data_o[33] = bypass_data_o_33_sv2v_reg;
  assign bypass_data_o[32] = bypass_data_o_32_sv2v_reg;
  assign bypass_data_o[31] = bypass_data_o_31_sv2v_reg;
  assign bypass_data_o[30] = bypass_data_o_30_sv2v_reg;
  assign bypass_data_o[29] = bypass_data_o_29_sv2v_reg;
  assign bypass_data_o[28] = bypass_data_o_28_sv2v_reg;
  assign bypass_data_o[27] = bypass_data_o_27_sv2v_reg;
  assign bypass_data_o[26] = bypass_data_o_26_sv2v_reg;
  assign bypass_data_o[25] = bypass_data_o_25_sv2v_reg;
  assign bypass_data_o[24] = bypass_data_o_24_sv2v_reg;
  assign bypass_data_o[23] = bypass_data_o_23_sv2v_reg;
  assign bypass_data_o[22] = bypass_data_o_22_sv2v_reg;
  assign bypass_data_o[21] = bypass_data_o_21_sv2v_reg;
  assign bypass_data_o[20] = bypass_data_o_20_sv2v_reg;
  assign bypass_data_o[19] = bypass_data_o_19_sv2v_reg;
  assign bypass_data_o[18] = bypass_data_o_18_sv2v_reg;
  assign bypass_data_o[17] = bypass_data_o_17_sv2v_reg;
  assign bypass_data_o[16] = bypass_data_o_16_sv2v_reg;
  assign bypass_data_o[15] = bypass_data_o_15_sv2v_reg;
  assign bypass_data_o[14] = bypass_data_o_14_sv2v_reg;
  assign bypass_data_o[13] = bypass_data_o_13_sv2v_reg;
  assign bypass_data_o[12] = bypass_data_o_12_sv2v_reg;
  assign bypass_data_o[11] = bypass_data_o_11_sv2v_reg;
  assign bypass_data_o[10] = bypass_data_o_10_sv2v_reg;
  assign bypass_data_o[9] = bypass_data_o_9_sv2v_reg;
  assign bypass_data_o[8] = bypass_data_o_8_sv2v_reg;
  assign bypass_data_o[7] = bypass_data_o_7_sv2v_reg;
  assign bypass_data_o[6] = bypass_data_o_6_sv2v_reg;
  assign bypass_data_o[5] = bypass_data_o_5_sv2v_reg;
  assign bypass_data_o[4] = bypass_data_o_4_sv2v_reg;
  assign bypass_data_o[3] = bypass_data_o_3_sv2v_reg;
  assign bypass_data_o[2] = bypass_data_o_2_sv2v_reg;
  assign bypass_data_o[1] = bypass_data_o_1_sv2v_reg;
  assign bypass_data_o[0] = bypass_data_o_0_sv2v_reg;
  assign bypass_mask_o[15] = bypass_mask_o_15_sv2v_reg;
  assign bypass_mask_o[14] = bypass_mask_o_14_sv2v_reg;
  assign bypass_mask_o[13] = bypass_mask_o_13_sv2v_reg;
  assign bypass_mask_o[12] = bypass_mask_o_12_sv2v_reg;
  assign bypass_mask_o[11] = bypass_mask_o_11_sv2v_reg;
  assign bypass_mask_o[10] = bypass_mask_o_10_sv2v_reg;
  assign bypass_mask_o[9] = bypass_mask_o_9_sv2v_reg;
  assign bypass_mask_o[8] = bypass_mask_o_8_sv2v_reg;
  assign bypass_mask_o[7] = bypass_mask_o_7_sv2v_reg;
  assign bypass_mask_o[6] = bypass_mask_o_6_sv2v_reg;
  assign bypass_mask_o[5] = bypass_mask_o_5_sv2v_reg;
  assign bypass_mask_o[4] = bypass_mask_o_4_sv2v_reg;
  assign bypass_mask_o[3] = bypass_mask_o_3_sv2v_reg;
  assign bypass_mask_o[2] = bypass_mask_o_2_sv2v_reg;
  assign bypass_mask_o[1] = bypass_mask_o_1_sv2v_reg;
  assign bypass_mask_o[0] = bypass_mask_o_0_sv2v_reg;

  bsg_cache_buffer_queue_000000b4
  q0
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .data_i(sbuf_entry_i),
    .v_o(v_o),
    .data_o(sbuf_entry_o),
    .yumi_i(yumi_i),
    .el0_valid_o(el0_valid),
    .el1_valid_o(el1_valid),
    .el0_snoop_o(el0),
    .el1_snoop_o(el1),
    .empty_o(empty_o),
    .full_o(full_o)
  );

  assign tag_hit0_n = bypass_addr_i[32:4] == el0[179:151];
  assign tag_hit1_n = bypass_addr_i[32:4] == el1[179:151];
  assign tag_hit2_n = bypass_addr_i[32:4] == sbuf_entry_i[179:151];

  bsg_mux_segmented_00000010_8
  mux_segmented_merge0
  (
    .data0_i(el1[146:19]),
    .data1_i(el0[146:19]),
    .sel_i({ _2_net__15_, _2_net__14_, _2_net__13_, _2_net__12_, _2_net__11_, _2_net__10_, _2_net__9_, _2_net__8_, _2_net__7_, _2_net__6_, _2_net__5_, _2_net__4_, _2_net__3_, _2_net__2_, _2_net__1_, _2_net__0_ }),
    .data_o(el0or1_data)
  );


  bsg_mux_segmented_00000010_8
  mux_segmented_merge1
  (
    .data0_i(el0or1_data),
    .data1_i(sbuf_entry_i[146:19]),
    .sel_i({ _4_net__15_, _4_net__14_, _4_net__13_, _4_net__12_, _4_net__11_, _4_net__10_, _4_net__9_, _4_net__8_, _4_net__7_, _4_net__6_, _4_net__5_, _4_net__4_, _4_net__3_, _4_net__2_, _4_net__1_, _4_net__0_ }),
    .data_o(bypass_data_n)
  );

  assign { N3, N2 } = (N0)? { 1'b1, 1'b1 } : 
                      (N1)? { 1'b0, 1'b0 } : 1'b0;
  assign N0 = bypass_v_i;
  assign tag_hit0x4[15] = tag_hit0_n & el0_valid;
  assign tag_hit1x4[15] = tag_hit1_n & el1_valid;
  assign tag_hit2x4[15] = tag_hit2_n & v_i;
  assign bypass_mask_n[15] = N6 | N7;
  assign N6 = N4 | N5;
  assign N4 = tag_hit0x4[15] & el0[18];
  assign N5 = tag_hit1x4[15] & el1[18];
  assign N7 = tag_hit2x4[15] & sbuf_entry_i[18];
  assign bypass_mask_n[14] = N10 | N11;
  assign N10 = N8 | N9;
  assign N8 = tag_hit0x4[15] & el0[17];
  assign N9 = tag_hit1x4[15] & el1[17];
  assign N11 = tag_hit2x4[15] & sbuf_entry_i[17];
  assign bypass_mask_n[13] = N14 | N15;
  assign N14 = N12 | N13;
  assign N12 = tag_hit0x4[15] & el0[16];
  assign N13 = tag_hit1x4[15] & el1[16];
  assign N15 = tag_hit2x4[15] & sbuf_entry_i[16];
  assign bypass_mask_n[12] = N18 | N19;
  assign N18 = N16 | N17;
  assign N16 = tag_hit0x4[15] & el0[15];
  assign N17 = tag_hit1x4[15] & el1[15];
  assign N19 = tag_hit2x4[15] & sbuf_entry_i[15];
  assign bypass_mask_n[11] = N22 | N23;
  assign N22 = N20 | N21;
  assign N20 = tag_hit0x4[15] & el0[14];
  assign N21 = tag_hit1x4[15] & el1[14];
  assign N23 = tag_hit2x4[15] & sbuf_entry_i[14];
  assign bypass_mask_n[10] = N26 | N27;
  assign N26 = N24 | N25;
  assign N24 = tag_hit0x4[15] & el0[13];
  assign N25 = tag_hit1x4[15] & el1[13];
  assign N27 = tag_hit2x4[15] & sbuf_entry_i[13];
  assign bypass_mask_n[9] = N30 | N31;
  assign N30 = N28 | N29;
  assign N28 = tag_hit0x4[15] & el0[12];
  assign N29 = tag_hit1x4[15] & el1[12];
  assign N31 = tag_hit2x4[15] & sbuf_entry_i[12];
  assign bypass_mask_n[8] = N34 | N35;
  assign N34 = N32 | N33;
  assign N32 = tag_hit0x4[15] & el0[11];
  assign N33 = tag_hit1x4[15] & el1[11];
  assign N35 = tag_hit2x4[15] & sbuf_entry_i[11];
  assign bypass_mask_n[7] = N38 | N39;
  assign N38 = N36 | N37;
  assign N36 = tag_hit0x4[15] & el0[10];
  assign N37 = tag_hit1x4[15] & el1[10];
  assign N39 = tag_hit2x4[15] & sbuf_entry_i[10];
  assign bypass_mask_n[6] = N42 | N43;
  assign N42 = N40 | N41;
  assign N40 = tag_hit0x4[15] & el0[9];
  assign N41 = tag_hit1x4[15] & el1[9];
  assign N43 = tag_hit2x4[15] & sbuf_entry_i[9];
  assign bypass_mask_n[5] = N46 | N47;
  assign N46 = N44 | N45;
  assign N44 = tag_hit0x4[15] & el0[8];
  assign N45 = tag_hit1x4[15] & el1[8];
  assign N47 = tag_hit2x4[15] & sbuf_entry_i[8];
  assign bypass_mask_n[4] = N50 | N51;
  assign N50 = N48 | N49;
  assign N48 = tag_hit0x4[15] & el0[7];
  assign N49 = tag_hit1x4[15] & el1[7];
  assign N51 = tag_hit2x4[15] & sbuf_entry_i[7];
  assign bypass_mask_n[3] = N54 | N55;
  assign N54 = N52 | N53;
  assign N52 = tag_hit0x4[15] & el0[6];
  assign N53 = tag_hit1x4[15] & el1[6];
  assign N55 = tag_hit2x4[15] & sbuf_entry_i[6];
  assign bypass_mask_n[2] = N58 | N59;
  assign N58 = N56 | N57;
  assign N56 = tag_hit0x4[15] & el0[5];
  assign N57 = tag_hit1x4[15] & el1[5];
  assign N59 = tag_hit2x4[15] & sbuf_entry_i[5];
  assign bypass_mask_n[1] = N62 | N63;
  assign N62 = N60 | N61;
  assign N60 = tag_hit0x4[15] & el0[4];
  assign N61 = tag_hit1x4[15] & el1[4];
  assign N63 = tag_hit2x4[15] & sbuf_entry_i[4];
  assign bypass_mask_n[0] = N66 | N67;
  assign N66 = N64 | N65;
  assign N64 = tag_hit0x4[15] & el0[3];
  assign N65 = tag_hit1x4[15] & el1[3];
  assign N67 = tag_hit2x4[15] & sbuf_entry_i[3];
  assign _2_net__15_ = tag_hit0x4[15] & el0[18];
  assign _2_net__14_ = tag_hit0x4[15] & el0[17];
  assign _2_net__13_ = tag_hit0x4[15] & el0[16];
  assign _2_net__12_ = tag_hit0x4[15] & el0[15];
  assign _2_net__11_ = tag_hit0x4[15] & el0[14];
  assign _2_net__10_ = tag_hit0x4[15] & el0[13];
  assign _2_net__9_ = tag_hit0x4[15] & el0[12];
  assign _2_net__8_ = tag_hit0x4[15] & el0[11];
  assign _2_net__7_ = tag_hit0x4[15] & el0[10];
  assign _2_net__6_ = tag_hit0x4[15] & el0[9];
  assign _2_net__5_ = tag_hit0x4[15] & el0[8];
  assign _2_net__4_ = tag_hit0x4[15] & el0[7];
  assign _2_net__3_ = tag_hit0x4[15] & el0[6];
  assign _2_net__2_ = tag_hit0x4[15] & el0[5];
  assign _2_net__1_ = tag_hit0x4[15] & el0[4];
  assign _2_net__0_ = tag_hit0x4[15] & el0[3];
  assign _4_net__15_ = tag_hit2x4[15] & sbuf_entry_i[18];
  assign _4_net__14_ = tag_hit2x4[15] & sbuf_entry_i[17];
  assign _4_net__13_ = tag_hit2x4[15] & sbuf_entry_i[16];
  assign _4_net__12_ = tag_hit2x4[15] & sbuf_entry_i[15];
  assign _4_net__11_ = tag_hit2x4[15] & sbuf_entry_i[14];
  assign _4_net__10_ = tag_hit2x4[15] & sbuf_entry_i[13];
  assign _4_net__9_ = tag_hit2x4[15] & sbuf_entry_i[12];
  assign _4_net__8_ = tag_hit2x4[15] & sbuf_entry_i[11];
  assign _4_net__7_ = tag_hit2x4[15] & sbuf_entry_i[10];
  assign _4_net__6_ = tag_hit2x4[15] & sbuf_entry_i[9];
  assign _4_net__5_ = tag_hit2x4[15] & sbuf_entry_i[8];
  assign _4_net__4_ = tag_hit2x4[15] & sbuf_entry_i[7];
  assign _4_net__3_ = tag_hit2x4[15] & sbuf_entry_i[6];
  assign _4_net__2_ = tag_hit2x4[15] & sbuf_entry_i[5];
  assign _4_net__1_ = tag_hit2x4[15] & sbuf_entry_i[4];
  assign _4_net__0_ = tag_hit2x4[15] & sbuf_entry_i[3];
  assign N1 = ~bypass_v_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      bypass_data_o_127_sv2v_reg <= 1'b0;
      bypass_data_o_126_sv2v_reg <= 1'b0;
      bypass_data_o_125_sv2v_reg <= 1'b0;
      bypass_data_o_124_sv2v_reg <= 1'b0;
      bypass_data_o_123_sv2v_reg <= 1'b0;
      bypass_data_o_122_sv2v_reg <= 1'b0;
      bypass_data_o_121_sv2v_reg <= 1'b0;
      bypass_data_o_120_sv2v_reg <= 1'b0;
      bypass_data_o_119_sv2v_reg <= 1'b0;
      bypass_data_o_118_sv2v_reg <= 1'b0;
      bypass_data_o_117_sv2v_reg <= 1'b0;
      bypass_data_o_116_sv2v_reg <= 1'b0;
      bypass_data_o_115_sv2v_reg <= 1'b0;
      bypass_data_o_114_sv2v_reg <= 1'b0;
      bypass_data_o_113_sv2v_reg <= 1'b0;
      bypass_data_o_112_sv2v_reg <= 1'b0;
      bypass_data_o_111_sv2v_reg <= 1'b0;
      bypass_data_o_110_sv2v_reg <= 1'b0;
      bypass_data_o_109_sv2v_reg <= 1'b0;
      bypass_data_o_108_sv2v_reg <= 1'b0;
      bypass_data_o_107_sv2v_reg <= 1'b0;
      bypass_data_o_106_sv2v_reg <= 1'b0;
      bypass_data_o_105_sv2v_reg <= 1'b0;
      bypass_data_o_104_sv2v_reg <= 1'b0;
      bypass_data_o_103_sv2v_reg <= 1'b0;
      bypass_data_o_102_sv2v_reg <= 1'b0;
      bypass_data_o_101_sv2v_reg <= 1'b0;
      bypass_data_o_100_sv2v_reg <= 1'b0;
      bypass_data_o_99_sv2v_reg <= 1'b0;
      bypass_data_o_98_sv2v_reg <= 1'b0;
      bypass_data_o_97_sv2v_reg <= 1'b0;
      bypass_data_o_96_sv2v_reg <= 1'b0;
      bypass_data_o_95_sv2v_reg <= 1'b0;
      bypass_data_o_94_sv2v_reg <= 1'b0;
      bypass_data_o_93_sv2v_reg <= 1'b0;
      bypass_data_o_92_sv2v_reg <= 1'b0;
      bypass_data_o_91_sv2v_reg <= 1'b0;
      bypass_data_o_90_sv2v_reg <= 1'b0;
      bypass_data_o_89_sv2v_reg <= 1'b0;
      bypass_data_o_88_sv2v_reg <= 1'b0;
      bypass_data_o_87_sv2v_reg <= 1'b0;
      bypass_data_o_86_sv2v_reg <= 1'b0;
      bypass_data_o_85_sv2v_reg <= 1'b0;
      bypass_data_o_84_sv2v_reg <= 1'b0;
      bypass_data_o_83_sv2v_reg <= 1'b0;
      bypass_data_o_82_sv2v_reg <= 1'b0;
      bypass_data_o_81_sv2v_reg <= 1'b0;
      bypass_data_o_80_sv2v_reg <= 1'b0;
      bypass_data_o_79_sv2v_reg <= 1'b0;
      bypass_data_o_78_sv2v_reg <= 1'b0;
      bypass_data_o_77_sv2v_reg <= 1'b0;
      bypass_data_o_76_sv2v_reg <= 1'b0;
      bypass_data_o_75_sv2v_reg <= 1'b0;
      bypass_data_o_74_sv2v_reg <= 1'b0;
      bypass_data_o_73_sv2v_reg <= 1'b0;
      bypass_data_o_72_sv2v_reg <= 1'b0;
      bypass_data_o_71_sv2v_reg <= 1'b0;
      bypass_data_o_70_sv2v_reg <= 1'b0;
      bypass_data_o_69_sv2v_reg <= 1'b0;
      bypass_data_o_68_sv2v_reg <= 1'b0;
      bypass_data_o_67_sv2v_reg <= 1'b0;
      bypass_data_o_66_sv2v_reg <= 1'b0;
      bypass_data_o_65_sv2v_reg <= 1'b0;
      bypass_data_o_64_sv2v_reg <= 1'b0;
      bypass_data_o_63_sv2v_reg <= 1'b0;
      bypass_data_o_62_sv2v_reg <= 1'b0;
      bypass_data_o_61_sv2v_reg <= 1'b0;
      bypass_data_o_60_sv2v_reg <= 1'b0;
      bypass_data_o_59_sv2v_reg <= 1'b0;
      bypass_data_o_58_sv2v_reg <= 1'b0;
      bypass_data_o_57_sv2v_reg <= 1'b0;
      bypass_data_o_56_sv2v_reg <= 1'b0;
      bypass_data_o_55_sv2v_reg <= 1'b0;
      bypass_data_o_54_sv2v_reg <= 1'b0;
      bypass_data_o_53_sv2v_reg <= 1'b0;
      bypass_data_o_52_sv2v_reg <= 1'b0;
      bypass_data_o_51_sv2v_reg <= 1'b0;
      bypass_data_o_50_sv2v_reg <= 1'b0;
      bypass_data_o_49_sv2v_reg <= 1'b0;
      bypass_data_o_48_sv2v_reg <= 1'b0;
      bypass_data_o_47_sv2v_reg <= 1'b0;
      bypass_data_o_46_sv2v_reg <= 1'b0;
      bypass_data_o_45_sv2v_reg <= 1'b0;
      bypass_data_o_44_sv2v_reg <= 1'b0;
      bypass_data_o_43_sv2v_reg <= 1'b0;
      bypass_data_o_42_sv2v_reg <= 1'b0;
      bypass_data_o_41_sv2v_reg <= 1'b0;
      bypass_data_o_40_sv2v_reg <= 1'b0;
      bypass_data_o_39_sv2v_reg <= 1'b0;
      bypass_data_o_38_sv2v_reg <= 1'b0;
      bypass_data_o_37_sv2v_reg <= 1'b0;
      bypass_data_o_36_sv2v_reg <= 1'b0;
      bypass_data_o_35_sv2v_reg <= 1'b0;
      bypass_data_o_34_sv2v_reg <= 1'b0;
      bypass_data_o_33_sv2v_reg <= 1'b0;
      bypass_data_o_32_sv2v_reg <= 1'b0;
      bypass_data_o_31_sv2v_reg <= 1'b0;
      bypass_data_o_30_sv2v_reg <= 1'b0;
      bypass_data_o_29_sv2v_reg <= 1'b0;
      bypass_mask_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      bypass_data_o_127_sv2v_reg <= bypass_data_n[127];
      bypass_data_o_126_sv2v_reg <= bypass_data_n[126];
      bypass_data_o_125_sv2v_reg <= bypass_data_n[125];
      bypass_data_o_124_sv2v_reg <= bypass_data_n[124];
      bypass_data_o_123_sv2v_reg <= bypass_data_n[123];
      bypass_data_o_122_sv2v_reg <= bypass_data_n[122];
      bypass_data_o_121_sv2v_reg <= bypass_data_n[121];
      bypass_data_o_120_sv2v_reg <= bypass_data_n[120];
      bypass_data_o_119_sv2v_reg <= bypass_data_n[119];
      bypass_data_o_118_sv2v_reg <= bypass_data_n[118];
      bypass_data_o_117_sv2v_reg <= bypass_data_n[117];
      bypass_data_o_116_sv2v_reg <= bypass_data_n[116];
      bypass_data_o_115_sv2v_reg <= bypass_data_n[115];
      bypass_data_o_114_sv2v_reg <= bypass_data_n[114];
      bypass_data_o_113_sv2v_reg <= bypass_data_n[113];
      bypass_data_o_112_sv2v_reg <= bypass_data_n[112];
      bypass_data_o_111_sv2v_reg <= bypass_data_n[111];
      bypass_data_o_110_sv2v_reg <= bypass_data_n[110];
      bypass_data_o_109_sv2v_reg <= bypass_data_n[109];
      bypass_data_o_108_sv2v_reg <= bypass_data_n[108];
      bypass_data_o_107_sv2v_reg <= bypass_data_n[107];
      bypass_data_o_106_sv2v_reg <= bypass_data_n[106];
      bypass_data_o_105_sv2v_reg <= bypass_data_n[105];
      bypass_data_o_104_sv2v_reg <= bypass_data_n[104];
      bypass_data_o_103_sv2v_reg <= bypass_data_n[103];
      bypass_data_o_102_sv2v_reg <= bypass_data_n[102];
      bypass_data_o_101_sv2v_reg <= bypass_data_n[101];
      bypass_data_o_100_sv2v_reg <= bypass_data_n[100];
      bypass_data_o_99_sv2v_reg <= bypass_data_n[99];
      bypass_data_o_98_sv2v_reg <= bypass_data_n[98];
      bypass_data_o_97_sv2v_reg <= bypass_data_n[97];
      bypass_data_o_96_sv2v_reg <= bypass_data_n[96];
      bypass_data_o_95_sv2v_reg <= bypass_data_n[95];
      bypass_data_o_94_sv2v_reg <= bypass_data_n[94];
      bypass_data_o_93_sv2v_reg <= bypass_data_n[93];
      bypass_data_o_92_sv2v_reg <= bypass_data_n[92];
      bypass_data_o_91_sv2v_reg <= bypass_data_n[91];
      bypass_data_o_90_sv2v_reg <= bypass_data_n[90];
      bypass_data_o_89_sv2v_reg <= bypass_data_n[89];
      bypass_data_o_88_sv2v_reg <= bypass_data_n[88];
      bypass_data_o_87_sv2v_reg <= bypass_data_n[87];
      bypass_data_o_86_sv2v_reg <= bypass_data_n[86];
      bypass_data_o_85_sv2v_reg <= bypass_data_n[85];
      bypass_data_o_84_sv2v_reg <= bypass_data_n[84];
      bypass_data_o_83_sv2v_reg <= bypass_data_n[83];
      bypass_data_o_82_sv2v_reg <= bypass_data_n[82];
      bypass_data_o_81_sv2v_reg <= bypass_data_n[81];
      bypass_data_o_80_sv2v_reg <= bypass_data_n[80];
      bypass_data_o_79_sv2v_reg <= bypass_data_n[79];
      bypass_data_o_78_sv2v_reg <= bypass_data_n[78];
      bypass_data_o_77_sv2v_reg <= bypass_data_n[77];
      bypass_data_o_76_sv2v_reg <= bypass_data_n[76];
      bypass_data_o_75_sv2v_reg <= bypass_data_n[75];
      bypass_data_o_74_sv2v_reg <= bypass_data_n[74];
      bypass_data_o_73_sv2v_reg <= bypass_data_n[73];
      bypass_data_o_72_sv2v_reg <= bypass_data_n[72];
      bypass_data_o_71_sv2v_reg <= bypass_data_n[71];
      bypass_data_o_70_sv2v_reg <= bypass_data_n[70];
      bypass_data_o_69_sv2v_reg <= bypass_data_n[69];
      bypass_data_o_68_sv2v_reg <= bypass_data_n[68];
      bypass_data_o_67_sv2v_reg <= bypass_data_n[67];
      bypass_data_o_66_sv2v_reg <= bypass_data_n[66];
      bypass_data_o_65_sv2v_reg <= bypass_data_n[65];
      bypass_data_o_64_sv2v_reg <= bypass_data_n[64];
      bypass_data_o_63_sv2v_reg <= bypass_data_n[63];
      bypass_data_o_62_sv2v_reg <= bypass_data_n[62];
      bypass_data_o_61_sv2v_reg <= bypass_data_n[61];
      bypass_data_o_60_sv2v_reg <= bypass_data_n[60];
      bypass_data_o_59_sv2v_reg <= bypass_data_n[59];
      bypass_data_o_58_sv2v_reg <= bypass_data_n[58];
      bypass_data_o_57_sv2v_reg <= bypass_data_n[57];
      bypass_data_o_56_sv2v_reg <= bypass_data_n[56];
      bypass_data_o_55_sv2v_reg <= bypass_data_n[55];
      bypass_data_o_54_sv2v_reg <= bypass_data_n[54];
      bypass_data_o_53_sv2v_reg <= bypass_data_n[53];
      bypass_data_o_52_sv2v_reg <= bypass_data_n[52];
      bypass_data_o_51_sv2v_reg <= bypass_data_n[51];
      bypass_data_o_50_sv2v_reg <= bypass_data_n[50];
      bypass_data_o_49_sv2v_reg <= bypass_data_n[49];
      bypass_data_o_48_sv2v_reg <= bypass_data_n[48];
      bypass_data_o_47_sv2v_reg <= bypass_data_n[47];
      bypass_data_o_46_sv2v_reg <= bypass_data_n[46];
      bypass_data_o_45_sv2v_reg <= bypass_data_n[45];
      bypass_data_o_44_sv2v_reg <= bypass_data_n[44];
      bypass_data_o_43_sv2v_reg <= bypass_data_n[43];
      bypass_data_o_42_sv2v_reg <= bypass_data_n[42];
      bypass_data_o_41_sv2v_reg <= bypass_data_n[41];
      bypass_data_o_40_sv2v_reg <= bypass_data_n[40];
      bypass_data_o_39_sv2v_reg <= bypass_data_n[39];
      bypass_data_o_38_sv2v_reg <= bypass_data_n[38];
      bypass_data_o_37_sv2v_reg <= bypass_data_n[37];
      bypass_data_o_36_sv2v_reg <= bypass_data_n[36];
      bypass_data_o_35_sv2v_reg <= bypass_data_n[35];
      bypass_data_o_34_sv2v_reg <= bypass_data_n[34];
      bypass_data_o_33_sv2v_reg <= bypass_data_n[33];
      bypass_data_o_32_sv2v_reg <= bypass_data_n[32];
      bypass_data_o_31_sv2v_reg <= bypass_data_n[31];
      bypass_data_o_30_sv2v_reg <= bypass_data_n[30];
      bypass_data_o_29_sv2v_reg <= bypass_data_n[29];
      bypass_mask_o_0_sv2v_reg <= bypass_mask_n[0];
    end 
    if(reset_i) begin
      bypass_data_o_28_sv2v_reg <= 1'b0;
      bypass_data_o_27_sv2v_reg <= 1'b0;
      bypass_data_o_26_sv2v_reg <= 1'b0;
      bypass_data_o_25_sv2v_reg <= 1'b0;
      bypass_data_o_24_sv2v_reg <= 1'b0;
      bypass_data_o_23_sv2v_reg <= 1'b0;
      bypass_data_o_22_sv2v_reg <= 1'b0;
      bypass_data_o_21_sv2v_reg <= 1'b0;
      bypass_data_o_20_sv2v_reg <= 1'b0;
      bypass_data_o_19_sv2v_reg <= 1'b0;
      bypass_data_o_18_sv2v_reg <= 1'b0;
      bypass_data_o_17_sv2v_reg <= 1'b0;
      bypass_data_o_16_sv2v_reg <= 1'b0;
      bypass_data_o_15_sv2v_reg <= 1'b0;
      bypass_data_o_14_sv2v_reg <= 1'b0;
      bypass_data_o_13_sv2v_reg <= 1'b0;
      bypass_data_o_12_sv2v_reg <= 1'b0;
      bypass_data_o_11_sv2v_reg <= 1'b0;
      bypass_data_o_10_sv2v_reg <= 1'b0;
      bypass_data_o_9_sv2v_reg <= 1'b0;
      bypass_data_o_8_sv2v_reg <= 1'b0;
      bypass_data_o_7_sv2v_reg <= 1'b0;
      bypass_data_o_6_sv2v_reg <= 1'b0;
      bypass_data_o_5_sv2v_reg <= 1'b0;
      bypass_data_o_4_sv2v_reg <= 1'b0;
      bypass_data_o_3_sv2v_reg <= 1'b0;
      bypass_data_o_2_sv2v_reg <= 1'b0;
      bypass_data_o_1_sv2v_reg <= 1'b0;
      bypass_data_o_0_sv2v_reg <= 1'b0;
      bypass_mask_o_15_sv2v_reg <= 1'b0;
      bypass_mask_o_14_sv2v_reg <= 1'b0;
      bypass_mask_o_13_sv2v_reg <= 1'b0;
      bypass_mask_o_12_sv2v_reg <= 1'b0;
      bypass_mask_o_11_sv2v_reg <= 1'b0;
      bypass_mask_o_10_sv2v_reg <= 1'b0;
      bypass_mask_o_9_sv2v_reg <= 1'b0;
      bypass_mask_o_8_sv2v_reg <= 1'b0;
      bypass_mask_o_7_sv2v_reg <= 1'b0;
      bypass_mask_o_6_sv2v_reg <= 1'b0;
      bypass_mask_o_5_sv2v_reg <= 1'b0;
      bypass_mask_o_4_sv2v_reg <= 1'b0;
      bypass_mask_o_3_sv2v_reg <= 1'b0;
      bypass_mask_o_2_sv2v_reg <= 1'b0;
      bypass_mask_o_1_sv2v_reg <= 1'b0;
    end else if(N3) begin
      bypass_data_o_28_sv2v_reg <= bypass_data_n[28];
      bypass_data_o_27_sv2v_reg <= bypass_data_n[27];
      bypass_data_o_26_sv2v_reg <= bypass_data_n[26];
      bypass_data_o_25_sv2v_reg <= bypass_data_n[25];
      bypass_data_o_24_sv2v_reg <= bypass_data_n[24];
      bypass_data_o_23_sv2v_reg <= bypass_data_n[23];
      bypass_data_o_22_sv2v_reg <= bypass_data_n[22];
      bypass_data_o_21_sv2v_reg <= bypass_data_n[21];
      bypass_data_o_20_sv2v_reg <= bypass_data_n[20];
      bypass_data_o_19_sv2v_reg <= bypass_data_n[19];
      bypass_data_o_18_sv2v_reg <= bypass_data_n[18];
      bypass_data_o_17_sv2v_reg <= bypass_data_n[17];
      bypass_data_o_16_sv2v_reg <= bypass_data_n[16];
      bypass_data_o_15_sv2v_reg <= bypass_data_n[15];
      bypass_data_o_14_sv2v_reg <= bypass_data_n[14];
      bypass_data_o_13_sv2v_reg <= bypass_data_n[13];
      bypass_data_o_12_sv2v_reg <= bypass_data_n[12];
      bypass_data_o_11_sv2v_reg <= bypass_data_n[11];
      bypass_data_o_10_sv2v_reg <= bypass_data_n[10];
      bypass_data_o_9_sv2v_reg <= bypass_data_n[9];
      bypass_data_o_8_sv2v_reg <= bypass_data_n[8];
      bypass_data_o_7_sv2v_reg <= bypass_data_n[7];
      bypass_data_o_6_sv2v_reg <= bypass_data_n[6];
      bypass_data_o_5_sv2v_reg <= bypass_data_n[5];
      bypass_data_o_4_sv2v_reg <= bypass_data_n[4];
      bypass_data_o_3_sv2v_reg <= bypass_data_n[3];
      bypass_data_o_2_sv2v_reg <= bypass_data_n[2];
      bypass_data_o_1_sv2v_reg <= bypass_data_n[1];
      bypass_data_o_0_sv2v_reg <= bypass_data_n[0];
      bypass_mask_o_15_sv2v_reg <= bypass_mask_n[15];
      bypass_mask_o_14_sv2v_reg <= bypass_mask_n[14];
      bypass_mask_o_13_sv2v_reg <= bypass_mask_n[13];
      bypass_mask_o_12_sv2v_reg <= bypass_mask_n[12];
      bypass_mask_o_11_sv2v_reg <= bypass_mask_n[11];
      bypass_mask_o_10_sv2v_reg <= bypass_mask_n[10];
      bypass_mask_o_9_sv2v_reg <= bypass_mask_n[9];
      bypass_mask_o_8_sv2v_reg <= bypass_mask_n[8];
      bypass_mask_o_7_sv2v_reg <= bypass_mask_n[7];
      bypass_mask_o_6_sv2v_reg <= bypass_mask_n[6];
      bypass_mask_o_5_sv2v_reg <= bypass_mask_n[5];
      bypass_mask_o_4_sv2v_reg <= bypass_mask_n[4];
      bypass_mask_o_3_sv2v_reg <= bypass_mask_n[3];
      bypass_mask_o_2_sv2v_reg <= bypass_mask_n[2];
      bypass_mask_o_1_sv2v_reg <= bypass_mask_n[1];
    end 
  end


endmodule



module bsg_decode_00000001
(
  i,
  o
);

  input [0:0] i;
  output [0:0] o;
  wire [0:0] o;
  assign o[0] = 1'b1;

endmodule



module bsg_mux_00000080_00000004
(
  data_i,
  sel_i,
  data_o
);

  input [511:0] data_i;
  input [1:0] sel_i;
  output [127:0] data_o;
  wire [127:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[127] = (N2)? data_i[127] : 
                       (N4)? data_i[255] : 
                       (N3)? data_i[383] : 
                       (N5)? data_i[511] : 1'b0;
  assign data_o[126] = (N2)? data_i[126] : 
                       (N4)? data_i[254] : 
                       (N3)? data_i[382] : 
                       (N5)? data_i[510] : 1'b0;
  assign data_o[125] = (N2)? data_i[125] : 
                       (N4)? data_i[253] : 
                       (N3)? data_i[381] : 
                       (N5)? data_i[509] : 1'b0;
  assign data_o[124] = (N2)? data_i[124] : 
                       (N4)? data_i[252] : 
                       (N3)? data_i[380] : 
                       (N5)? data_i[508] : 1'b0;
  assign data_o[123] = (N2)? data_i[123] : 
                       (N4)? data_i[251] : 
                       (N3)? data_i[379] : 
                       (N5)? data_i[507] : 1'b0;
  assign data_o[122] = (N2)? data_i[122] : 
                       (N4)? data_i[250] : 
                       (N3)? data_i[378] : 
                       (N5)? data_i[506] : 1'b0;
  assign data_o[121] = (N2)? data_i[121] : 
                       (N4)? data_i[249] : 
                       (N3)? data_i[377] : 
                       (N5)? data_i[505] : 1'b0;
  assign data_o[120] = (N2)? data_i[120] : 
                       (N4)? data_i[248] : 
                       (N3)? data_i[376] : 
                       (N5)? data_i[504] : 1'b0;
  assign data_o[119] = (N2)? data_i[119] : 
                       (N4)? data_i[247] : 
                       (N3)? data_i[375] : 
                       (N5)? data_i[503] : 1'b0;
  assign data_o[118] = (N2)? data_i[118] : 
                       (N4)? data_i[246] : 
                       (N3)? data_i[374] : 
                       (N5)? data_i[502] : 1'b0;
  assign data_o[117] = (N2)? data_i[117] : 
                       (N4)? data_i[245] : 
                       (N3)? data_i[373] : 
                       (N5)? data_i[501] : 1'b0;
  assign data_o[116] = (N2)? data_i[116] : 
                       (N4)? data_i[244] : 
                       (N3)? data_i[372] : 
                       (N5)? data_i[500] : 1'b0;
  assign data_o[115] = (N2)? data_i[115] : 
                       (N4)? data_i[243] : 
                       (N3)? data_i[371] : 
                       (N5)? data_i[499] : 1'b0;
  assign data_o[114] = (N2)? data_i[114] : 
                       (N4)? data_i[242] : 
                       (N3)? data_i[370] : 
                       (N5)? data_i[498] : 1'b0;
  assign data_o[113] = (N2)? data_i[113] : 
                       (N4)? data_i[241] : 
                       (N3)? data_i[369] : 
                       (N5)? data_i[497] : 1'b0;
  assign data_o[112] = (N2)? data_i[112] : 
                       (N4)? data_i[240] : 
                       (N3)? data_i[368] : 
                       (N5)? data_i[496] : 1'b0;
  assign data_o[111] = (N2)? data_i[111] : 
                       (N4)? data_i[239] : 
                       (N3)? data_i[367] : 
                       (N5)? data_i[495] : 1'b0;
  assign data_o[110] = (N2)? data_i[110] : 
                       (N4)? data_i[238] : 
                       (N3)? data_i[366] : 
                       (N5)? data_i[494] : 1'b0;
  assign data_o[109] = (N2)? data_i[109] : 
                       (N4)? data_i[237] : 
                       (N3)? data_i[365] : 
                       (N5)? data_i[493] : 1'b0;
  assign data_o[108] = (N2)? data_i[108] : 
                       (N4)? data_i[236] : 
                       (N3)? data_i[364] : 
                       (N5)? data_i[492] : 1'b0;
  assign data_o[107] = (N2)? data_i[107] : 
                       (N4)? data_i[235] : 
                       (N3)? data_i[363] : 
                       (N5)? data_i[491] : 1'b0;
  assign data_o[106] = (N2)? data_i[106] : 
                       (N4)? data_i[234] : 
                       (N3)? data_i[362] : 
                       (N5)? data_i[490] : 1'b0;
  assign data_o[105] = (N2)? data_i[105] : 
                       (N4)? data_i[233] : 
                       (N3)? data_i[361] : 
                       (N5)? data_i[489] : 1'b0;
  assign data_o[104] = (N2)? data_i[104] : 
                       (N4)? data_i[232] : 
                       (N3)? data_i[360] : 
                       (N5)? data_i[488] : 1'b0;
  assign data_o[103] = (N2)? data_i[103] : 
                       (N4)? data_i[231] : 
                       (N3)? data_i[359] : 
                       (N5)? data_i[487] : 1'b0;
  assign data_o[102] = (N2)? data_i[102] : 
                       (N4)? data_i[230] : 
                       (N3)? data_i[358] : 
                       (N5)? data_i[486] : 1'b0;
  assign data_o[101] = (N2)? data_i[101] : 
                       (N4)? data_i[229] : 
                       (N3)? data_i[357] : 
                       (N5)? data_i[485] : 1'b0;
  assign data_o[100] = (N2)? data_i[100] : 
                       (N4)? data_i[228] : 
                       (N3)? data_i[356] : 
                       (N5)? data_i[484] : 1'b0;
  assign data_o[99] = (N2)? data_i[99] : 
                      (N4)? data_i[227] : 
                      (N3)? data_i[355] : 
                      (N5)? data_i[483] : 1'b0;
  assign data_o[98] = (N2)? data_i[98] : 
                      (N4)? data_i[226] : 
                      (N3)? data_i[354] : 
                      (N5)? data_i[482] : 1'b0;
  assign data_o[97] = (N2)? data_i[97] : 
                      (N4)? data_i[225] : 
                      (N3)? data_i[353] : 
                      (N5)? data_i[481] : 1'b0;
  assign data_o[96] = (N2)? data_i[96] : 
                      (N4)? data_i[224] : 
                      (N3)? data_i[352] : 
                      (N5)? data_i[480] : 1'b0;
  assign data_o[95] = (N2)? data_i[95] : 
                      (N4)? data_i[223] : 
                      (N3)? data_i[351] : 
                      (N5)? data_i[479] : 1'b0;
  assign data_o[94] = (N2)? data_i[94] : 
                      (N4)? data_i[222] : 
                      (N3)? data_i[350] : 
                      (N5)? data_i[478] : 1'b0;
  assign data_o[93] = (N2)? data_i[93] : 
                      (N4)? data_i[221] : 
                      (N3)? data_i[349] : 
                      (N5)? data_i[477] : 1'b0;
  assign data_o[92] = (N2)? data_i[92] : 
                      (N4)? data_i[220] : 
                      (N3)? data_i[348] : 
                      (N5)? data_i[476] : 1'b0;
  assign data_o[91] = (N2)? data_i[91] : 
                      (N4)? data_i[219] : 
                      (N3)? data_i[347] : 
                      (N5)? data_i[475] : 1'b0;
  assign data_o[90] = (N2)? data_i[90] : 
                      (N4)? data_i[218] : 
                      (N3)? data_i[346] : 
                      (N5)? data_i[474] : 1'b0;
  assign data_o[89] = (N2)? data_i[89] : 
                      (N4)? data_i[217] : 
                      (N3)? data_i[345] : 
                      (N5)? data_i[473] : 1'b0;
  assign data_o[88] = (N2)? data_i[88] : 
                      (N4)? data_i[216] : 
                      (N3)? data_i[344] : 
                      (N5)? data_i[472] : 1'b0;
  assign data_o[87] = (N2)? data_i[87] : 
                      (N4)? data_i[215] : 
                      (N3)? data_i[343] : 
                      (N5)? data_i[471] : 1'b0;
  assign data_o[86] = (N2)? data_i[86] : 
                      (N4)? data_i[214] : 
                      (N3)? data_i[342] : 
                      (N5)? data_i[470] : 1'b0;
  assign data_o[85] = (N2)? data_i[85] : 
                      (N4)? data_i[213] : 
                      (N3)? data_i[341] : 
                      (N5)? data_i[469] : 1'b0;
  assign data_o[84] = (N2)? data_i[84] : 
                      (N4)? data_i[212] : 
                      (N3)? data_i[340] : 
                      (N5)? data_i[468] : 1'b0;
  assign data_o[83] = (N2)? data_i[83] : 
                      (N4)? data_i[211] : 
                      (N3)? data_i[339] : 
                      (N5)? data_i[467] : 1'b0;
  assign data_o[82] = (N2)? data_i[82] : 
                      (N4)? data_i[210] : 
                      (N3)? data_i[338] : 
                      (N5)? data_i[466] : 1'b0;
  assign data_o[81] = (N2)? data_i[81] : 
                      (N4)? data_i[209] : 
                      (N3)? data_i[337] : 
                      (N5)? data_i[465] : 1'b0;
  assign data_o[80] = (N2)? data_i[80] : 
                      (N4)? data_i[208] : 
                      (N3)? data_i[336] : 
                      (N5)? data_i[464] : 1'b0;
  assign data_o[79] = (N2)? data_i[79] : 
                      (N4)? data_i[207] : 
                      (N3)? data_i[335] : 
                      (N5)? data_i[463] : 1'b0;
  assign data_o[78] = (N2)? data_i[78] : 
                      (N4)? data_i[206] : 
                      (N3)? data_i[334] : 
                      (N5)? data_i[462] : 1'b0;
  assign data_o[77] = (N2)? data_i[77] : 
                      (N4)? data_i[205] : 
                      (N3)? data_i[333] : 
                      (N5)? data_i[461] : 1'b0;
  assign data_o[76] = (N2)? data_i[76] : 
                      (N4)? data_i[204] : 
                      (N3)? data_i[332] : 
                      (N5)? data_i[460] : 1'b0;
  assign data_o[75] = (N2)? data_i[75] : 
                      (N4)? data_i[203] : 
                      (N3)? data_i[331] : 
                      (N5)? data_i[459] : 1'b0;
  assign data_o[74] = (N2)? data_i[74] : 
                      (N4)? data_i[202] : 
                      (N3)? data_i[330] : 
                      (N5)? data_i[458] : 1'b0;
  assign data_o[73] = (N2)? data_i[73] : 
                      (N4)? data_i[201] : 
                      (N3)? data_i[329] : 
                      (N5)? data_i[457] : 1'b0;
  assign data_o[72] = (N2)? data_i[72] : 
                      (N4)? data_i[200] : 
                      (N3)? data_i[328] : 
                      (N5)? data_i[456] : 1'b0;
  assign data_o[71] = (N2)? data_i[71] : 
                      (N4)? data_i[199] : 
                      (N3)? data_i[327] : 
                      (N5)? data_i[455] : 1'b0;
  assign data_o[70] = (N2)? data_i[70] : 
                      (N4)? data_i[198] : 
                      (N3)? data_i[326] : 
                      (N5)? data_i[454] : 1'b0;
  assign data_o[69] = (N2)? data_i[69] : 
                      (N4)? data_i[197] : 
                      (N3)? data_i[325] : 
                      (N5)? data_i[453] : 1'b0;
  assign data_o[68] = (N2)? data_i[68] : 
                      (N4)? data_i[196] : 
                      (N3)? data_i[324] : 
                      (N5)? data_i[452] : 1'b0;
  assign data_o[67] = (N2)? data_i[67] : 
                      (N4)? data_i[195] : 
                      (N3)? data_i[323] : 
                      (N5)? data_i[451] : 1'b0;
  assign data_o[66] = (N2)? data_i[66] : 
                      (N4)? data_i[194] : 
                      (N3)? data_i[322] : 
                      (N5)? data_i[450] : 1'b0;
  assign data_o[65] = (N2)? data_i[65] : 
                      (N4)? data_i[193] : 
                      (N3)? data_i[321] : 
                      (N5)? data_i[449] : 1'b0;
  assign data_o[64] = (N2)? data_i[64] : 
                      (N4)? data_i[192] : 
                      (N3)? data_i[320] : 
                      (N5)? data_i[448] : 1'b0;
  assign data_o[63] = (N2)? data_i[63] : 
                      (N4)? data_i[191] : 
                      (N3)? data_i[319] : 
                      (N5)? data_i[447] : 1'b0;
  assign data_o[62] = (N2)? data_i[62] : 
                      (N4)? data_i[190] : 
                      (N3)? data_i[318] : 
                      (N5)? data_i[446] : 1'b0;
  assign data_o[61] = (N2)? data_i[61] : 
                      (N4)? data_i[189] : 
                      (N3)? data_i[317] : 
                      (N5)? data_i[445] : 1'b0;
  assign data_o[60] = (N2)? data_i[60] : 
                      (N4)? data_i[188] : 
                      (N3)? data_i[316] : 
                      (N5)? data_i[444] : 1'b0;
  assign data_o[59] = (N2)? data_i[59] : 
                      (N4)? data_i[187] : 
                      (N3)? data_i[315] : 
                      (N5)? data_i[443] : 1'b0;
  assign data_o[58] = (N2)? data_i[58] : 
                      (N4)? data_i[186] : 
                      (N3)? data_i[314] : 
                      (N5)? data_i[442] : 1'b0;
  assign data_o[57] = (N2)? data_i[57] : 
                      (N4)? data_i[185] : 
                      (N3)? data_i[313] : 
                      (N5)? data_i[441] : 1'b0;
  assign data_o[56] = (N2)? data_i[56] : 
                      (N4)? data_i[184] : 
                      (N3)? data_i[312] : 
                      (N5)? data_i[440] : 1'b0;
  assign data_o[55] = (N2)? data_i[55] : 
                      (N4)? data_i[183] : 
                      (N3)? data_i[311] : 
                      (N5)? data_i[439] : 1'b0;
  assign data_o[54] = (N2)? data_i[54] : 
                      (N4)? data_i[182] : 
                      (N3)? data_i[310] : 
                      (N5)? data_i[438] : 1'b0;
  assign data_o[53] = (N2)? data_i[53] : 
                      (N4)? data_i[181] : 
                      (N3)? data_i[309] : 
                      (N5)? data_i[437] : 1'b0;
  assign data_o[52] = (N2)? data_i[52] : 
                      (N4)? data_i[180] : 
                      (N3)? data_i[308] : 
                      (N5)? data_i[436] : 1'b0;
  assign data_o[51] = (N2)? data_i[51] : 
                      (N4)? data_i[179] : 
                      (N3)? data_i[307] : 
                      (N5)? data_i[435] : 1'b0;
  assign data_o[50] = (N2)? data_i[50] : 
                      (N4)? data_i[178] : 
                      (N3)? data_i[306] : 
                      (N5)? data_i[434] : 1'b0;
  assign data_o[49] = (N2)? data_i[49] : 
                      (N4)? data_i[177] : 
                      (N3)? data_i[305] : 
                      (N5)? data_i[433] : 1'b0;
  assign data_o[48] = (N2)? data_i[48] : 
                      (N4)? data_i[176] : 
                      (N3)? data_i[304] : 
                      (N5)? data_i[432] : 1'b0;
  assign data_o[47] = (N2)? data_i[47] : 
                      (N4)? data_i[175] : 
                      (N3)? data_i[303] : 
                      (N5)? data_i[431] : 1'b0;
  assign data_o[46] = (N2)? data_i[46] : 
                      (N4)? data_i[174] : 
                      (N3)? data_i[302] : 
                      (N5)? data_i[430] : 1'b0;
  assign data_o[45] = (N2)? data_i[45] : 
                      (N4)? data_i[173] : 
                      (N3)? data_i[301] : 
                      (N5)? data_i[429] : 1'b0;
  assign data_o[44] = (N2)? data_i[44] : 
                      (N4)? data_i[172] : 
                      (N3)? data_i[300] : 
                      (N5)? data_i[428] : 1'b0;
  assign data_o[43] = (N2)? data_i[43] : 
                      (N4)? data_i[171] : 
                      (N3)? data_i[299] : 
                      (N5)? data_i[427] : 1'b0;
  assign data_o[42] = (N2)? data_i[42] : 
                      (N4)? data_i[170] : 
                      (N3)? data_i[298] : 
                      (N5)? data_i[426] : 1'b0;
  assign data_o[41] = (N2)? data_i[41] : 
                      (N4)? data_i[169] : 
                      (N3)? data_i[297] : 
                      (N5)? data_i[425] : 1'b0;
  assign data_o[40] = (N2)? data_i[40] : 
                      (N4)? data_i[168] : 
                      (N3)? data_i[296] : 
                      (N5)? data_i[424] : 1'b0;
  assign data_o[39] = (N2)? data_i[39] : 
                      (N4)? data_i[167] : 
                      (N3)? data_i[295] : 
                      (N5)? data_i[423] : 1'b0;
  assign data_o[38] = (N2)? data_i[38] : 
                      (N4)? data_i[166] : 
                      (N3)? data_i[294] : 
                      (N5)? data_i[422] : 1'b0;
  assign data_o[37] = (N2)? data_i[37] : 
                      (N4)? data_i[165] : 
                      (N3)? data_i[293] : 
                      (N5)? data_i[421] : 1'b0;
  assign data_o[36] = (N2)? data_i[36] : 
                      (N4)? data_i[164] : 
                      (N3)? data_i[292] : 
                      (N5)? data_i[420] : 1'b0;
  assign data_o[35] = (N2)? data_i[35] : 
                      (N4)? data_i[163] : 
                      (N3)? data_i[291] : 
                      (N5)? data_i[419] : 1'b0;
  assign data_o[34] = (N2)? data_i[34] : 
                      (N4)? data_i[162] : 
                      (N3)? data_i[290] : 
                      (N5)? data_i[418] : 1'b0;
  assign data_o[33] = (N2)? data_i[33] : 
                      (N4)? data_i[161] : 
                      (N3)? data_i[289] : 
                      (N5)? data_i[417] : 1'b0;
  assign data_o[32] = (N2)? data_i[32] : 
                      (N4)? data_i[160] : 
                      (N3)? data_i[288] : 
                      (N5)? data_i[416] : 1'b0;
  assign data_o[31] = (N2)? data_i[31] : 
                      (N4)? data_i[159] : 
                      (N3)? data_i[287] : 
                      (N5)? data_i[415] : 1'b0;
  assign data_o[30] = (N2)? data_i[30] : 
                      (N4)? data_i[158] : 
                      (N3)? data_i[286] : 
                      (N5)? data_i[414] : 1'b0;
  assign data_o[29] = (N2)? data_i[29] : 
                      (N4)? data_i[157] : 
                      (N3)? data_i[285] : 
                      (N5)? data_i[413] : 1'b0;
  assign data_o[28] = (N2)? data_i[28] : 
                      (N4)? data_i[156] : 
                      (N3)? data_i[284] : 
                      (N5)? data_i[412] : 1'b0;
  assign data_o[27] = (N2)? data_i[27] : 
                      (N4)? data_i[155] : 
                      (N3)? data_i[283] : 
                      (N5)? data_i[411] : 1'b0;
  assign data_o[26] = (N2)? data_i[26] : 
                      (N4)? data_i[154] : 
                      (N3)? data_i[282] : 
                      (N5)? data_i[410] : 1'b0;
  assign data_o[25] = (N2)? data_i[25] : 
                      (N4)? data_i[153] : 
                      (N3)? data_i[281] : 
                      (N5)? data_i[409] : 1'b0;
  assign data_o[24] = (N2)? data_i[24] : 
                      (N4)? data_i[152] : 
                      (N3)? data_i[280] : 
                      (N5)? data_i[408] : 1'b0;
  assign data_o[23] = (N2)? data_i[23] : 
                      (N4)? data_i[151] : 
                      (N3)? data_i[279] : 
                      (N5)? data_i[407] : 1'b0;
  assign data_o[22] = (N2)? data_i[22] : 
                      (N4)? data_i[150] : 
                      (N3)? data_i[278] : 
                      (N5)? data_i[406] : 1'b0;
  assign data_o[21] = (N2)? data_i[21] : 
                      (N4)? data_i[149] : 
                      (N3)? data_i[277] : 
                      (N5)? data_i[405] : 1'b0;
  assign data_o[20] = (N2)? data_i[20] : 
                      (N4)? data_i[148] : 
                      (N3)? data_i[276] : 
                      (N5)? data_i[404] : 1'b0;
  assign data_o[19] = (N2)? data_i[19] : 
                      (N4)? data_i[147] : 
                      (N3)? data_i[275] : 
                      (N5)? data_i[403] : 1'b0;
  assign data_o[18] = (N2)? data_i[18] : 
                      (N4)? data_i[146] : 
                      (N3)? data_i[274] : 
                      (N5)? data_i[402] : 1'b0;
  assign data_o[17] = (N2)? data_i[17] : 
                      (N4)? data_i[145] : 
                      (N3)? data_i[273] : 
                      (N5)? data_i[401] : 1'b0;
  assign data_o[16] = (N2)? data_i[16] : 
                      (N4)? data_i[144] : 
                      (N3)? data_i[272] : 
                      (N5)? data_i[400] : 1'b0;
  assign data_o[15] = (N2)? data_i[15] : 
                      (N4)? data_i[143] : 
                      (N3)? data_i[271] : 
                      (N5)? data_i[399] : 1'b0;
  assign data_o[14] = (N2)? data_i[14] : 
                      (N4)? data_i[142] : 
                      (N3)? data_i[270] : 
                      (N5)? data_i[398] : 1'b0;
  assign data_o[13] = (N2)? data_i[13] : 
                      (N4)? data_i[141] : 
                      (N3)? data_i[269] : 
                      (N5)? data_i[397] : 1'b0;
  assign data_o[12] = (N2)? data_i[12] : 
                      (N4)? data_i[140] : 
                      (N3)? data_i[268] : 
                      (N5)? data_i[396] : 1'b0;
  assign data_o[11] = (N2)? data_i[11] : 
                      (N4)? data_i[139] : 
                      (N3)? data_i[267] : 
                      (N5)? data_i[395] : 1'b0;
  assign data_o[10] = (N2)? data_i[10] : 
                      (N4)? data_i[138] : 
                      (N3)? data_i[266] : 
                      (N5)? data_i[394] : 1'b0;
  assign data_o[9] = (N2)? data_i[9] : 
                     (N4)? data_i[137] : 
                     (N3)? data_i[265] : 
                     (N5)? data_i[393] : 1'b0;
  assign data_o[8] = (N2)? data_i[8] : 
                     (N4)? data_i[136] : 
                     (N3)? data_i[264] : 
                     (N5)? data_i[392] : 1'b0;
  assign data_o[7] = (N2)? data_i[7] : 
                     (N4)? data_i[135] : 
                     (N3)? data_i[263] : 
                     (N5)? data_i[391] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] : 
                     (N4)? data_i[134] : 
                     (N3)? data_i[262] : 
                     (N5)? data_i[390] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] : 
                     (N4)? data_i[133] : 
                     (N3)? data_i[261] : 
                     (N5)? data_i[389] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] : 
                     (N4)? data_i[132] : 
                     (N3)? data_i[260] : 
                     (N5)? data_i[388] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] : 
                     (N4)? data_i[131] : 
                     (N3)? data_i[259] : 
                     (N5)? data_i[387] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] : 
                     (N4)? data_i[130] : 
                     (N3)? data_i[258] : 
                     (N5)? data_i[386] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N4)? data_i[129] : 
                     (N3)? data_i[257] : 
                     (N5)? data_i[385] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[128] : 
                     (N3)? data_i[256] : 
                     (N5)? data_i[384] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_mux_00000010_00000004
(
  data_i,
  sel_i,
  data_o
);

  input [63:0] data_i;
  input [1:0] sel_i;
  output [15:0] data_o;
  wire [15:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[15] = (N2)? data_i[15] : 
                      (N4)? data_i[31] : 
                      (N3)? data_i[47] : 
                      (N5)? data_i[63] : 1'b0;
  assign data_o[14] = (N2)? data_i[14] : 
                      (N4)? data_i[30] : 
                      (N3)? data_i[46] : 
                      (N5)? data_i[62] : 1'b0;
  assign data_o[13] = (N2)? data_i[13] : 
                      (N4)? data_i[29] : 
                      (N3)? data_i[45] : 
                      (N5)? data_i[61] : 1'b0;
  assign data_o[12] = (N2)? data_i[12] : 
                      (N4)? data_i[28] : 
                      (N3)? data_i[44] : 
                      (N5)? data_i[60] : 1'b0;
  assign data_o[11] = (N2)? data_i[11] : 
                      (N4)? data_i[27] : 
                      (N3)? data_i[43] : 
                      (N5)? data_i[59] : 1'b0;
  assign data_o[10] = (N2)? data_i[10] : 
                      (N4)? data_i[26] : 
                      (N3)? data_i[42] : 
                      (N5)? data_i[58] : 1'b0;
  assign data_o[9] = (N2)? data_i[9] : 
                     (N4)? data_i[25] : 
                     (N3)? data_i[41] : 
                     (N5)? data_i[57] : 1'b0;
  assign data_o[8] = (N2)? data_i[8] : 
                     (N4)? data_i[24] : 
                     (N3)? data_i[40] : 
                     (N5)? data_i[56] : 1'b0;
  assign data_o[7] = (N2)? data_i[7] : 
                     (N4)? data_i[23] : 
                     (N3)? data_i[39] : 
                     (N5)? data_i[55] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] : 
                     (N4)? data_i[22] : 
                     (N3)? data_i[38] : 
                     (N5)? data_i[54] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] : 
                     (N4)? data_i[21] : 
                     (N3)? data_i[37] : 
                     (N5)? data_i[53] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] : 
                     (N4)? data_i[20] : 
                     (N3)? data_i[36] : 
                     (N5)? data_i[52] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] : 
                     (N4)? data_i[19] : 
                     (N3)? data_i[35] : 
                     (N5)? data_i[51] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] : 
                     (N4)? data_i[18] : 
                     (N3)? data_i[34] : 
                     (N5)? data_i[50] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N4)? data_i[17] : 
                     (N3)? data_i[33] : 
                     (N5)? data_i[49] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[16] : 
                     (N3)? data_i[32] : 
                     (N5)? data_i[48] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_decode_00000010
(
  i,
  o
);

  input [3:0] i;
  output [15:0] o;
  wire [15:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_decode_00000004
(
  i,
  o
);

  input [1:0] i;
  output [3:0] o;
  wire [3:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_cache_buffer_queue_00000024
(
  clk_i,
  reset_i,
  v_i,
  data_i,
  v_o,
  data_o,
  yumi_i,
  el0_valid_o,
  el1_valid_o,
  el0_snoop_o,
  el1_snoop_o,
  empty_o,
  full_o
);

  input [35:0] data_i;
  output [35:0] data_o;
  output [35:0] el0_snoop_o;
  output [35:0] el1_snoop_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output v_o;
  output el0_valid_o;
  output el1_valid_o;
  output empty_o;
  output full_o;
  wire [35:0] data_o,el0_snoop_o,el1_snoop_o;
  wire v_o,el0_valid_o,el1_valid_o,empty_o,full_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,
  N11,N12,N13,N14,N15,el0_enable,el1_enable,mux0_sel,mux1_sel,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62;
  wire [1:0] num_els_r;
  reg num_els_r_1_sv2v_reg,num_els_r_0_sv2v_reg,el0_snoop_o_35_sv2v_reg,
  el0_snoop_o_34_sv2v_reg,el0_snoop_o_33_sv2v_reg,el0_snoop_o_32_sv2v_reg,
  el0_snoop_o_31_sv2v_reg,el0_snoop_o_30_sv2v_reg,el0_snoop_o_29_sv2v_reg,el0_snoop_o_28_sv2v_reg,
  el0_snoop_o_27_sv2v_reg,el0_snoop_o_26_sv2v_reg,el0_snoop_o_25_sv2v_reg,
  el0_snoop_o_24_sv2v_reg,el0_snoop_o_23_sv2v_reg,el0_snoop_o_22_sv2v_reg,
  el0_snoop_o_21_sv2v_reg,el0_snoop_o_20_sv2v_reg,el0_snoop_o_19_sv2v_reg,el0_snoop_o_18_sv2v_reg,
  el0_snoop_o_17_sv2v_reg,el0_snoop_o_16_sv2v_reg,el0_snoop_o_15_sv2v_reg,
  el0_snoop_o_14_sv2v_reg,el0_snoop_o_13_sv2v_reg,el0_snoop_o_12_sv2v_reg,
  el0_snoop_o_11_sv2v_reg,el0_snoop_o_10_sv2v_reg,el0_snoop_o_9_sv2v_reg,el0_snoop_o_8_sv2v_reg,
  el0_snoop_o_7_sv2v_reg,el0_snoop_o_6_sv2v_reg,el0_snoop_o_5_sv2v_reg,
  el0_snoop_o_4_sv2v_reg,el0_snoop_o_3_sv2v_reg,el0_snoop_o_2_sv2v_reg,el0_snoop_o_1_sv2v_reg,
  el0_snoop_o_0_sv2v_reg,el1_snoop_o_35_sv2v_reg,el1_snoop_o_34_sv2v_reg,
  el1_snoop_o_33_sv2v_reg,el1_snoop_o_32_sv2v_reg,el1_snoop_o_31_sv2v_reg,el1_snoop_o_30_sv2v_reg,
  el1_snoop_o_29_sv2v_reg,el1_snoop_o_28_sv2v_reg,el1_snoop_o_27_sv2v_reg,
  el1_snoop_o_26_sv2v_reg,el1_snoop_o_25_sv2v_reg,el1_snoop_o_24_sv2v_reg,
  el1_snoop_o_23_sv2v_reg,el1_snoop_o_22_sv2v_reg,el1_snoop_o_21_sv2v_reg,el1_snoop_o_20_sv2v_reg,
  el1_snoop_o_19_sv2v_reg,el1_snoop_o_18_sv2v_reg,el1_snoop_o_17_sv2v_reg,
  el1_snoop_o_16_sv2v_reg,el1_snoop_o_15_sv2v_reg,el1_snoop_o_14_sv2v_reg,
  el1_snoop_o_13_sv2v_reg,el1_snoop_o_12_sv2v_reg,el1_snoop_o_11_sv2v_reg,el1_snoop_o_10_sv2v_reg,
  el1_snoop_o_9_sv2v_reg,el1_snoop_o_8_sv2v_reg,el1_snoop_o_7_sv2v_reg,
  el1_snoop_o_6_sv2v_reg,el1_snoop_o_5_sv2v_reg,el1_snoop_o_4_sv2v_reg,
  el1_snoop_o_3_sv2v_reg,el1_snoop_o_2_sv2v_reg,el1_snoop_o_1_sv2v_reg,el1_snoop_o_0_sv2v_reg;
  assign num_els_r[1] = num_els_r_1_sv2v_reg;
  assign num_els_r[0] = num_els_r_0_sv2v_reg;
  assign el0_snoop_o[35] = el0_snoop_o_35_sv2v_reg;
  assign el0_snoop_o[34] = el0_snoop_o_34_sv2v_reg;
  assign el0_snoop_o[33] = el0_snoop_o_33_sv2v_reg;
  assign el0_snoop_o[32] = el0_snoop_o_32_sv2v_reg;
  assign el0_snoop_o[31] = el0_snoop_o_31_sv2v_reg;
  assign el0_snoop_o[30] = el0_snoop_o_30_sv2v_reg;
  assign el0_snoop_o[29] = el0_snoop_o_29_sv2v_reg;
  assign el0_snoop_o[28] = el0_snoop_o_28_sv2v_reg;
  assign el0_snoop_o[27] = el0_snoop_o_27_sv2v_reg;
  assign el0_snoop_o[26] = el0_snoop_o_26_sv2v_reg;
  assign el0_snoop_o[25] = el0_snoop_o_25_sv2v_reg;
  assign el0_snoop_o[24] = el0_snoop_o_24_sv2v_reg;
  assign el0_snoop_o[23] = el0_snoop_o_23_sv2v_reg;
  assign el0_snoop_o[22] = el0_snoop_o_22_sv2v_reg;
  assign el0_snoop_o[21] = el0_snoop_o_21_sv2v_reg;
  assign el0_snoop_o[20] = el0_snoop_o_20_sv2v_reg;
  assign el0_snoop_o[19] = el0_snoop_o_19_sv2v_reg;
  assign el0_snoop_o[18] = el0_snoop_o_18_sv2v_reg;
  assign el0_snoop_o[17] = el0_snoop_o_17_sv2v_reg;
  assign el0_snoop_o[16] = el0_snoop_o_16_sv2v_reg;
  assign el0_snoop_o[15] = el0_snoop_o_15_sv2v_reg;
  assign el0_snoop_o[14] = el0_snoop_o_14_sv2v_reg;
  assign el0_snoop_o[13] = el0_snoop_o_13_sv2v_reg;
  assign el0_snoop_o[12] = el0_snoop_o_12_sv2v_reg;
  assign el0_snoop_o[11] = el0_snoop_o_11_sv2v_reg;
  assign el0_snoop_o[10] = el0_snoop_o_10_sv2v_reg;
  assign el0_snoop_o[9] = el0_snoop_o_9_sv2v_reg;
  assign el0_snoop_o[8] = el0_snoop_o_8_sv2v_reg;
  assign el0_snoop_o[7] = el0_snoop_o_7_sv2v_reg;
  assign el0_snoop_o[6] = el0_snoop_o_6_sv2v_reg;
  assign el0_snoop_o[5] = el0_snoop_o_5_sv2v_reg;
  assign el0_snoop_o[4] = el0_snoop_o_4_sv2v_reg;
  assign el0_snoop_o[3] = el0_snoop_o_3_sv2v_reg;
  assign el0_snoop_o[2] = el0_snoop_o_2_sv2v_reg;
  assign el0_snoop_o[1] = el0_snoop_o_1_sv2v_reg;
  assign el0_snoop_o[0] = el0_snoop_o_0_sv2v_reg;
  assign el1_snoop_o[35] = el1_snoop_o_35_sv2v_reg;
  assign el1_snoop_o[34] = el1_snoop_o_34_sv2v_reg;
  assign el1_snoop_o[33] = el1_snoop_o_33_sv2v_reg;
  assign el1_snoop_o[32] = el1_snoop_o_32_sv2v_reg;
  assign el1_snoop_o[31] = el1_snoop_o_31_sv2v_reg;
  assign el1_snoop_o[30] = el1_snoop_o_30_sv2v_reg;
  assign el1_snoop_o[29] = el1_snoop_o_29_sv2v_reg;
  assign el1_snoop_o[28] = el1_snoop_o_28_sv2v_reg;
  assign el1_snoop_o[27] = el1_snoop_o_27_sv2v_reg;
  assign el1_snoop_o[26] = el1_snoop_o_26_sv2v_reg;
  assign el1_snoop_o[25] = el1_snoop_o_25_sv2v_reg;
  assign el1_snoop_o[24] = el1_snoop_o_24_sv2v_reg;
  assign el1_snoop_o[23] = el1_snoop_o_23_sv2v_reg;
  assign el1_snoop_o[22] = el1_snoop_o_22_sv2v_reg;
  assign el1_snoop_o[21] = el1_snoop_o_21_sv2v_reg;
  assign el1_snoop_o[20] = el1_snoop_o_20_sv2v_reg;
  assign el1_snoop_o[19] = el1_snoop_o_19_sv2v_reg;
  assign el1_snoop_o[18] = el1_snoop_o_18_sv2v_reg;
  assign el1_snoop_o[17] = el1_snoop_o_17_sv2v_reg;
  assign el1_snoop_o[16] = el1_snoop_o_16_sv2v_reg;
  assign el1_snoop_o[15] = el1_snoop_o_15_sv2v_reg;
  assign el1_snoop_o[14] = el1_snoop_o_14_sv2v_reg;
  assign el1_snoop_o[13] = el1_snoop_o_13_sv2v_reg;
  assign el1_snoop_o[12] = el1_snoop_o_12_sv2v_reg;
  assign el1_snoop_o[11] = el1_snoop_o_11_sv2v_reg;
  assign el1_snoop_o[10] = el1_snoop_o_10_sv2v_reg;
  assign el1_snoop_o[9] = el1_snoop_o_9_sv2v_reg;
  assign el1_snoop_o[8] = el1_snoop_o_8_sv2v_reg;
  assign el1_snoop_o[7] = el1_snoop_o_7_sv2v_reg;
  assign el1_snoop_o[6] = el1_snoop_o_6_sv2v_reg;
  assign el1_snoop_o[5] = el1_snoop_o_5_sv2v_reg;
  assign el1_snoop_o[4] = el1_snoop_o_4_sv2v_reg;
  assign el1_snoop_o[3] = el1_snoop_o_3_sv2v_reg;
  assign el1_snoop_o[2] = el1_snoop_o_2_sv2v_reg;
  assign el1_snoop_o[1] = el1_snoop_o_1_sv2v_reg;
  assign el1_snoop_o[0] = el1_snoop_o_0_sv2v_reg;
  assign N10 = N8 & N9;
  assign N11 = num_els_r[1] | N9;
  assign N13 = N8 | num_els_r[0];
  assign N15 = num_els_r[1] & num_els_r[0];
  assign { N20, N19 } = num_els_r + v_i;
  assign { N23, N22 } = { N20, N19 } - N21;
  assign v_o = (N0)? v_i : 
               (N1)? 1'b1 : 
               (N2)? 1'b1 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = N10;
  assign N1 = N12;
  assign N2 = N14;
  assign N3 = N15;
  assign empty_o = (N0)? 1'b1 : 
                   (N1)? 1'b0 : 
                   (N2)? 1'b0 : 
                   (N3)? 1'b0 : 1'b0;
  assign full_o = (N0)? 1'b0 : 
                  (N1)? 1'b0 : 
                  (N2)? 1'b1 : 
                  (N3)? 1'b0 : 1'b0;
  assign el0_valid_o = (N0)? 1'b0 : 
                       (N1)? 1'b0 : 
                       (N2)? 1'b1 : 
                       (N3)? 1'b0 : 1'b0;
  assign el1_valid_o = (N0)? 1'b0 : 
                       (N1)? 1'b1 : 
                       (N2)? 1'b1 : 
                       (N3)? 1'b0 : 1'b0;
  assign el0_enable = (N0)? 1'b0 : 
                      (N1)? N16 : 
                      (N2)? N17 : 
                      (N3)? 1'b0 : 1'b0;
  assign el1_enable = (N0)? N16 : 
                      (N1)? N17 : 
                      (N2)? yumi_i : 
                      (N3)? 1'b0 : 1'b0;
  assign mux0_sel = (N0)? 1'b0 : 
                    (N1)? 1'b0 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b0 : 1'b0;
  assign mux1_sel = (N0)? 1'b0 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b0 : 1'b0;
  assign { N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25 } = (N4)? el0_snoop_o : 
                                                                                                                                                                                                  (N5)? data_i : 1'b0;
  assign N4 = mux0_sel;
  assign N5 = N24;
  assign data_o = (N6)? el1_snoop_o : 
                  (N7)? data_i : 1'b0;
  assign N6 = mux1_sel;
  assign N7 = N61;
  assign N8 = ~num_els_r[1];
  assign N9 = ~num_els_r[0];
  assign N12 = ~N11;
  assign N14 = ~N13;
  assign N16 = v_i & N62;
  assign N62 = ~yumi_i;
  assign N17 = v_i & yumi_i;
  assign N18 = ~reset_i;
  assign N21 = v_o & yumi_i;
  assign N24 = ~mux0_sel;
  assign N61 = ~mux1_sel;

  always @(posedge clk_i) begin
    if(reset_i) begin
      num_els_r_1_sv2v_reg <= 1'b0;
      num_els_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      num_els_r_1_sv2v_reg <= N23;
      num_els_r_0_sv2v_reg <= N22;
    end 
    if(el0_enable) begin
      el0_snoop_o_35_sv2v_reg <= data_i[35];
      el0_snoop_o_34_sv2v_reg <= data_i[34];
      el0_snoop_o_33_sv2v_reg <= data_i[33];
      el0_snoop_o_32_sv2v_reg <= data_i[32];
      el0_snoop_o_31_sv2v_reg <= data_i[31];
      el0_snoop_o_30_sv2v_reg <= data_i[30];
      el0_snoop_o_29_sv2v_reg <= data_i[29];
      el0_snoop_o_28_sv2v_reg <= data_i[28];
      el0_snoop_o_27_sv2v_reg <= data_i[27];
      el0_snoop_o_26_sv2v_reg <= data_i[26];
      el0_snoop_o_25_sv2v_reg <= data_i[25];
      el0_snoop_o_24_sv2v_reg <= data_i[24];
      el0_snoop_o_23_sv2v_reg <= data_i[23];
      el0_snoop_o_22_sv2v_reg <= data_i[22];
      el0_snoop_o_21_sv2v_reg <= data_i[21];
      el0_snoop_o_20_sv2v_reg <= data_i[20];
      el0_snoop_o_19_sv2v_reg <= data_i[19];
      el0_snoop_o_18_sv2v_reg <= data_i[18];
      el0_snoop_o_17_sv2v_reg <= data_i[17];
      el0_snoop_o_16_sv2v_reg <= data_i[16];
      el0_snoop_o_15_sv2v_reg <= data_i[15];
      el0_snoop_o_14_sv2v_reg <= data_i[14];
      el0_snoop_o_13_sv2v_reg <= data_i[13];
      el0_snoop_o_12_sv2v_reg <= data_i[12];
      el0_snoop_o_11_sv2v_reg <= data_i[11];
      el0_snoop_o_10_sv2v_reg <= data_i[10];
      el0_snoop_o_9_sv2v_reg <= data_i[9];
      el0_snoop_o_8_sv2v_reg <= data_i[8];
      el0_snoop_o_7_sv2v_reg <= data_i[7];
      el0_snoop_o_6_sv2v_reg <= data_i[6];
      el0_snoop_o_5_sv2v_reg <= data_i[5];
      el0_snoop_o_4_sv2v_reg <= data_i[4];
      el0_snoop_o_3_sv2v_reg <= data_i[3];
      el0_snoop_o_2_sv2v_reg <= data_i[2];
      el0_snoop_o_1_sv2v_reg <= data_i[1];
      el0_snoop_o_0_sv2v_reg <= data_i[0];
    end 
    if(el1_enable) begin
      el1_snoop_o_35_sv2v_reg <= N60;
      el1_snoop_o_34_sv2v_reg <= N59;
      el1_snoop_o_33_sv2v_reg <= N58;
      el1_snoop_o_32_sv2v_reg <= N57;
      el1_snoop_o_31_sv2v_reg <= N56;
      el1_snoop_o_30_sv2v_reg <= N55;
      el1_snoop_o_29_sv2v_reg <= N54;
      el1_snoop_o_28_sv2v_reg <= N53;
      el1_snoop_o_27_sv2v_reg <= N52;
      el1_snoop_o_26_sv2v_reg <= N51;
      el1_snoop_o_25_sv2v_reg <= N50;
      el1_snoop_o_24_sv2v_reg <= N49;
      el1_snoop_o_23_sv2v_reg <= N48;
      el1_snoop_o_22_sv2v_reg <= N47;
      el1_snoop_o_21_sv2v_reg <= N46;
      el1_snoop_o_20_sv2v_reg <= N45;
      el1_snoop_o_19_sv2v_reg <= N44;
      el1_snoop_o_18_sv2v_reg <= N43;
      el1_snoop_o_17_sv2v_reg <= N42;
      el1_snoop_o_16_sv2v_reg <= N41;
      el1_snoop_o_15_sv2v_reg <= N40;
      el1_snoop_o_14_sv2v_reg <= N39;
      el1_snoop_o_13_sv2v_reg <= N38;
      el1_snoop_o_12_sv2v_reg <= N37;
      el1_snoop_o_11_sv2v_reg <= N36;
      el1_snoop_o_10_sv2v_reg <= N35;
      el1_snoop_o_9_sv2v_reg <= N34;
      el1_snoop_o_8_sv2v_reg <= N33;
      el1_snoop_o_7_sv2v_reg <= N32;
      el1_snoop_o_6_sv2v_reg <= N31;
      el1_snoop_o_5_sv2v_reg <= N30;
      el1_snoop_o_4_sv2v_reg <= N29;
      el1_snoop_o_3_sv2v_reg <= N28;
      el1_snoop_o_2_sv2v_reg <= N27;
      el1_snoop_o_1_sv2v_reg <= N26;
      el1_snoop_o_0_sv2v_reg <= N25;
    end 
  end


endmodule



module bsg_cache_tbuf_00000080_00000021_00000008
(
  clk_i,
  reset_i,
  addr_i,
  way_i,
  v_i,
  addr_o,
  way_o,
  v_o,
  yumi_i,
  empty_o,
  full_o,
  bypass_addr_i,
  bypass_v_i,
  bypass_track_o
);

  input [32:0] addr_i;
  input [2:0] way_i;
  output [32:0] addr_o;
  output [2:0] way_o;
  input [32:0] bypass_addr_i;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input bypass_v_i;
  output v_o;
  output empty_o;
  output full_o;
  output bypass_track_o;
  wire [32:0] addr_o,el1_addr,el0_addr;
  wire [2:0] way_o,el1_way,el0_way;
  wire v_o,empty_o,full_o,bypass_track_o,N0,el0_valid,el1_valid,tag_hit0_n,tag_hit1_n,
  tag_hit2_n,tag_hit0,tag_hit1,tag_hit2,bypass_track_n,N1,N2,N3;
  reg bypass_track_o_sv2v_reg;
  assign bypass_track_o = bypass_track_o_sv2v_reg;

  bsg_cache_buffer_queue_00000024
  q0
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .data_i({ addr_i, way_i }),
    .v_o(v_o),
    .data_o({ addr_o, way_o }),
    .yumi_i(yumi_i),
    .el0_valid_o(el0_valid),
    .el1_valid_o(el1_valid),
    .el0_snoop_o({ el0_addr, el0_way }),
    .el1_snoop_o({ el1_addr, el1_way }),
    .empty_o(empty_o),
    .full_o(full_o)
  );

  assign tag_hit0_n = bypass_addr_i[32:4] == el0_addr[32:4];
  assign tag_hit1_n = bypass_addr_i[32:4] == el1_addr[32:4];
  assign tag_hit2_n = bypass_addr_i[32:4] == addr_i[32:4];
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = bypass_v_i;
  assign tag_hit0 = tag_hit0_n & el0_valid;
  assign tag_hit1 = tag_hit1_n & el1_valid;
  assign tag_hit2 = tag_hit2_n & v_i;
  assign bypass_track_n = N3 | tag_hit2;
  assign N3 = tag_hit0 | tag_hit1;
  assign N1 = ~bypass_v_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      bypass_track_o_sv2v_reg <= 1'b0;
    end else if(N2) begin
      bypass_track_o_sv2v_reg <= bypass_track_n;
    end 
  end


endmodule



module bsg_expand_bitmask_00000010_8
(
  i,
  o
);

  input [15:0] i;
  output [127:0] o;
  wire [127:0] o;
  wire o_127_,o_119_,o_111_,o_103_,o_95_,o_87_,o_79_,o_71_,o_63_,o_55_,o_47_,o_39_,
  o_31_,o_23_,o_15_,o_7_;
  assign o_127_ = i[15];
  assign o[120] = o_127_;
  assign o[121] = o_127_;
  assign o[122] = o_127_;
  assign o[123] = o_127_;
  assign o[124] = o_127_;
  assign o[125] = o_127_;
  assign o[126] = o_127_;
  assign o[127] = o_127_;
  assign o_119_ = i[14];
  assign o[112] = o_119_;
  assign o[113] = o_119_;
  assign o[114] = o_119_;
  assign o[115] = o_119_;
  assign o[116] = o_119_;
  assign o[117] = o_119_;
  assign o[118] = o_119_;
  assign o[119] = o_119_;
  assign o_111_ = i[13];
  assign o[104] = o_111_;
  assign o[105] = o_111_;
  assign o[106] = o_111_;
  assign o[107] = o_111_;
  assign o[108] = o_111_;
  assign o[109] = o_111_;
  assign o[110] = o_111_;
  assign o[111] = o_111_;
  assign o_103_ = i[12];
  assign o[96] = o_103_;
  assign o[97] = o_103_;
  assign o[98] = o_103_;
  assign o[99] = o_103_;
  assign o[100] = o_103_;
  assign o[101] = o_103_;
  assign o[102] = o_103_;
  assign o[103] = o_103_;
  assign o_95_ = i[11];
  assign o[88] = o_95_;
  assign o[89] = o_95_;
  assign o[90] = o_95_;
  assign o[91] = o_95_;
  assign o[92] = o_95_;
  assign o[93] = o_95_;
  assign o[94] = o_95_;
  assign o[95] = o_95_;
  assign o_87_ = i[10];
  assign o[80] = o_87_;
  assign o[81] = o_87_;
  assign o[82] = o_87_;
  assign o[83] = o_87_;
  assign o[84] = o_87_;
  assign o[85] = o_87_;
  assign o[86] = o_87_;
  assign o[87] = o_87_;
  assign o_79_ = i[9];
  assign o[72] = o_79_;
  assign o[73] = o_79_;
  assign o[74] = o_79_;
  assign o[75] = o_79_;
  assign o[76] = o_79_;
  assign o[77] = o_79_;
  assign o[78] = o_79_;
  assign o[79] = o_79_;
  assign o_71_ = i[8];
  assign o[64] = o_71_;
  assign o[65] = o_71_;
  assign o[66] = o_71_;
  assign o[67] = o_71_;
  assign o[68] = o_71_;
  assign o[69] = o_71_;
  assign o[70] = o_71_;
  assign o[71] = o_71_;
  assign o_63_ = i[7];
  assign o[56] = o_63_;
  assign o[57] = o_63_;
  assign o[58] = o_63_;
  assign o[59] = o_63_;
  assign o[60] = o_63_;
  assign o[61] = o_63_;
  assign o[62] = o_63_;
  assign o[63] = o_63_;
  assign o_55_ = i[6];
  assign o[48] = o_55_;
  assign o[49] = o_55_;
  assign o[50] = o_55_;
  assign o[51] = o_55_;
  assign o[52] = o_55_;
  assign o[53] = o_55_;
  assign o[54] = o_55_;
  assign o[55] = o_55_;
  assign o_47_ = i[5];
  assign o[40] = o_47_;
  assign o[41] = o_47_;
  assign o[42] = o_47_;
  assign o[43] = o_47_;
  assign o[44] = o_47_;
  assign o[45] = o_47_;
  assign o[46] = o_47_;
  assign o[47] = o_47_;
  assign o_39_ = i[4];
  assign o[32] = o_39_;
  assign o[33] = o_39_;
  assign o[34] = o_39_;
  assign o[35] = o_39_;
  assign o[36] = o_39_;
  assign o[37] = o_39_;
  assign o[38] = o_39_;
  assign o[39] = o_39_;
  assign o_31_ = i[3];
  assign o[24] = o_31_;
  assign o[25] = o_31_;
  assign o[26] = o_31_;
  assign o[27] = o_31_;
  assign o[28] = o_31_;
  assign o[29] = o_31_;
  assign o[30] = o_31_;
  assign o[31] = o_31_;
  assign o_23_ = i[2];
  assign o[16] = o_23_;
  assign o[17] = o_23_;
  assign o[18] = o_23_;
  assign o[19] = o_23_;
  assign o[20] = o_23_;
  assign o[21] = o_23_;
  assign o[22] = o_23_;
  assign o[23] = o_23_;
  assign o_15_ = i[1];
  assign o[8] = o_15_;
  assign o[9] = o_15_;
  assign o[10] = o_15_;
  assign o[11] = o_15_;
  assign o[12] = o_15_;
  assign o[13] = o_15_;
  assign o[14] = o_15_;
  assign o[15] = o_15_;
  assign o_7_ = i[0];
  assign o[0] = o_7_;
  assign o[1] = o_7_;
  assign o[2] = o_7_;
  assign o[3] = o_7_;
  assign o[4] = o_7_;
  assign o[5] = o_7_;
  assign o[6] = o_7_;
  assign o[7] = o_7_;

endmodule



module bsg_mux_8_00000010
(
  data_i,
  sel_i,
  data_o
);

  input [127:0] data_i;
  input [3:0] sel_i;
  output [7:0] data_o;
  wire [7:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31;
  assign data_o[7] = (N16)? data_i[7] : 
                     (N18)? data_i[15] : 
                     (N20)? data_i[23] : 
                     (N22)? data_i[31] : 
                     (N24)? data_i[39] : 
                     (N26)? data_i[47] : 
                     (N28)? data_i[55] : 
                     (N30)? data_i[63] : 
                     (N17)? data_i[71] : 
                     (N19)? data_i[79] : 
                     (N21)? data_i[87] : 
                     (N23)? data_i[95] : 
                     (N25)? data_i[103] : 
                     (N27)? data_i[111] : 
                     (N29)? data_i[119] : 
                     (N31)? data_i[127] : 1'b0;
  assign data_o[6] = (N16)? data_i[6] : 
                     (N18)? data_i[14] : 
                     (N20)? data_i[22] : 
                     (N22)? data_i[30] : 
                     (N24)? data_i[38] : 
                     (N26)? data_i[46] : 
                     (N28)? data_i[54] : 
                     (N30)? data_i[62] : 
                     (N17)? data_i[70] : 
                     (N19)? data_i[78] : 
                     (N21)? data_i[86] : 
                     (N23)? data_i[94] : 
                     (N25)? data_i[102] : 
                     (N27)? data_i[110] : 
                     (N29)? data_i[118] : 
                     (N31)? data_i[126] : 1'b0;
  assign data_o[5] = (N16)? data_i[5] : 
                     (N18)? data_i[13] : 
                     (N20)? data_i[21] : 
                     (N22)? data_i[29] : 
                     (N24)? data_i[37] : 
                     (N26)? data_i[45] : 
                     (N28)? data_i[53] : 
                     (N30)? data_i[61] : 
                     (N17)? data_i[69] : 
                     (N19)? data_i[77] : 
                     (N21)? data_i[85] : 
                     (N23)? data_i[93] : 
                     (N25)? data_i[101] : 
                     (N27)? data_i[109] : 
                     (N29)? data_i[117] : 
                     (N31)? data_i[125] : 1'b0;
  assign data_o[4] = (N16)? data_i[4] : 
                     (N18)? data_i[12] : 
                     (N20)? data_i[20] : 
                     (N22)? data_i[28] : 
                     (N24)? data_i[36] : 
                     (N26)? data_i[44] : 
                     (N28)? data_i[52] : 
                     (N30)? data_i[60] : 
                     (N17)? data_i[68] : 
                     (N19)? data_i[76] : 
                     (N21)? data_i[84] : 
                     (N23)? data_i[92] : 
                     (N25)? data_i[100] : 
                     (N27)? data_i[108] : 
                     (N29)? data_i[116] : 
                     (N31)? data_i[124] : 1'b0;
  assign data_o[3] = (N16)? data_i[3] : 
                     (N18)? data_i[11] : 
                     (N20)? data_i[19] : 
                     (N22)? data_i[27] : 
                     (N24)? data_i[35] : 
                     (N26)? data_i[43] : 
                     (N28)? data_i[51] : 
                     (N30)? data_i[59] : 
                     (N17)? data_i[67] : 
                     (N19)? data_i[75] : 
                     (N21)? data_i[83] : 
                     (N23)? data_i[91] : 
                     (N25)? data_i[99] : 
                     (N27)? data_i[107] : 
                     (N29)? data_i[115] : 
                     (N31)? data_i[123] : 1'b0;
  assign data_o[2] = (N16)? data_i[2] : 
                     (N18)? data_i[10] : 
                     (N20)? data_i[18] : 
                     (N22)? data_i[26] : 
                     (N24)? data_i[34] : 
                     (N26)? data_i[42] : 
                     (N28)? data_i[50] : 
                     (N30)? data_i[58] : 
                     (N17)? data_i[66] : 
                     (N19)? data_i[74] : 
                     (N21)? data_i[82] : 
                     (N23)? data_i[90] : 
                     (N25)? data_i[98] : 
                     (N27)? data_i[106] : 
                     (N29)? data_i[114] : 
                     (N31)? data_i[122] : 1'b0;
  assign data_o[1] = (N16)? data_i[1] : 
                     (N18)? data_i[9] : 
                     (N20)? data_i[17] : 
                     (N22)? data_i[25] : 
                     (N24)? data_i[33] : 
                     (N26)? data_i[41] : 
                     (N28)? data_i[49] : 
                     (N30)? data_i[57] : 
                     (N17)? data_i[65] : 
                     (N19)? data_i[73] : 
                     (N21)? data_i[81] : 
                     (N23)? data_i[89] : 
                     (N25)? data_i[97] : 
                     (N27)? data_i[105] : 
                     (N29)? data_i[113] : 
                     (N31)? data_i[121] : 1'b0;
  assign data_o[0] = (N16)? data_i[0] : 
                     (N18)? data_i[8] : 
                     (N20)? data_i[16] : 
                     (N22)? data_i[24] : 
                     (N24)? data_i[32] : 
                     (N26)? data_i[40] : 
                     (N28)? data_i[48] : 
                     (N30)? data_i[56] : 
                     (N17)? data_i[64] : 
                     (N19)? data_i[72] : 
                     (N21)? data_i[80] : 
                     (N23)? data_i[88] : 
                     (N25)? data_i[96] : 
                     (N27)? data_i[104] : 
                     (N29)? data_i[112] : 
                     (N31)? data_i[120] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];
  assign N6 = ~sel_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & sel_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & sel_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & sel_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & sel_i[2];
  assign N15 = ~sel_i[3];
  assign N16 = N7 & N15;
  assign N17 = N7 & sel_i[3];
  assign N18 = N9 & N15;
  assign N19 = N9 & sel_i[3];
  assign N20 = N11 & N15;
  assign N21 = N11 & sel_i[3];
  assign N22 = N13 & N15;
  assign N23 = N13 & sel_i[3];
  assign N24 = N8 & N15;
  assign N25 = N8 & sel_i[3];
  assign N26 = N10 & N15;
  assign N27 = N10 & sel_i[3];
  assign N28 = N12 & N15;
  assign N29 = N12 & sel_i[3];
  assign N30 = N14 & N15;
  assign N31 = N14 & sel_i[3];

endmodule



module bsg_mux_16_00000008
(
  data_i,
  sel_i,
  data_o
);

  input [127:0] data_i;
  input [2:0] sel_i;
  output [15:0] data_o;
  wire [15:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;
  assign data_o[15] = (N7)? data_i[15] : 
                      (N9)? data_i[31] : 
                      (N11)? data_i[47] : 
                      (N13)? data_i[63] : 
                      (N8)? data_i[79] : 
                      (N10)? data_i[95] : 
                      (N12)? data_i[111] : 
                      (N14)? data_i[127] : 1'b0;
  assign data_o[14] = (N7)? data_i[14] : 
                      (N9)? data_i[30] : 
                      (N11)? data_i[46] : 
                      (N13)? data_i[62] : 
                      (N8)? data_i[78] : 
                      (N10)? data_i[94] : 
                      (N12)? data_i[110] : 
                      (N14)? data_i[126] : 1'b0;
  assign data_o[13] = (N7)? data_i[13] : 
                      (N9)? data_i[29] : 
                      (N11)? data_i[45] : 
                      (N13)? data_i[61] : 
                      (N8)? data_i[77] : 
                      (N10)? data_i[93] : 
                      (N12)? data_i[109] : 
                      (N14)? data_i[125] : 1'b0;
  assign data_o[12] = (N7)? data_i[12] : 
                      (N9)? data_i[28] : 
                      (N11)? data_i[44] : 
                      (N13)? data_i[60] : 
                      (N8)? data_i[76] : 
                      (N10)? data_i[92] : 
                      (N12)? data_i[108] : 
                      (N14)? data_i[124] : 1'b0;
  assign data_o[11] = (N7)? data_i[11] : 
                      (N9)? data_i[27] : 
                      (N11)? data_i[43] : 
                      (N13)? data_i[59] : 
                      (N8)? data_i[75] : 
                      (N10)? data_i[91] : 
                      (N12)? data_i[107] : 
                      (N14)? data_i[123] : 1'b0;
  assign data_o[10] = (N7)? data_i[10] : 
                      (N9)? data_i[26] : 
                      (N11)? data_i[42] : 
                      (N13)? data_i[58] : 
                      (N8)? data_i[74] : 
                      (N10)? data_i[90] : 
                      (N12)? data_i[106] : 
                      (N14)? data_i[122] : 1'b0;
  assign data_o[9] = (N7)? data_i[9] : 
                     (N9)? data_i[25] : 
                     (N11)? data_i[41] : 
                     (N13)? data_i[57] : 
                     (N8)? data_i[73] : 
                     (N10)? data_i[89] : 
                     (N12)? data_i[105] : 
                     (N14)? data_i[121] : 1'b0;
  assign data_o[8] = (N7)? data_i[8] : 
                     (N9)? data_i[24] : 
                     (N11)? data_i[40] : 
                     (N13)? data_i[56] : 
                     (N8)? data_i[72] : 
                     (N10)? data_i[88] : 
                     (N12)? data_i[104] : 
                     (N14)? data_i[120] : 1'b0;
  assign data_o[7] = (N7)? data_i[7] : 
                     (N9)? data_i[23] : 
                     (N11)? data_i[39] : 
                     (N13)? data_i[55] : 
                     (N8)? data_i[71] : 
                     (N10)? data_i[87] : 
                     (N12)? data_i[103] : 
                     (N14)? data_i[119] : 1'b0;
  assign data_o[6] = (N7)? data_i[6] : 
                     (N9)? data_i[22] : 
                     (N11)? data_i[38] : 
                     (N13)? data_i[54] : 
                     (N8)? data_i[70] : 
                     (N10)? data_i[86] : 
                     (N12)? data_i[102] : 
                     (N14)? data_i[118] : 1'b0;
  assign data_o[5] = (N7)? data_i[5] : 
                     (N9)? data_i[21] : 
                     (N11)? data_i[37] : 
                     (N13)? data_i[53] : 
                     (N8)? data_i[69] : 
                     (N10)? data_i[85] : 
                     (N12)? data_i[101] : 
                     (N14)? data_i[117] : 1'b0;
  assign data_o[4] = (N7)? data_i[4] : 
                     (N9)? data_i[20] : 
                     (N11)? data_i[36] : 
                     (N13)? data_i[52] : 
                     (N8)? data_i[68] : 
                     (N10)? data_i[84] : 
                     (N12)? data_i[100] : 
                     (N14)? data_i[116] : 1'b0;
  assign data_o[3] = (N7)? data_i[3] : 
                     (N9)? data_i[19] : 
                     (N11)? data_i[35] : 
                     (N13)? data_i[51] : 
                     (N8)? data_i[67] : 
                     (N10)? data_i[83] : 
                     (N12)? data_i[99] : 
                     (N14)? data_i[115] : 1'b0;
  assign data_o[2] = (N7)? data_i[2] : 
                     (N9)? data_i[18] : 
                     (N11)? data_i[34] : 
                     (N13)? data_i[50] : 
                     (N8)? data_i[66] : 
                     (N10)? data_i[82] : 
                     (N12)? data_i[98] : 
                     (N14)? data_i[114] : 1'b0;
  assign data_o[1] = (N7)? data_i[1] : 
                     (N9)? data_i[17] : 
                     (N11)? data_i[33] : 
                     (N13)? data_i[49] : 
                     (N8)? data_i[65] : 
                     (N10)? data_i[81] : 
                     (N12)? data_i[97] : 
                     (N14)? data_i[113] : 1'b0;
  assign data_o[0] = (N7)? data_i[0] : 
                     (N9)? data_i[16] : 
                     (N11)? data_i[32] : 
                     (N13)? data_i[48] : 
                     (N8)? data_i[64] : 
                     (N10)? data_i[80] : 
                     (N12)? data_i[96] : 
                     (N14)? data_i[112] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];
  assign N6 = ~sel_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & sel_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & sel_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & sel_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & sel_i[2];

endmodule



module bsg_mux_32_00000004
(
  data_i,
  sel_i,
  data_o
);

  input [127:0] data_i;
  input [1:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[31] = (N2)? data_i[31] : 
                      (N4)? data_i[63] : 
                      (N3)? data_i[95] : 
                      (N5)? data_i[127] : 1'b0;
  assign data_o[30] = (N2)? data_i[30] : 
                      (N4)? data_i[62] : 
                      (N3)? data_i[94] : 
                      (N5)? data_i[126] : 1'b0;
  assign data_o[29] = (N2)? data_i[29] : 
                      (N4)? data_i[61] : 
                      (N3)? data_i[93] : 
                      (N5)? data_i[125] : 1'b0;
  assign data_o[28] = (N2)? data_i[28] : 
                      (N4)? data_i[60] : 
                      (N3)? data_i[92] : 
                      (N5)? data_i[124] : 1'b0;
  assign data_o[27] = (N2)? data_i[27] : 
                      (N4)? data_i[59] : 
                      (N3)? data_i[91] : 
                      (N5)? data_i[123] : 1'b0;
  assign data_o[26] = (N2)? data_i[26] : 
                      (N4)? data_i[58] : 
                      (N3)? data_i[90] : 
                      (N5)? data_i[122] : 1'b0;
  assign data_o[25] = (N2)? data_i[25] : 
                      (N4)? data_i[57] : 
                      (N3)? data_i[89] : 
                      (N5)? data_i[121] : 1'b0;
  assign data_o[24] = (N2)? data_i[24] : 
                      (N4)? data_i[56] : 
                      (N3)? data_i[88] : 
                      (N5)? data_i[120] : 1'b0;
  assign data_o[23] = (N2)? data_i[23] : 
                      (N4)? data_i[55] : 
                      (N3)? data_i[87] : 
                      (N5)? data_i[119] : 1'b0;
  assign data_o[22] = (N2)? data_i[22] : 
                      (N4)? data_i[54] : 
                      (N3)? data_i[86] : 
                      (N5)? data_i[118] : 1'b0;
  assign data_o[21] = (N2)? data_i[21] : 
                      (N4)? data_i[53] : 
                      (N3)? data_i[85] : 
                      (N5)? data_i[117] : 1'b0;
  assign data_o[20] = (N2)? data_i[20] : 
                      (N4)? data_i[52] : 
                      (N3)? data_i[84] : 
                      (N5)? data_i[116] : 1'b0;
  assign data_o[19] = (N2)? data_i[19] : 
                      (N4)? data_i[51] : 
                      (N3)? data_i[83] : 
                      (N5)? data_i[115] : 1'b0;
  assign data_o[18] = (N2)? data_i[18] : 
                      (N4)? data_i[50] : 
                      (N3)? data_i[82] : 
                      (N5)? data_i[114] : 1'b0;
  assign data_o[17] = (N2)? data_i[17] : 
                      (N4)? data_i[49] : 
                      (N3)? data_i[81] : 
                      (N5)? data_i[113] : 1'b0;
  assign data_o[16] = (N2)? data_i[16] : 
                      (N4)? data_i[48] : 
                      (N3)? data_i[80] : 
                      (N5)? data_i[112] : 1'b0;
  assign data_o[15] = (N2)? data_i[15] : 
                      (N4)? data_i[47] : 
                      (N3)? data_i[79] : 
                      (N5)? data_i[111] : 1'b0;
  assign data_o[14] = (N2)? data_i[14] : 
                      (N4)? data_i[46] : 
                      (N3)? data_i[78] : 
                      (N5)? data_i[110] : 1'b0;
  assign data_o[13] = (N2)? data_i[13] : 
                      (N4)? data_i[45] : 
                      (N3)? data_i[77] : 
                      (N5)? data_i[109] : 1'b0;
  assign data_o[12] = (N2)? data_i[12] : 
                      (N4)? data_i[44] : 
                      (N3)? data_i[76] : 
                      (N5)? data_i[108] : 1'b0;
  assign data_o[11] = (N2)? data_i[11] : 
                      (N4)? data_i[43] : 
                      (N3)? data_i[75] : 
                      (N5)? data_i[107] : 1'b0;
  assign data_o[10] = (N2)? data_i[10] : 
                      (N4)? data_i[42] : 
                      (N3)? data_i[74] : 
                      (N5)? data_i[106] : 1'b0;
  assign data_o[9] = (N2)? data_i[9] : 
                     (N4)? data_i[41] : 
                     (N3)? data_i[73] : 
                     (N5)? data_i[105] : 1'b0;
  assign data_o[8] = (N2)? data_i[8] : 
                     (N4)? data_i[40] : 
                     (N3)? data_i[72] : 
                     (N5)? data_i[104] : 1'b0;
  assign data_o[7] = (N2)? data_i[7] : 
                     (N4)? data_i[39] : 
                     (N3)? data_i[71] : 
                     (N5)? data_i[103] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] : 
                     (N4)? data_i[38] : 
                     (N3)? data_i[70] : 
                     (N5)? data_i[102] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] : 
                     (N4)? data_i[37] : 
                     (N3)? data_i[69] : 
                     (N5)? data_i[101] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] : 
                     (N4)? data_i[36] : 
                     (N3)? data_i[68] : 
                     (N5)? data_i[100] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] : 
                     (N4)? data_i[35] : 
                     (N3)? data_i[67] : 
                     (N5)? data_i[99] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] : 
                     (N4)? data_i[34] : 
                     (N3)? data_i[66] : 
                     (N5)? data_i[98] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N4)? data_i[33] : 
                     (N3)? data_i[65] : 
                     (N5)? data_i[97] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[32] : 
                     (N3)? data_i[64] : 
                     (N5)? data_i[96] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_mux_64_00000002
(
  data_i,
  sel_i,
  data_o
);

  input [127:0] data_i;
  input [0:0] sel_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1;
  assign data_o[63] = (N1)? data_i[63] : 
                      (N0)? data_i[127] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[62] = (N1)? data_i[62] : 
                      (N0)? data_i[126] : 1'b0;
  assign data_o[61] = (N1)? data_i[61] : 
                      (N0)? data_i[125] : 1'b0;
  assign data_o[60] = (N1)? data_i[60] : 
                      (N0)? data_i[124] : 1'b0;
  assign data_o[59] = (N1)? data_i[59] : 
                      (N0)? data_i[123] : 1'b0;
  assign data_o[58] = (N1)? data_i[58] : 
                      (N0)? data_i[122] : 1'b0;
  assign data_o[57] = (N1)? data_i[57] : 
                      (N0)? data_i[121] : 1'b0;
  assign data_o[56] = (N1)? data_i[56] : 
                      (N0)? data_i[120] : 1'b0;
  assign data_o[55] = (N1)? data_i[55] : 
                      (N0)? data_i[119] : 1'b0;
  assign data_o[54] = (N1)? data_i[54] : 
                      (N0)? data_i[118] : 1'b0;
  assign data_o[53] = (N1)? data_i[53] : 
                      (N0)? data_i[117] : 1'b0;
  assign data_o[52] = (N1)? data_i[52] : 
                      (N0)? data_i[116] : 1'b0;
  assign data_o[51] = (N1)? data_i[51] : 
                      (N0)? data_i[115] : 1'b0;
  assign data_o[50] = (N1)? data_i[50] : 
                      (N0)? data_i[114] : 1'b0;
  assign data_o[49] = (N1)? data_i[49] : 
                      (N0)? data_i[113] : 1'b0;
  assign data_o[48] = (N1)? data_i[48] : 
                      (N0)? data_i[112] : 1'b0;
  assign data_o[47] = (N1)? data_i[47] : 
                      (N0)? data_i[111] : 1'b0;
  assign data_o[46] = (N1)? data_i[46] : 
                      (N0)? data_i[110] : 1'b0;
  assign data_o[45] = (N1)? data_i[45] : 
                      (N0)? data_i[109] : 1'b0;
  assign data_o[44] = (N1)? data_i[44] : 
                      (N0)? data_i[108] : 1'b0;
  assign data_o[43] = (N1)? data_i[43] : 
                      (N0)? data_i[107] : 1'b0;
  assign data_o[42] = (N1)? data_i[42] : 
                      (N0)? data_i[106] : 1'b0;
  assign data_o[41] = (N1)? data_i[41] : 
                      (N0)? data_i[105] : 1'b0;
  assign data_o[40] = (N1)? data_i[40] : 
                      (N0)? data_i[104] : 1'b0;
  assign data_o[39] = (N1)? data_i[39] : 
                      (N0)? data_i[103] : 1'b0;
  assign data_o[38] = (N1)? data_i[38] : 
                      (N0)? data_i[102] : 1'b0;
  assign data_o[37] = (N1)? data_i[37] : 
                      (N0)? data_i[101] : 1'b0;
  assign data_o[36] = (N1)? data_i[36] : 
                      (N0)? data_i[100] : 1'b0;
  assign data_o[35] = (N1)? data_i[35] : 
                      (N0)? data_i[99] : 1'b0;
  assign data_o[34] = (N1)? data_i[34] : 
                      (N0)? data_i[98] : 1'b0;
  assign data_o[33] = (N1)? data_i[33] : 
                      (N0)? data_i[97] : 1'b0;
  assign data_o[32] = (N1)? data_i[32] : 
                      (N0)? data_i[96] : 1'b0;
  assign data_o[31] = (N1)? data_i[31] : 
                      (N0)? data_i[95] : 1'b0;
  assign data_o[30] = (N1)? data_i[30] : 
                      (N0)? data_i[94] : 1'b0;
  assign data_o[29] = (N1)? data_i[29] : 
                      (N0)? data_i[93] : 1'b0;
  assign data_o[28] = (N1)? data_i[28] : 
                      (N0)? data_i[92] : 1'b0;
  assign data_o[27] = (N1)? data_i[27] : 
                      (N0)? data_i[91] : 1'b0;
  assign data_o[26] = (N1)? data_i[26] : 
                      (N0)? data_i[90] : 1'b0;
  assign data_o[25] = (N1)? data_i[25] : 
                      (N0)? data_i[89] : 1'b0;
  assign data_o[24] = (N1)? data_i[24] : 
                      (N0)? data_i[88] : 1'b0;
  assign data_o[23] = (N1)? data_i[23] : 
                      (N0)? data_i[87] : 1'b0;
  assign data_o[22] = (N1)? data_i[22] : 
                      (N0)? data_i[86] : 1'b0;
  assign data_o[21] = (N1)? data_i[21] : 
                      (N0)? data_i[85] : 1'b0;
  assign data_o[20] = (N1)? data_i[20] : 
                      (N0)? data_i[84] : 1'b0;
  assign data_o[19] = (N1)? data_i[19] : 
                      (N0)? data_i[83] : 1'b0;
  assign data_o[18] = (N1)? data_i[18] : 
                      (N0)? data_i[82] : 1'b0;
  assign data_o[17] = (N1)? data_i[17] : 
                      (N0)? data_i[81] : 1'b0;
  assign data_o[16] = (N1)? data_i[16] : 
                      (N0)? data_i[80] : 1'b0;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[79] : 1'b0;
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[78] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[77] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[76] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[75] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[74] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[73] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[72] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[71] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[70] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[69] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[68] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[67] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[66] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[65] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[64] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_cache_00000021_00000080_00000004_00000080_00000008_1_1_00000080
(
  clk_i,
  reset_i,
  cache_pkt_i,
  v_i,
  yumi_o,
  data_o,
  v_o,
  yumi_i,
  dma_pkt_o,
  dma_pkt_v_o,
  dma_pkt_yumi_i,
  dma_data_i,
  dma_data_v_i,
  dma_data_ready_and_o,
  dma_data_o,
  dma_data_v_o,
  dma_data_yumi_i,
  v_we_o
);

  input [182:0] cache_pkt_i;
  output [127:0] data_o;
  output [37:0] dma_pkt_o;
  input [127:0] dma_data_i;
  output [127:0] dma_data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input dma_pkt_yumi_i;
  input dma_data_v_i;
  input dma_data_yumi_i;
  output yumi_o;
  output v_o;
  output dma_pkt_v_o;
  output dma_data_ready_and_o;
  output dma_data_v_o;
  output v_we_o;
  wire [127:0] data_o,dma_data_o,data_tl_r,data_mem_w_mask_li,data_v_r,snoop_word_lo,
  dma_data_mem_w_mask_lo,bypass_data_lo,sbuf_data_mem_w_mask,sbuf_data_in,
  ld_data_way_picked,ld_data_offset_picked,bypass_data_masked,snoop_or_ld_data,expanded_mask_v,
  ld_data_masked,ld_data_final_lo;
  wire [37:0] dma_pkt_o;
  wire yumi_o,v_o,dma_pkt_v_o,dma_data_ready_and_o,dma_data_v_o,v_we_o,N0,N1,N3,N4,N5,
  N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,
  N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,
  N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
  N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,tl_we,sbuf_hazard,N77,N78,v_tl_r,N79,N80,
  N81,N82,N83,N84,tag_mem_v_li,tag_mem_w_li,data_mem_v_li,data_mem_w_li,
  track_mem_v_li,track_mem_w_li,N85,N86,N87,v_v_r,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,
  N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,
  N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,tag_hit_found,N125,N126,N127,
  partial_st,N128,N129,N130,partial_st_tl,N131,N132,N133,N134,partial_st_v,
  ld_st_amo_tag_miss,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,bypass_track_lo,
  track_miss,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,
  N175,N176,tagfl_hit,aflinv_hit,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
  N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,alock_miss,N197,N198,N199,
  N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,
  aunlock_hit,miss_v,retval_op_v,stat_mem_v_li,stat_mem_w_li,sbuf_empty_lo,
  tbuf_empty_lo,dma_done_li,miss_track_data_we_lo,miss_stat_mem_v_lo,miss_stat_mem_w_lo,
  miss_tag_mem_v_lo,miss_tag_mem_w_lo,miss_track_mem_v_lo,miss_track_mem_w_lo,
  recover_lo,miss_done_lo,_1_net_,select_snoop_data_r_lo,dma_data_mem_v_lo,
  dma_data_mem_w_lo,dma_evict_lo,sbuf_entry_li_data__127_,sbuf_entry_li_data__126_,
  sbuf_entry_li_data__125_,sbuf_entry_li_data__124_,sbuf_entry_li_data__123_,
  sbuf_entry_li_data__122_,sbuf_entry_li_data__121_,sbuf_entry_li_data__120_,sbuf_entry_li_data__119_,
  sbuf_entry_li_data__118_,sbuf_entry_li_data__117_,sbuf_entry_li_data__116_,
  sbuf_entry_li_data__115_,sbuf_entry_li_data__114_,sbuf_entry_li_data__113_,
  sbuf_entry_li_data__112_,sbuf_entry_li_data__111_,sbuf_entry_li_data__110_,
  sbuf_entry_li_data__109_,sbuf_entry_li_data__108_,sbuf_entry_li_data__107_,
  sbuf_entry_li_data__106_,sbuf_entry_li_data__105_,sbuf_entry_li_data__104_,sbuf_entry_li_data__103_,
  sbuf_entry_li_data__102_,sbuf_entry_li_data__101_,sbuf_entry_li_data__100_,
  sbuf_entry_li_data__99_,sbuf_entry_li_data__98_,sbuf_entry_li_data__97_,
  sbuf_entry_li_data__96_,sbuf_entry_li_data__95_,sbuf_entry_li_data__94_,
  sbuf_entry_li_data__93_,sbuf_entry_li_data__92_,sbuf_entry_li_data__91_,sbuf_entry_li_data__90_,
  sbuf_entry_li_data__89_,sbuf_entry_li_data__88_,sbuf_entry_li_data__87_,
  sbuf_entry_li_data__86_,sbuf_entry_li_data__85_,sbuf_entry_li_data__84_,
  sbuf_entry_li_data__83_,sbuf_entry_li_data__82_,sbuf_entry_li_data__81_,sbuf_entry_li_data__80_,
  sbuf_entry_li_data__79_,sbuf_entry_li_data__78_,sbuf_entry_li_data__77_,
  sbuf_entry_li_data__76_,sbuf_entry_li_data__75_,sbuf_entry_li_data__74_,
  sbuf_entry_li_data__73_,sbuf_entry_li_data__72_,sbuf_entry_li_data__71_,sbuf_entry_li_data__70_,
  sbuf_entry_li_data__69_,sbuf_entry_li_data__68_,sbuf_entry_li_data__67_,
  sbuf_entry_li_data__66_,sbuf_entry_li_data__65_,sbuf_entry_li_data__64_,
  sbuf_entry_li_data__63_,sbuf_entry_li_data__62_,sbuf_entry_li_data__61_,sbuf_entry_li_data__60_,
  sbuf_entry_li_data__59_,sbuf_entry_li_data__58_,sbuf_entry_li_data__57_,
  sbuf_entry_li_data__56_,sbuf_entry_li_data__55_,sbuf_entry_li_data__54_,
  sbuf_entry_li_data__53_,sbuf_entry_li_data__52_,sbuf_entry_li_data__51_,sbuf_entry_li_data__50_,
  sbuf_entry_li_data__49_,sbuf_entry_li_data__48_,sbuf_entry_li_data__47_,
  sbuf_entry_li_data__46_,sbuf_entry_li_data__45_,sbuf_entry_li_data__44_,
  sbuf_entry_li_data__43_,sbuf_entry_li_data__42_,sbuf_entry_li_data__41_,sbuf_entry_li_data__40_,
  sbuf_entry_li_data__39_,sbuf_entry_li_data__38_,sbuf_entry_li_data__37_,
  sbuf_entry_li_data__36_,sbuf_entry_li_data__35_,sbuf_entry_li_data__34_,
  sbuf_entry_li_data__33_,sbuf_entry_li_data__32_,sbuf_entry_li_data__31_,sbuf_entry_li_data__30_,
  sbuf_entry_li_data__29_,sbuf_entry_li_data__28_,sbuf_entry_li_data__27_,
  sbuf_entry_li_data__26_,sbuf_entry_li_data__25_,sbuf_entry_li_data__24_,
  sbuf_entry_li_data__23_,sbuf_entry_li_data__22_,sbuf_entry_li_data__21_,sbuf_entry_li_data__20_,
  sbuf_entry_li_data__19_,sbuf_entry_li_data__18_,sbuf_entry_li_data__17_,
  sbuf_entry_li_data__16_,sbuf_entry_li_data__15_,sbuf_entry_li_data__14_,
  sbuf_entry_li_data__13_,sbuf_entry_li_data__12_,sbuf_entry_li_data__11_,sbuf_entry_li_data__10_,
  sbuf_entry_li_data__9_,sbuf_entry_li_data__8_,sbuf_entry_li_data__7_,
  sbuf_entry_li_data__6_,sbuf_entry_li_data__5_,sbuf_entry_li_data__4_,sbuf_entry_li_data__3_,
  sbuf_entry_li_data__2_,sbuf_entry_li_data__1_,sbuf_entry_li_data__0_,
  sbuf_entry_li_mask__15_,sbuf_entry_li_mask__14_,sbuf_entry_li_mask__13_,
  sbuf_entry_li_mask__12_,sbuf_entry_li_mask__11_,sbuf_entry_li_mask__10_,sbuf_entry_li_mask__9_,
  sbuf_entry_li_mask__8_,sbuf_entry_li_mask__7_,sbuf_entry_li_mask__6_,
  sbuf_entry_li_mask__5_,sbuf_entry_li_mask__4_,sbuf_entry_li_mask__3_,sbuf_entry_li_mask__2_,
  sbuf_entry_li_mask__1_,sbuf_entry_li_mask__0_,sbuf_entry_li_way_id__2_,
  sbuf_entry_li_way_id__1_,sbuf_entry_li_way_id__0_,sbuf_v_li,sbuf_v_lo,sbuf_yumi_li,sbuf_full_lo,
  sbuf_bypass_v_li,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
  ld_data_final_li_3__127_,ld_data_final_li_3__126_,ld_data_final_li_3__125_,
  ld_data_final_li_3__124_,ld_data_final_li_3__123_,ld_data_final_li_3__122_,
  ld_data_final_li_3__121_,ld_data_final_li_3__120_,ld_data_final_li_3__119_,ld_data_final_li_3__118_,
  ld_data_final_li_3__117_,ld_data_final_li_3__116_,ld_data_final_li_3__115_,
  ld_data_final_li_3__114_,ld_data_final_li_3__113_,ld_data_final_li_3__112_,
  ld_data_final_li_3__111_,ld_data_final_li_3__110_,ld_data_final_li_3__109_,
  ld_data_final_li_3__108_,ld_data_final_li_3__107_,ld_data_final_li_3__106_,
  ld_data_final_li_3__105_,ld_data_final_li_3__104_,ld_data_final_li_3__103_,ld_data_final_li_3__102_,
  ld_data_final_li_3__101_,ld_data_final_li_3__100_,ld_data_final_li_3__99_,
  ld_data_final_li_3__98_,ld_data_final_li_3__97_,ld_data_final_li_3__96_,
  ld_data_final_li_3__95_,ld_data_final_li_3__94_,ld_data_final_li_3__93_,ld_data_final_li_3__92_,
  ld_data_final_li_3__91_,ld_data_final_li_3__90_,ld_data_final_li_3__89_,
  ld_data_final_li_3__88_,ld_data_final_li_3__87_,ld_data_final_li_3__86_,
  ld_data_final_li_3__85_,ld_data_final_li_3__84_,ld_data_final_li_3__83_,ld_data_final_li_3__82_,
  ld_data_final_li_3__81_,ld_data_final_li_3__80_,ld_data_final_li_3__79_,
  ld_data_final_li_3__78_,ld_data_final_li_3__77_,ld_data_final_li_3__76_,
  ld_data_final_li_3__75_,ld_data_final_li_3__74_,ld_data_final_li_3__73_,ld_data_final_li_3__72_,
  ld_data_final_li_3__71_,ld_data_final_li_3__70_,ld_data_final_li_3__69_,
  ld_data_final_li_3__68_,ld_data_final_li_3__67_,ld_data_final_li_3__66_,
  ld_data_final_li_3__65_,ld_data_final_li_3__64_,ld_data_final_li_2__127_,
  ld_data_final_li_2__126_,ld_data_final_li_2__125_,ld_data_final_li_2__124_,ld_data_final_li_2__123_,
  ld_data_final_li_2__122_,ld_data_final_li_2__121_,ld_data_final_li_2__120_,
  ld_data_final_li_2__119_,ld_data_final_li_2__118_,ld_data_final_li_2__117_,
  ld_data_final_li_2__116_,ld_data_final_li_2__115_,ld_data_final_li_2__114_,
  ld_data_final_li_2__113_,ld_data_final_li_2__112_,ld_data_final_li_2__111_,
  ld_data_final_li_2__110_,ld_data_final_li_2__109_,ld_data_final_li_2__108_,ld_data_final_li_2__107_,
  ld_data_final_li_2__106_,ld_data_final_li_2__105_,ld_data_final_li_2__104_,
  ld_data_final_li_2__103_,ld_data_final_li_2__102_,ld_data_final_li_2__101_,
  ld_data_final_li_2__100_,ld_data_final_li_2__99_,ld_data_final_li_2__98_,
  ld_data_final_li_2__97_,ld_data_final_li_2__96_,ld_data_final_li_2__95_,ld_data_final_li_2__94_,
  ld_data_final_li_2__93_,ld_data_final_li_2__92_,ld_data_final_li_2__91_,
  ld_data_final_li_2__90_,ld_data_final_li_2__89_,ld_data_final_li_2__88_,
  ld_data_final_li_2__87_,ld_data_final_li_2__86_,ld_data_final_li_2__85_,ld_data_final_li_2__84_,
  ld_data_final_li_2__83_,ld_data_final_li_2__82_,ld_data_final_li_2__81_,
  ld_data_final_li_2__80_,ld_data_final_li_2__79_,ld_data_final_li_2__78_,
  ld_data_final_li_2__77_,ld_data_final_li_2__76_,ld_data_final_li_2__75_,ld_data_final_li_2__74_,
  ld_data_final_li_2__73_,ld_data_final_li_2__72_,ld_data_final_li_2__71_,
  ld_data_final_li_2__70_,ld_data_final_li_2__69_,ld_data_final_li_2__68_,
  ld_data_final_li_2__67_,ld_data_final_li_2__66_,ld_data_final_li_2__65_,ld_data_final_li_2__64_,
  ld_data_final_li_2__63_,ld_data_final_li_2__62_,ld_data_final_li_2__61_,
  ld_data_final_li_2__60_,ld_data_final_li_2__59_,ld_data_final_li_2__58_,
  ld_data_final_li_2__57_,ld_data_final_li_2__56_,ld_data_final_li_2__55_,ld_data_final_li_2__54_,
  ld_data_final_li_2__53_,ld_data_final_li_2__52_,ld_data_final_li_2__51_,
  ld_data_final_li_2__50_,ld_data_final_li_2__49_,ld_data_final_li_2__48_,
  ld_data_final_li_2__47_,ld_data_final_li_2__46_,ld_data_final_li_2__45_,ld_data_final_li_2__44_,
  ld_data_final_li_2__43_,ld_data_final_li_2__42_,ld_data_final_li_2__41_,
  ld_data_final_li_2__40_,ld_data_final_li_2__39_,ld_data_final_li_2__38_,
  ld_data_final_li_2__37_,ld_data_final_li_2__36_,ld_data_final_li_2__35_,ld_data_final_li_2__34_,
  ld_data_final_li_2__33_,ld_data_final_li_2__32_,ld_data_final_li_1__127_,
  ld_data_final_li_1__126_,ld_data_final_li_1__125_,ld_data_final_li_1__124_,
  ld_data_final_li_1__123_,ld_data_final_li_1__122_,ld_data_final_li_1__121_,
  ld_data_final_li_1__120_,ld_data_final_li_1__119_,ld_data_final_li_1__118_,ld_data_final_li_1__117_,
  ld_data_final_li_1__116_,ld_data_final_li_1__115_,ld_data_final_li_1__114_,
  ld_data_final_li_1__113_,ld_data_final_li_1__112_,ld_data_final_li_1__111_,
  ld_data_final_li_1__110_,ld_data_final_li_1__109_,ld_data_final_li_1__108_,
  ld_data_final_li_1__107_,ld_data_final_li_1__106_,ld_data_final_li_1__105_,
  ld_data_final_li_1__104_,ld_data_final_li_1__103_,ld_data_final_li_1__102_,ld_data_final_li_1__101_,
  ld_data_final_li_1__100_,ld_data_final_li_1__99_,ld_data_final_li_1__98_,
  ld_data_final_li_1__97_,ld_data_final_li_1__96_,ld_data_final_li_1__95_,
  ld_data_final_li_1__94_,ld_data_final_li_1__93_,ld_data_final_li_1__92_,ld_data_final_li_1__91_,
  ld_data_final_li_1__90_,ld_data_final_li_1__89_,ld_data_final_li_1__88_,
  ld_data_final_li_1__87_,ld_data_final_li_1__86_,ld_data_final_li_1__85_,
  ld_data_final_li_1__84_,ld_data_final_li_1__83_,ld_data_final_li_1__82_,ld_data_final_li_1__81_,
  ld_data_final_li_1__80_,ld_data_final_li_1__79_,ld_data_final_li_1__78_,
  ld_data_final_li_1__77_,ld_data_final_li_1__76_,ld_data_final_li_1__75_,
  ld_data_final_li_1__74_,ld_data_final_li_1__73_,ld_data_final_li_1__72_,ld_data_final_li_1__71_,
  ld_data_final_li_1__70_,ld_data_final_li_1__69_,ld_data_final_li_1__68_,
  ld_data_final_li_1__67_,ld_data_final_li_1__66_,ld_data_final_li_1__65_,
  ld_data_final_li_1__64_,ld_data_final_li_1__63_,ld_data_final_li_1__62_,ld_data_final_li_1__61_,
  ld_data_final_li_1__60_,ld_data_final_li_1__59_,ld_data_final_li_1__58_,
  ld_data_final_li_1__57_,ld_data_final_li_1__56_,ld_data_final_li_1__55_,
  ld_data_final_li_1__54_,ld_data_final_li_1__53_,ld_data_final_li_1__52_,ld_data_final_li_1__51_,
  ld_data_final_li_1__50_,ld_data_final_li_1__49_,ld_data_final_li_1__48_,
  ld_data_final_li_1__47_,ld_data_final_li_1__46_,ld_data_final_li_1__45_,
  ld_data_final_li_1__44_,ld_data_final_li_1__43_,ld_data_final_li_1__42_,ld_data_final_li_1__41_,
  ld_data_final_li_1__40_,ld_data_final_li_1__39_,ld_data_final_li_1__38_,
  ld_data_final_li_1__37_,ld_data_final_li_1__36_,ld_data_final_li_1__35_,
  ld_data_final_li_1__34_,ld_data_final_li_1__33_,ld_data_final_li_1__32_,ld_data_final_li_1__31_,
  ld_data_final_li_1__30_,ld_data_final_li_1__29_,ld_data_final_li_1__28_,
  ld_data_final_li_1__27_,ld_data_final_li_1__26_,ld_data_final_li_1__25_,
  ld_data_final_li_1__24_,ld_data_final_li_1__23_,ld_data_final_li_1__22_,ld_data_final_li_1__21_,
  ld_data_final_li_1__20_,ld_data_final_li_1__19_,ld_data_final_li_1__18_,
  ld_data_final_li_1__17_,ld_data_final_li_1__16_,ld_data_final_li_0__127_,
  ld_data_final_li_0__126_,ld_data_final_li_0__125_,ld_data_final_li_0__124_,
  ld_data_final_li_0__123_,ld_data_final_li_0__122_,ld_data_final_li_0__121_,ld_data_final_li_0__120_,
  ld_data_final_li_0__119_,ld_data_final_li_0__118_,ld_data_final_li_0__117_,
  ld_data_final_li_0__116_,ld_data_final_li_0__115_,ld_data_final_li_0__114_,
  ld_data_final_li_0__113_,ld_data_final_li_0__112_,ld_data_final_li_0__111_,
  ld_data_final_li_0__110_,ld_data_final_li_0__109_,ld_data_final_li_0__108_,
  ld_data_final_li_0__107_,ld_data_final_li_0__106_,ld_data_final_li_0__105_,ld_data_final_li_0__104_,
  ld_data_final_li_0__103_,ld_data_final_li_0__102_,ld_data_final_li_0__101_,
  ld_data_final_li_0__100_,ld_data_final_li_0__99_,ld_data_final_li_0__98_,
  ld_data_final_li_0__97_,ld_data_final_li_0__96_,ld_data_final_li_0__95_,
  ld_data_final_li_0__94_,ld_data_final_li_0__93_,ld_data_final_li_0__92_,ld_data_final_li_0__91_,
  ld_data_final_li_0__90_,ld_data_final_li_0__89_,ld_data_final_li_0__88_,
  ld_data_final_li_0__87_,ld_data_final_li_0__86_,ld_data_final_li_0__85_,
  ld_data_final_li_0__84_,ld_data_final_li_0__83_,ld_data_final_li_0__82_,ld_data_final_li_0__81_,
  ld_data_final_li_0__80_,ld_data_final_li_0__79_,ld_data_final_li_0__78_,
  ld_data_final_li_0__77_,ld_data_final_li_0__76_,ld_data_final_li_0__75_,
  ld_data_final_li_0__74_,ld_data_final_li_0__73_,ld_data_final_li_0__72_,ld_data_final_li_0__71_,
  ld_data_final_li_0__70_,ld_data_final_li_0__69_,ld_data_final_li_0__68_,
  ld_data_final_li_0__67_,ld_data_final_li_0__66_,ld_data_final_li_0__65_,
  ld_data_final_li_0__64_,ld_data_final_li_0__63_,ld_data_final_li_0__62_,ld_data_final_li_0__61_,
  ld_data_final_li_0__60_,ld_data_final_li_0__59_,ld_data_final_li_0__58_,
  ld_data_final_li_0__57_,ld_data_final_li_0__56_,ld_data_final_li_0__55_,
  ld_data_final_li_0__54_,ld_data_final_li_0__53_,ld_data_final_li_0__52_,ld_data_final_li_0__51_,
  ld_data_final_li_0__50_,ld_data_final_li_0__49_,ld_data_final_li_0__48_,
  ld_data_final_li_0__47_,ld_data_final_li_0__46_,ld_data_final_li_0__45_,
  ld_data_final_li_0__44_,ld_data_final_li_0__43_,ld_data_final_li_0__42_,ld_data_final_li_0__41_,
  ld_data_final_li_0__40_,ld_data_final_li_0__39_,ld_data_final_li_0__38_,
  ld_data_final_li_0__37_,ld_data_final_li_0__36_,ld_data_final_li_0__35_,
  ld_data_final_li_0__34_,ld_data_final_li_0__33_,ld_data_final_li_0__32_,ld_data_final_li_0__31_,
  ld_data_final_li_0__30_,ld_data_final_li_0__29_,ld_data_final_li_0__28_,
  ld_data_final_li_0__27_,ld_data_final_li_0__26_,ld_data_final_li_0__25_,
  ld_data_final_li_0__24_,ld_data_final_li_0__23_,ld_data_final_li_0__22_,ld_data_final_li_0__21_,
  ld_data_final_li_0__20_,ld_data_final_li_0__19_,ld_data_final_li_0__18_,
  ld_data_final_li_0__17_,ld_data_final_li_0__16_,ld_data_final_li_0__15_,
  ld_data_final_li_0__14_,ld_data_final_li_0__13_,ld_data_final_li_0__12_,ld_data_final_li_0__11_,
  ld_data_final_li_0__10_,ld_data_final_li_0__9_,ld_data_final_li_0__8_,N354,N355,N356,
  N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,
  N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,
  N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,
  N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,
  N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,
  N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,
  N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,
  N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,
  N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,
  N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,
  N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,
  N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,
  N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,
  N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,
  N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,
  N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,
  N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,
  N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,
  N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,
  N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,
  N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,
  N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,
  N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,
  N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,
  N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,
  N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,
  N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,
  N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,
  N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,
  N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,
  N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,
  N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,
  N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,
  N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,
  N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,
  N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,
  N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,
  N949,N950,tbuf_v_li,tbuf_v_lo,tbuf_yumi_li,tbuf_full_lo,tbuf_bypass_v_li,N951,
  N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,N966,N967,
  N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,N982,N983,
  N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,N998,N999,
  N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012,
  N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,
  N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038,N1039,
  N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,
  N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,
  N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079,
  N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091,N1092,
  N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,
  N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118,N1119,
  N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,N1131,N1132,
  N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,
  N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
  N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,N1171,N1172,
  N1173,N1174,N1175,tl_ready,N1176,N1177,tagst_write_en,N1178,N1179,N1180,N1181,N1182,
  N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,
  N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,
  N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,
  N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,
  N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,
  N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,
  N1263,N1264,N1265,N1266,N1267,N2,N1268,N1269,N1270,N1271,N1272,N1273,N1274,
  N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,
  N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,
  N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,
  N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,
  N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,
  N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,
  N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,
  N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,
  N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,
  N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,
  N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,
  N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,
  N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,
  N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461;
  wire [20:0] decode,decode_tl_r,decode_v_r;
  wire [15:0] mask_tl_r,mask_v_r,bypass_mask_lo,sbuf_expand_mask,sbuf_mask_in,
  \sbuf_in_sel_0_.decode_lo ,\ld_data_sel_1_.byte_sel ;
  wire [32:0] addr_tl_r,addr_v_r,dma_addr_lo,tbuf_addr_lo;
  wire [6:0] tag_mem_addr_li,track_mem_addr_li,stat_mem_addr_li,miss_stat_mem_addr_lo,
  miss_tag_mem_addr_lo,miss_track_mem_addr_lo,plru_decode_data_lo,plru_decode_mask_lo;
  wire [175:0] tag_mem_data_li,tag_mem_w_mask_li,tag_mem_data_lo,miss_tag_mem_data_lo,
  miss_tag_mem_w_mask_lo;
  wire [8:0] data_mem_addr_li,dma_data_mem_addr_lo;
  wire [1023:0] data_mem_data_li,data_mem_data_lo,ld_data_v_r,dma_data_mem_data_lo;
  wire [31:0] track_mem_data_li,track_mem_w_mask_li,track_mem_data_lo,track_data_v_r,
  miss_track_mem_w_mask_lo,miss_track_mem_data_lo,\sbuf_in_sel_2_.slice_data ,
  tbuf_track_mem_w_mask;
  wire [7:0] valid_v_r,lock_v_r,tag_hit_v,sbuf_way_decode,\sbuf_in_sel_1_.decode_lo ,
  tbuf_way_decode,\ld_data_sel_0_.byte_sel ,addr_way_decode;
  wire [159:0] tag_v_r;
  wire [2:0] tag_hit_way_id,dma_way_lo,chosen_way_lo,tbuf_way_li,tbuf_way_lo;
  wire [14:0] stat_mem_data_li,stat_mem_w_mask_li,stat_mem_data_lo,miss_stat_mem_data_lo,
  miss_stat_mem_w_mask_lo;
  wire [3:0] dma_cmd_lo,\sbuf_in_sel_2_.decode_lo ,tbuf_word_offset_decode;
  wire [179:0] sbuf_entry_lo;
  wire [0:0] sbuf_burst_offset_decode;
  wire [63:0] sbuf_mask_in_mux_li,atomic_reg_data,\atomic_64.amo64_mem_in ,atomic_mem_data,
  atomic_alu_result,atomic_result,\sbuf_in_sel_3_.slice_data ;
  wire [63:32] \atomic_64.amo32_mem_in ;
  wire [1:0] \sbuf_in_sel_3_.decode_lo ;
  reg data_tl_r_127_sv2v_reg,data_tl_r_126_sv2v_reg,data_tl_r_125_sv2v_reg,
  data_tl_r_124_sv2v_reg,data_tl_r_123_sv2v_reg,data_tl_r_122_sv2v_reg,
  data_tl_r_121_sv2v_reg,data_tl_r_120_sv2v_reg,data_tl_r_119_sv2v_reg,data_tl_r_118_sv2v_reg,
  data_tl_r_117_sv2v_reg,data_tl_r_116_sv2v_reg,data_tl_r_115_sv2v_reg,
  data_tl_r_114_sv2v_reg,data_tl_r_113_sv2v_reg,data_tl_r_112_sv2v_reg,data_tl_r_111_sv2v_reg,
  data_tl_r_110_sv2v_reg,data_tl_r_109_sv2v_reg,data_tl_r_108_sv2v_reg,
  data_tl_r_107_sv2v_reg,data_tl_r_106_sv2v_reg,data_tl_r_105_sv2v_reg,data_tl_r_104_sv2v_reg,
  data_tl_r_103_sv2v_reg,data_tl_r_102_sv2v_reg,data_tl_r_101_sv2v_reg,
  data_tl_r_100_sv2v_reg,data_tl_r_99_sv2v_reg,data_tl_r_98_sv2v_reg,data_tl_r_97_sv2v_reg,
  data_tl_r_96_sv2v_reg,data_tl_r_95_sv2v_reg,data_tl_r_94_sv2v_reg,data_tl_r_93_sv2v_reg,
  data_tl_r_92_sv2v_reg,data_tl_r_91_sv2v_reg,data_tl_r_90_sv2v_reg,
  data_tl_r_89_sv2v_reg,data_tl_r_88_sv2v_reg,data_tl_r_87_sv2v_reg,data_tl_r_86_sv2v_reg,
  data_tl_r_85_sv2v_reg,data_tl_r_84_sv2v_reg,data_tl_r_83_sv2v_reg,data_tl_r_82_sv2v_reg,
  data_tl_r_81_sv2v_reg,data_tl_r_80_sv2v_reg,data_tl_r_79_sv2v_reg,
  data_tl_r_78_sv2v_reg,data_tl_r_77_sv2v_reg,data_tl_r_76_sv2v_reg,data_tl_r_75_sv2v_reg,
  data_tl_r_74_sv2v_reg,data_tl_r_73_sv2v_reg,data_tl_r_72_sv2v_reg,
  data_tl_r_71_sv2v_reg,data_tl_r_70_sv2v_reg,data_tl_r_69_sv2v_reg,data_tl_r_68_sv2v_reg,
  data_tl_r_67_sv2v_reg,data_tl_r_66_sv2v_reg,data_tl_r_65_sv2v_reg,data_tl_r_64_sv2v_reg,
  data_tl_r_63_sv2v_reg,data_tl_r_62_sv2v_reg,data_tl_r_61_sv2v_reg,
  data_tl_r_60_sv2v_reg,data_tl_r_59_sv2v_reg,data_tl_r_58_sv2v_reg,data_tl_r_57_sv2v_reg,
  data_tl_r_56_sv2v_reg,data_tl_r_55_sv2v_reg,data_tl_r_54_sv2v_reg,data_tl_r_53_sv2v_reg,
  data_tl_r_52_sv2v_reg,data_tl_r_51_sv2v_reg,data_tl_r_50_sv2v_reg,
  data_tl_r_49_sv2v_reg,data_tl_r_48_sv2v_reg,data_tl_r_47_sv2v_reg,data_tl_r_46_sv2v_reg,
  data_tl_r_45_sv2v_reg,data_tl_r_44_sv2v_reg,data_tl_r_43_sv2v_reg,data_tl_r_42_sv2v_reg,
  data_tl_r_41_sv2v_reg,data_tl_r_40_sv2v_reg,data_tl_r_39_sv2v_reg,
  data_tl_r_38_sv2v_reg,data_tl_r_37_sv2v_reg,data_tl_r_36_sv2v_reg,data_tl_r_35_sv2v_reg,
  data_tl_r_34_sv2v_reg,data_tl_r_33_sv2v_reg,data_tl_r_32_sv2v_reg,
  data_tl_r_31_sv2v_reg,data_tl_r_30_sv2v_reg,data_tl_r_29_sv2v_reg,data_tl_r_28_sv2v_reg,
  data_tl_r_27_sv2v_reg,data_tl_r_26_sv2v_reg,data_tl_r_25_sv2v_reg,data_tl_r_24_sv2v_reg,
  data_tl_r_23_sv2v_reg,data_tl_r_22_sv2v_reg,data_tl_r_21_sv2v_reg,
  data_tl_r_20_sv2v_reg,data_tl_r_19_sv2v_reg,data_tl_r_18_sv2v_reg,data_tl_r_17_sv2v_reg,
  data_tl_r_16_sv2v_reg,data_tl_r_15_sv2v_reg,data_tl_r_14_sv2v_reg,data_tl_r_13_sv2v_reg,
  data_tl_r_12_sv2v_reg,data_tl_r_11_sv2v_reg,data_tl_r_10_sv2v_reg,
  data_tl_r_9_sv2v_reg,data_tl_r_8_sv2v_reg,data_tl_r_7_sv2v_reg,data_tl_r_6_sv2v_reg,
  data_tl_r_5_sv2v_reg,data_tl_r_4_sv2v_reg,data_tl_r_3_sv2v_reg,data_tl_r_2_sv2v_reg,
  data_tl_r_1_sv2v_reg,data_tl_r_0_sv2v_reg,v_tl_r_sv2v_reg,decode_tl_r_20_sv2v_reg,
  decode_tl_r_19_sv2v_reg,decode_tl_r_18_sv2v_reg,decode_tl_r_17_sv2v_reg,
  decode_tl_r_16_sv2v_reg,decode_tl_r_15_sv2v_reg,decode_tl_r_14_sv2v_reg,
  decode_tl_r_13_sv2v_reg,decode_tl_r_12_sv2v_reg,decode_tl_r_11_sv2v_reg,decode_tl_r_10_sv2v_reg,
  decode_tl_r_9_sv2v_reg,decode_tl_r_8_sv2v_reg,decode_tl_r_7_sv2v_reg,
  decode_tl_r_6_sv2v_reg,decode_tl_r_5_sv2v_reg,decode_tl_r_4_sv2v_reg,decode_tl_r_3_sv2v_reg,
  decode_tl_r_2_sv2v_reg,decode_tl_r_1_sv2v_reg,decode_tl_r_0_sv2v_reg,
  mask_tl_r_15_sv2v_reg,mask_tl_r_14_sv2v_reg,mask_tl_r_13_sv2v_reg,mask_tl_r_12_sv2v_reg,
  mask_tl_r_11_sv2v_reg,mask_tl_r_10_sv2v_reg,mask_tl_r_9_sv2v_reg,mask_tl_r_8_sv2v_reg,
  mask_tl_r_7_sv2v_reg,mask_tl_r_6_sv2v_reg,mask_tl_r_5_sv2v_reg,
  mask_tl_r_4_sv2v_reg,mask_tl_r_3_sv2v_reg,mask_tl_r_2_sv2v_reg,mask_tl_r_1_sv2v_reg,
  mask_tl_r_0_sv2v_reg,addr_tl_r_32_sv2v_reg,addr_tl_r_31_sv2v_reg,addr_tl_r_30_sv2v_reg,
  addr_tl_r_29_sv2v_reg,addr_tl_r_28_sv2v_reg,addr_tl_r_27_sv2v_reg,addr_tl_r_26_sv2v_reg,
  addr_tl_r_25_sv2v_reg,addr_tl_r_24_sv2v_reg,addr_tl_r_23_sv2v_reg,
  addr_tl_r_22_sv2v_reg,addr_tl_r_21_sv2v_reg,addr_tl_r_20_sv2v_reg,addr_tl_r_19_sv2v_reg,
  addr_tl_r_18_sv2v_reg,addr_tl_r_17_sv2v_reg,addr_tl_r_16_sv2v_reg,
  addr_tl_r_15_sv2v_reg,addr_tl_r_14_sv2v_reg,addr_tl_r_13_sv2v_reg,addr_tl_r_12_sv2v_reg,
  addr_tl_r_11_sv2v_reg,addr_tl_r_10_sv2v_reg,addr_tl_r_9_sv2v_reg,addr_tl_r_8_sv2v_reg,
  addr_tl_r_7_sv2v_reg,addr_tl_r_6_sv2v_reg,addr_tl_r_5_sv2v_reg,addr_tl_r_4_sv2v_reg,
  addr_tl_r_3_sv2v_reg,addr_tl_r_2_sv2v_reg,addr_tl_r_1_sv2v_reg,
  addr_tl_r_0_sv2v_reg,ld_data_v_r_1023_sv2v_reg,ld_data_v_r_1022_sv2v_reg,ld_data_v_r_1021_sv2v_reg,
  ld_data_v_r_1020_sv2v_reg,ld_data_v_r_1019_sv2v_reg,ld_data_v_r_1018_sv2v_reg,
  ld_data_v_r_1017_sv2v_reg,ld_data_v_r_1016_sv2v_reg,ld_data_v_r_1015_sv2v_reg,
  ld_data_v_r_1014_sv2v_reg,ld_data_v_r_1013_sv2v_reg,ld_data_v_r_1012_sv2v_reg,
  ld_data_v_r_1011_sv2v_reg,ld_data_v_r_1010_sv2v_reg,ld_data_v_r_1009_sv2v_reg,
  ld_data_v_r_1008_sv2v_reg,ld_data_v_r_1007_sv2v_reg,ld_data_v_r_1006_sv2v_reg,
  ld_data_v_r_1005_sv2v_reg,ld_data_v_r_1004_sv2v_reg,ld_data_v_r_1003_sv2v_reg,
  ld_data_v_r_1002_sv2v_reg,ld_data_v_r_1001_sv2v_reg,ld_data_v_r_1000_sv2v_reg,
  ld_data_v_r_999_sv2v_reg,ld_data_v_r_998_sv2v_reg,ld_data_v_r_997_sv2v_reg,
  ld_data_v_r_996_sv2v_reg,ld_data_v_r_995_sv2v_reg,ld_data_v_r_994_sv2v_reg,
  ld_data_v_r_993_sv2v_reg,ld_data_v_r_992_sv2v_reg,ld_data_v_r_991_sv2v_reg,ld_data_v_r_990_sv2v_reg,
  ld_data_v_r_989_sv2v_reg,ld_data_v_r_988_sv2v_reg,ld_data_v_r_987_sv2v_reg,
  ld_data_v_r_986_sv2v_reg,ld_data_v_r_985_sv2v_reg,ld_data_v_r_984_sv2v_reg,
  ld_data_v_r_983_sv2v_reg,ld_data_v_r_982_sv2v_reg,ld_data_v_r_981_sv2v_reg,
  ld_data_v_r_980_sv2v_reg,ld_data_v_r_979_sv2v_reg,ld_data_v_r_978_sv2v_reg,
  ld_data_v_r_977_sv2v_reg,ld_data_v_r_976_sv2v_reg,ld_data_v_r_975_sv2v_reg,ld_data_v_r_974_sv2v_reg,
  ld_data_v_r_973_sv2v_reg,ld_data_v_r_972_sv2v_reg,ld_data_v_r_971_sv2v_reg,
  ld_data_v_r_970_sv2v_reg,ld_data_v_r_969_sv2v_reg,ld_data_v_r_968_sv2v_reg,
  ld_data_v_r_967_sv2v_reg,ld_data_v_r_966_sv2v_reg,ld_data_v_r_965_sv2v_reg,
  ld_data_v_r_964_sv2v_reg,ld_data_v_r_963_sv2v_reg,ld_data_v_r_962_sv2v_reg,
  ld_data_v_r_961_sv2v_reg,ld_data_v_r_960_sv2v_reg,ld_data_v_r_959_sv2v_reg,ld_data_v_r_958_sv2v_reg,
  ld_data_v_r_957_sv2v_reg,ld_data_v_r_956_sv2v_reg,ld_data_v_r_955_sv2v_reg,
  ld_data_v_r_954_sv2v_reg,ld_data_v_r_953_sv2v_reg,ld_data_v_r_952_sv2v_reg,
  ld_data_v_r_951_sv2v_reg,ld_data_v_r_950_sv2v_reg,ld_data_v_r_949_sv2v_reg,
  ld_data_v_r_948_sv2v_reg,ld_data_v_r_947_sv2v_reg,ld_data_v_r_946_sv2v_reg,
  ld_data_v_r_945_sv2v_reg,ld_data_v_r_944_sv2v_reg,ld_data_v_r_943_sv2v_reg,ld_data_v_r_942_sv2v_reg,
  ld_data_v_r_941_sv2v_reg,ld_data_v_r_940_sv2v_reg,ld_data_v_r_939_sv2v_reg,
  ld_data_v_r_938_sv2v_reg,ld_data_v_r_937_sv2v_reg,ld_data_v_r_936_sv2v_reg,
  ld_data_v_r_935_sv2v_reg,ld_data_v_r_934_sv2v_reg,ld_data_v_r_933_sv2v_reg,
  ld_data_v_r_932_sv2v_reg,ld_data_v_r_931_sv2v_reg,ld_data_v_r_930_sv2v_reg,
  ld_data_v_r_929_sv2v_reg,ld_data_v_r_928_sv2v_reg,ld_data_v_r_927_sv2v_reg,ld_data_v_r_926_sv2v_reg,
  ld_data_v_r_925_sv2v_reg,ld_data_v_r_924_sv2v_reg,ld_data_v_r_923_sv2v_reg,
  ld_data_v_r_922_sv2v_reg,ld_data_v_r_921_sv2v_reg,ld_data_v_r_920_sv2v_reg,
  ld_data_v_r_919_sv2v_reg,ld_data_v_r_918_sv2v_reg,ld_data_v_r_917_sv2v_reg,
  ld_data_v_r_916_sv2v_reg,ld_data_v_r_915_sv2v_reg,ld_data_v_r_914_sv2v_reg,
  ld_data_v_r_913_sv2v_reg,ld_data_v_r_912_sv2v_reg,ld_data_v_r_911_sv2v_reg,ld_data_v_r_910_sv2v_reg,
  ld_data_v_r_909_sv2v_reg,ld_data_v_r_908_sv2v_reg,ld_data_v_r_907_sv2v_reg,
  ld_data_v_r_906_sv2v_reg,ld_data_v_r_905_sv2v_reg,ld_data_v_r_904_sv2v_reg,
  ld_data_v_r_903_sv2v_reg,ld_data_v_r_902_sv2v_reg,ld_data_v_r_901_sv2v_reg,
  ld_data_v_r_900_sv2v_reg,ld_data_v_r_899_sv2v_reg,ld_data_v_r_898_sv2v_reg,
  ld_data_v_r_897_sv2v_reg,ld_data_v_r_896_sv2v_reg,ld_data_v_r_895_sv2v_reg,ld_data_v_r_894_sv2v_reg,
  ld_data_v_r_893_sv2v_reg,ld_data_v_r_892_sv2v_reg,ld_data_v_r_891_sv2v_reg,
  ld_data_v_r_890_sv2v_reg,ld_data_v_r_889_sv2v_reg,ld_data_v_r_888_sv2v_reg,
  ld_data_v_r_887_sv2v_reg,ld_data_v_r_886_sv2v_reg,ld_data_v_r_885_sv2v_reg,
  ld_data_v_r_884_sv2v_reg,ld_data_v_r_883_sv2v_reg,ld_data_v_r_882_sv2v_reg,
  ld_data_v_r_881_sv2v_reg,ld_data_v_r_880_sv2v_reg,ld_data_v_r_879_sv2v_reg,ld_data_v_r_878_sv2v_reg,
  ld_data_v_r_877_sv2v_reg,ld_data_v_r_876_sv2v_reg,ld_data_v_r_875_sv2v_reg,
  ld_data_v_r_874_sv2v_reg,ld_data_v_r_873_sv2v_reg,ld_data_v_r_872_sv2v_reg,
  ld_data_v_r_871_sv2v_reg,ld_data_v_r_870_sv2v_reg,ld_data_v_r_869_sv2v_reg,
  ld_data_v_r_868_sv2v_reg,ld_data_v_r_867_sv2v_reg,ld_data_v_r_866_sv2v_reg,
  ld_data_v_r_865_sv2v_reg,ld_data_v_r_864_sv2v_reg,ld_data_v_r_863_sv2v_reg,ld_data_v_r_862_sv2v_reg,
  ld_data_v_r_861_sv2v_reg,ld_data_v_r_860_sv2v_reg,ld_data_v_r_859_sv2v_reg,
  ld_data_v_r_858_sv2v_reg,ld_data_v_r_857_sv2v_reg,ld_data_v_r_856_sv2v_reg,
  ld_data_v_r_855_sv2v_reg,ld_data_v_r_854_sv2v_reg,ld_data_v_r_853_sv2v_reg,
  ld_data_v_r_852_sv2v_reg,ld_data_v_r_851_sv2v_reg,ld_data_v_r_850_sv2v_reg,
  ld_data_v_r_849_sv2v_reg,ld_data_v_r_848_sv2v_reg,ld_data_v_r_847_sv2v_reg,ld_data_v_r_846_sv2v_reg,
  ld_data_v_r_845_sv2v_reg,ld_data_v_r_844_sv2v_reg,ld_data_v_r_843_sv2v_reg,
  ld_data_v_r_842_sv2v_reg,ld_data_v_r_841_sv2v_reg,ld_data_v_r_840_sv2v_reg,
  ld_data_v_r_839_sv2v_reg,ld_data_v_r_838_sv2v_reg,ld_data_v_r_837_sv2v_reg,
  ld_data_v_r_836_sv2v_reg,ld_data_v_r_835_sv2v_reg,ld_data_v_r_834_sv2v_reg,
  ld_data_v_r_833_sv2v_reg,ld_data_v_r_832_sv2v_reg,ld_data_v_r_831_sv2v_reg,ld_data_v_r_830_sv2v_reg,
  ld_data_v_r_829_sv2v_reg,ld_data_v_r_828_sv2v_reg,ld_data_v_r_827_sv2v_reg,
  ld_data_v_r_826_sv2v_reg,ld_data_v_r_825_sv2v_reg,ld_data_v_r_824_sv2v_reg,
  ld_data_v_r_823_sv2v_reg,ld_data_v_r_822_sv2v_reg,ld_data_v_r_821_sv2v_reg,
  ld_data_v_r_820_sv2v_reg,ld_data_v_r_819_sv2v_reg,ld_data_v_r_818_sv2v_reg,
  ld_data_v_r_817_sv2v_reg,ld_data_v_r_816_sv2v_reg,ld_data_v_r_815_sv2v_reg,ld_data_v_r_814_sv2v_reg,
  ld_data_v_r_813_sv2v_reg,ld_data_v_r_812_sv2v_reg,ld_data_v_r_811_sv2v_reg,
  ld_data_v_r_810_sv2v_reg,ld_data_v_r_809_sv2v_reg,ld_data_v_r_808_sv2v_reg,
  ld_data_v_r_807_sv2v_reg,ld_data_v_r_806_sv2v_reg,ld_data_v_r_805_sv2v_reg,
  ld_data_v_r_804_sv2v_reg,ld_data_v_r_803_sv2v_reg,ld_data_v_r_802_sv2v_reg,
  ld_data_v_r_801_sv2v_reg,ld_data_v_r_800_sv2v_reg,ld_data_v_r_799_sv2v_reg,ld_data_v_r_798_sv2v_reg,
  ld_data_v_r_797_sv2v_reg,ld_data_v_r_796_sv2v_reg,ld_data_v_r_795_sv2v_reg,
  ld_data_v_r_794_sv2v_reg,ld_data_v_r_793_sv2v_reg,ld_data_v_r_792_sv2v_reg,
  ld_data_v_r_791_sv2v_reg,ld_data_v_r_790_sv2v_reg,ld_data_v_r_789_sv2v_reg,
  ld_data_v_r_788_sv2v_reg,ld_data_v_r_787_sv2v_reg,ld_data_v_r_786_sv2v_reg,
  ld_data_v_r_785_sv2v_reg,ld_data_v_r_784_sv2v_reg,ld_data_v_r_783_sv2v_reg,ld_data_v_r_782_sv2v_reg,
  ld_data_v_r_781_sv2v_reg,ld_data_v_r_780_sv2v_reg,ld_data_v_r_779_sv2v_reg,
  ld_data_v_r_778_sv2v_reg,ld_data_v_r_777_sv2v_reg,ld_data_v_r_776_sv2v_reg,
  ld_data_v_r_775_sv2v_reg,ld_data_v_r_774_sv2v_reg,ld_data_v_r_773_sv2v_reg,
  ld_data_v_r_772_sv2v_reg,ld_data_v_r_771_sv2v_reg,ld_data_v_r_770_sv2v_reg,
  ld_data_v_r_769_sv2v_reg,ld_data_v_r_768_sv2v_reg,ld_data_v_r_767_sv2v_reg,ld_data_v_r_766_sv2v_reg,
  ld_data_v_r_765_sv2v_reg,ld_data_v_r_764_sv2v_reg,ld_data_v_r_763_sv2v_reg,
  ld_data_v_r_762_sv2v_reg,ld_data_v_r_761_sv2v_reg,ld_data_v_r_760_sv2v_reg,
  ld_data_v_r_759_sv2v_reg,ld_data_v_r_758_sv2v_reg,ld_data_v_r_757_sv2v_reg,
  ld_data_v_r_756_sv2v_reg,ld_data_v_r_755_sv2v_reg,ld_data_v_r_754_sv2v_reg,
  ld_data_v_r_753_sv2v_reg,ld_data_v_r_752_sv2v_reg,ld_data_v_r_751_sv2v_reg,ld_data_v_r_750_sv2v_reg,
  ld_data_v_r_749_sv2v_reg,ld_data_v_r_748_sv2v_reg,ld_data_v_r_747_sv2v_reg,
  ld_data_v_r_746_sv2v_reg,ld_data_v_r_745_sv2v_reg,ld_data_v_r_744_sv2v_reg,
  ld_data_v_r_743_sv2v_reg,ld_data_v_r_742_sv2v_reg,ld_data_v_r_741_sv2v_reg,
  ld_data_v_r_740_sv2v_reg,ld_data_v_r_739_sv2v_reg,ld_data_v_r_738_sv2v_reg,
  ld_data_v_r_737_sv2v_reg,ld_data_v_r_736_sv2v_reg,ld_data_v_r_735_sv2v_reg,ld_data_v_r_734_sv2v_reg,
  ld_data_v_r_733_sv2v_reg,ld_data_v_r_732_sv2v_reg,ld_data_v_r_731_sv2v_reg,
  ld_data_v_r_730_sv2v_reg,ld_data_v_r_729_sv2v_reg,ld_data_v_r_728_sv2v_reg,
  ld_data_v_r_727_sv2v_reg,ld_data_v_r_726_sv2v_reg,ld_data_v_r_725_sv2v_reg,
  ld_data_v_r_724_sv2v_reg,ld_data_v_r_723_sv2v_reg,ld_data_v_r_722_sv2v_reg,
  ld_data_v_r_721_sv2v_reg,ld_data_v_r_720_sv2v_reg,ld_data_v_r_719_sv2v_reg,ld_data_v_r_718_sv2v_reg,
  ld_data_v_r_717_sv2v_reg,ld_data_v_r_716_sv2v_reg,ld_data_v_r_715_sv2v_reg,
  ld_data_v_r_714_sv2v_reg,ld_data_v_r_713_sv2v_reg,ld_data_v_r_712_sv2v_reg,
  ld_data_v_r_711_sv2v_reg,ld_data_v_r_710_sv2v_reg,ld_data_v_r_709_sv2v_reg,
  ld_data_v_r_708_sv2v_reg,ld_data_v_r_707_sv2v_reg,ld_data_v_r_706_sv2v_reg,
  ld_data_v_r_705_sv2v_reg,ld_data_v_r_704_sv2v_reg,ld_data_v_r_703_sv2v_reg,ld_data_v_r_702_sv2v_reg,
  ld_data_v_r_701_sv2v_reg,ld_data_v_r_700_sv2v_reg,ld_data_v_r_699_sv2v_reg,
  ld_data_v_r_698_sv2v_reg,ld_data_v_r_697_sv2v_reg,ld_data_v_r_696_sv2v_reg,
  ld_data_v_r_695_sv2v_reg,ld_data_v_r_694_sv2v_reg,ld_data_v_r_693_sv2v_reg,
  ld_data_v_r_692_sv2v_reg,ld_data_v_r_691_sv2v_reg,ld_data_v_r_690_sv2v_reg,
  ld_data_v_r_689_sv2v_reg,ld_data_v_r_688_sv2v_reg,ld_data_v_r_687_sv2v_reg,ld_data_v_r_686_sv2v_reg,
  ld_data_v_r_685_sv2v_reg,ld_data_v_r_684_sv2v_reg,ld_data_v_r_683_sv2v_reg,
  ld_data_v_r_682_sv2v_reg,ld_data_v_r_681_sv2v_reg,ld_data_v_r_680_sv2v_reg,
  ld_data_v_r_679_sv2v_reg,ld_data_v_r_678_sv2v_reg,ld_data_v_r_677_sv2v_reg,
  ld_data_v_r_676_sv2v_reg,ld_data_v_r_675_sv2v_reg,ld_data_v_r_674_sv2v_reg,
  ld_data_v_r_673_sv2v_reg,ld_data_v_r_672_sv2v_reg,ld_data_v_r_671_sv2v_reg,ld_data_v_r_670_sv2v_reg,
  ld_data_v_r_669_sv2v_reg,ld_data_v_r_668_sv2v_reg,ld_data_v_r_667_sv2v_reg,
  ld_data_v_r_666_sv2v_reg,ld_data_v_r_665_sv2v_reg,ld_data_v_r_664_sv2v_reg,
  ld_data_v_r_663_sv2v_reg,ld_data_v_r_662_sv2v_reg,ld_data_v_r_661_sv2v_reg,
  ld_data_v_r_660_sv2v_reg,ld_data_v_r_659_sv2v_reg,ld_data_v_r_658_sv2v_reg,
  ld_data_v_r_657_sv2v_reg,ld_data_v_r_656_sv2v_reg,ld_data_v_r_655_sv2v_reg,ld_data_v_r_654_sv2v_reg,
  ld_data_v_r_653_sv2v_reg,ld_data_v_r_652_sv2v_reg,ld_data_v_r_651_sv2v_reg,
  ld_data_v_r_650_sv2v_reg,ld_data_v_r_649_sv2v_reg,ld_data_v_r_648_sv2v_reg,
  ld_data_v_r_647_sv2v_reg,ld_data_v_r_646_sv2v_reg,ld_data_v_r_645_sv2v_reg,
  ld_data_v_r_644_sv2v_reg,ld_data_v_r_643_sv2v_reg,ld_data_v_r_642_sv2v_reg,
  ld_data_v_r_641_sv2v_reg,ld_data_v_r_640_sv2v_reg,ld_data_v_r_639_sv2v_reg,ld_data_v_r_638_sv2v_reg,
  ld_data_v_r_637_sv2v_reg,ld_data_v_r_636_sv2v_reg,ld_data_v_r_635_sv2v_reg,
  ld_data_v_r_634_sv2v_reg,ld_data_v_r_633_sv2v_reg,ld_data_v_r_632_sv2v_reg,
  ld_data_v_r_631_sv2v_reg,ld_data_v_r_630_sv2v_reg,ld_data_v_r_629_sv2v_reg,
  ld_data_v_r_628_sv2v_reg,ld_data_v_r_627_sv2v_reg,ld_data_v_r_626_sv2v_reg,
  ld_data_v_r_625_sv2v_reg,ld_data_v_r_624_sv2v_reg,ld_data_v_r_623_sv2v_reg,ld_data_v_r_622_sv2v_reg,
  ld_data_v_r_621_sv2v_reg,ld_data_v_r_620_sv2v_reg,ld_data_v_r_619_sv2v_reg,
  ld_data_v_r_618_sv2v_reg,ld_data_v_r_617_sv2v_reg,ld_data_v_r_616_sv2v_reg,
  ld_data_v_r_615_sv2v_reg,ld_data_v_r_614_sv2v_reg,ld_data_v_r_613_sv2v_reg,
  ld_data_v_r_612_sv2v_reg,ld_data_v_r_611_sv2v_reg,ld_data_v_r_610_sv2v_reg,
  ld_data_v_r_609_sv2v_reg,ld_data_v_r_608_sv2v_reg,ld_data_v_r_607_sv2v_reg,ld_data_v_r_606_sv2v_reg,
  ld_data_v_r_605_sv2v_reg,ld_data_v_r_604_sv2v_reg,ld_data_v_r_603_sv2v_reg,
  ld_data_v_r_602_sv2v_reg,ld_data_v_r_601_sv2v_reg,ld_data_v_r_600_sv2v_reg,
  ld_data_v_r_599_sv2v_reg,ld_data_v_r_598_sv2v_reg,ld_data_v_r_597_sv2v_reg,
  ld_data_v_r_596_sv2v_reg,ld_data_v_r_595_sv2v_reg,ld_data_v_r_594_sv2v_reg,
  ld_data_v_r_593_sv2v_reg,ld_data_v_r_592_sv2v_reg,ld_data_v_r_591_sv2v_reg,ld_data_v_r_590_sv2v_reg,
  ld_data_v_r_589_sv2v_reg,ld_data_v_r_588_sv2v_reg,ld_data_v_r_587_sv2v_reg,
  ld_data_v_r_586_sv2v_reg,ld_data_v_r_585_sv2v_reg,ld_data_v_r_584_sv2v_reg,
  ld_data_v_r_583_sv2v_reg,ld_data_v_r_582_sv2v_reg,ld_data_v_r_581_sv2v_reg,
  ld_data_v_r_580_sv2v_reg,ld_data_v_r_579_sv2v_reg,ld_data_v_r_578_sv2v_reg,
  ld_data_v_r_577_sv2v_reg,ld_data_v_r_576_sv2v_reg,ld_data_v_r_575_sv2v_reg,ld_data_v_r_574_sv2v_reg,
  ld_data_v_r_573_sv2v_reg,ld_data_v_r_572_sv2v_reg,ld_data_v_r_571_sv2v_reg,
  ld_data_v_r_570_sv2v_reg,ld_data_v_r_569_sv2v_reg,ld_data_v_r_568_sv2v_reg,
  ld_data_v_r_567_sv2v_reg,ld_data_v_r_566_sv2v_reg,ld_data_v_r_565_sv2v_reg,
  ld_data_v_r_564_sv2v_reg,ld_data_v_r_563_sv2v_reg,ld_data_v_r_562_sv2v_reg,
  ld_data_v_r_561_sv2v_reg,ld_data_v_r_560_sv2v_reg,ld_data_v_r_559_sv2v_reg,ld_data_v_r_558_sv2v_reg,
  ld_data_v_r_557_sv2v_reg,ld_data_v_r_556_sv2v_reg,ld_data_v_r_555_sv2v_reg,
  ld_data_v_r_554_sv2v_reg,ld_data_v_r_553_sv2v_reg,ld_data_v_r_552_sv2v_reg,
  ld_data_v_r_551_sv2v_reg,ld_data_v_r_550_sv2v_reg,ld_data_v_r_549_sv2v_reg,
  ld_data_v_r_548_sv2v_reg,ld_data_v_r_547_sv2v_reg,ld_data_v_r_546_sv2v_reg,
  ld_data_v_r_545_sv2v_reg,ld_data_v_r_544_sv2v_reg,ld_data_v_r_543_sv2v_reg,ld_data_v_r_542_sv2v_reg,
  ld_data_v_r_541_sv2v_reg,ld_data_v_r_540_sv2v_reg,ld_data_v_r_539_sv2v_reg,
  ld_data_v_r_538_sv2v_reg,ld_data_v_r_537_sv2v_reg,ld_data_v_r_536_sv2v_reg,
  ld_data_v_r_535_sv2v_reg,ld_data_v_r_534_sv2v_reg,ld_data_v_r_533_sv2v_reg,
  ld_data_v_r_532_sv2v_reg,ld_data_v_r_531_sv2v_reg,ld_data_v_r_530_sv2v_reg,
  ld_data_v_r_529_sv2v_reg,ld_data_v_r_528_sv2v_reg,ld_data_v_r_527_sv2v_reg,ld_data_v_r_526_sv2v_reg,
  ld_data_v_r_525_sv2v_reg,ld_data_v_r_524_sv2v_reg,ld_data_v_r_523_sv2v_reg,
  ld_data_v_r_522_sv2v_reg,ld_data_v_r_521_sv2v_reg,ld_data_v_r_520_sv2v_reg,
  ld_data_v_r_519_sv2v_reg,ld_data_v_r_518_sv2v_reg,ld_data_v_r_517_sv2v_reg,
  ld_data_v_r_516_sv2v_reg,ld_data_v_r_515_sv2v_reg,ld_data_v_r_514_sv2v_reg,
  ld_data_v_r_513_sv2v_reg,ld_data_v_r_512_sv2v_reg,ld_data_v_r_511_sv2v_reg,ld_data_v_r_510_sv2v_reg,
  ld_data_v_r_509_sv2v_reg,ld_data_v_r_508_sv2v_reg,ld_data_v_r_507_sv2v_reg,
  ld_data_v_r_506_sv2v_reg,ld_data_v_r_505_sv2v_reg,ld_data_v_r_504_sv2v_reg,
  ld_data_v_r_503_sv2v_reg,ld_data_v_r_502_sv2v_reg,ld_data_v_r_501_sv2v_reg,
  ld_data_v_r_500_sv2v_reg,ld_data_v_r_499_sv2v_reg,ld_data_v_r_498_sv2v_reg,
  ld_data_v_r_497_sv2v_reg,ld_data_v_r_496_sv2v_reg,ld_data_v_r_495_sv2v_reg,ld_data_v_r_494_sv2v_reg,
  ld_data_v_r_493_sv2v_reg,ld_data_v_r_492_sv2v_reg,ld_data_v_r_491_sv2v_reg,
  ld_data_v_r_490_sv2v_reg,ld_data_v_r_489_sv2v_reg,ld_data_v_r_488_sv2v_reg,
  ld_data_v_r_487_sv2v_reg,ld_data_v_r_486_sv2v_reg,ld_data_v_r_485_sv2v_reg,
  ld_data_v_r_484_sv2v_reg,ld_data_v_r_483_sv2v_reg,ld_data_v_r_482_sv2v_reg,
  ld_data_v_r_481_sv2v_reg,ld_data_v_r_480_sv2v_reg,ld_data_v_r_479_sv2v_reg,ld_data_v_r_478_sv2v_reg,
  ld_data_v_r_477_sv2v_reg,ld_data_v_r_476_sv2v_reg,ld_data_v_r_475_sv2v_reg,
  ld_data_v_r_474_sv2v_reg,ld_data_v_r_473_sv2v_reg,ld_data_v_r_472_sv2v_reg,
  ld_data_v_r_471_sv2v_reg,ld_data_v_r_470_sv2v_reg,ld_data_v_r_469_sv2v_reg,
  ld_data_v_r_468_sv2v_reg,ld_data_v_r_467_sv2v_reg,ld_data_v_r_466_sv2v_reg,
  ld_data_v_r_465_sv2v_reg,ld_data_v_r_464_sv2v_reg,ld_data_v_r_463_sv2v_reg,ld_data_v_r_462_sv2v_reg,
  ld_data_v_r_461_sv2v_reg,ld_data_v_r_460_sv2v_reg,ld_data_v_r_459_sv2v_reg,
  ld_data_v_r_458_sv2v_reg,ld_data_v_r_457_sv2v_reg,ld_data_v_r_456_sv2v_reg,
  ld_data_v_r_455_sv2v_reg,ld_data_v_r_454_sv2v_reg,ld_data_v_r_453_sv2v_reg,
  ld_data_v_r_452_sv2v_reg,ld_data_v_r_451_sv2v_reg,ld_data_v_r_450_sv2v_reg,
  ld_data_v_r_449_sv2v_reg,ld_data_v_r_448_sv2v_reg,ld_data_v_r_447_sv2v_reg,ld_data_v_r_446_sv2v_reg,
  ld_data_v_r_445_sv2v_reg,ld_data_v_r_444_sv2v_reg,ld_data_v_r_443_sv2v_reg,
  ld_data_v_r_442_sv2v_reg,ld_data_v_r_441_sv2v_reg,ld_data_v_r_440_sv2v_reg,
  ld_data_v_r_439_sv2v_reg,ld_data_v_r_438_sv2v_reg,ld_data_v_r_437_sv2v_reg,
  ld_data_v_r_436_sv2v_reg,ld_data_v_r_435_sv2v_reg,ld_data_v_r_434_sv2v_reg,
  ld_data_v_r_433_sv2v_reg,ld_data_v_r_432_sv2v_reg,ld_data_v_r_431_sv2v_reg,ld_data_v_r_430_sv2v_reg,
  ld_data_v_r_429_sv2v_reg,ld_data_v_r_428_sv2v_reg,ld_data_v_r_427_sv2v_reg,
  ld_data_v_r_426_sv2v_reg,ld_data_v_r_425_sv2v_reg,ld_data_v_r_424_sv2v_reg,
  ld_data_v_r_423_sv2v_reg,ld_data_v_r_422_sv2v_reg,ld_data_v_r_421_sv2v_reg,
  ld_data_v_r_420_sv2v_reg,ld_data_v_r_419_sv2v_reg,ld_data_v_r_418_sv2v_reg,
  ld_data_v_r_417_sv2v_reg,ld_data_v_r_416_sv2v_reg,ld_data_v_r_415_sv2v_reg,ld_data_v_r_414_sv2v_reg,
  ld_data_v_r_413_sv2v_reg,ld_data_v_r_412_sv2v_reg,ld_data_v_r_411_sv2v_reg,
  ld_data_v_r_410_sv2v_reg,ld_data_v_r_409_sv2v_reg,ld_data_v_r_408_sv2v_reg,
  ld_data_v_r_407_sv2v_reg,ld_data_v_r_406_sv2v_reg,ld_data_v_r_405_sv2v_reg,
  ld_data_v_r_404_sv2v_reg,ld_data_v_r_403_sv2v_reg,ld_data_v_r_402_sv2v_reg,
  ld_data_v_r_401_sv2v_reg,ld_data_v_r_400_sv2v_reg,ld_data_v_r_399_sv2v_reg,ld_data_v_r_398_sv2v_reg,
  ld_data_v_r_397_sv2v_reg,ld_data_v_r_396_sv2v_reg,ld_data_v_r_395_sv2v_reg,
  ld_data_v_r_394_sv2v_reg,ld_data_v_r_393_sv2v_reg,ld_data_v_r_392_sv2v_reg,
  ld_data_v_r_391_sv2v_reg,ld_data_v_r_390_sv2v_reg,ld_data_v_r_389_sv2v_reg,
  ld_data_v_r_388_sv2v_reg,ld_data_v_r_387_sv2v_reg,ld_data_v_r_386_sv2v_reg,
  ld_data_v_r_385_sv2v_reg,ld_data_v_r_384_sv2v_reg,ld_data_v_r_383_sv2v_reg,ld_data_v_r_382_sv2v_reg,
  ld_data_v_r_381_sv2v_reg,ld_data_v_r_380_sv2v_reg,ld_data_v_r_379_sv2v_reg,
  ld_data_v_r_378_sv2v_reg,ld_data_v_r_377_sv2v_reg,ld_data_v_r_376_sv2v_reg,
  ld_data_v_r_375_sv2v_reg,ld_data_v_r_374_sv2v_reg,ld_data_v_r_373_sv2v_reg,
  ld_data_v_r_372_sv2v_reg,ld_data_v_r_371_sv2v_reg,ld_data_v_r_370_sv2v_reg,
  ld_data_v_r_369_sv2v_reg,ld_data_v_r_368_sv2v_reg,ld_data_v_r_367_sv2v_reg,ld_data_v_r_366_sv2v_reg,
  ld_data_v_r_365_sv2v_reg,ld_data_v_r_364_sv2v_reg,ld_data_v_r_363_sv2v_reg,
  ld_data_v_r_362_sv2v_reg,ld_data_v_r_361_sv2v_reg,ld_data_v_r_360_sv2v_reg,
  ld_data_v_r_359_sv2v_reg,ld_data_v_r_358_sv2v_reg,ld_data_v_r_357_sv2v_reg,
  ld_data_v_r_356_sv2v_reg,ld_data_v_r_355_sv2v_reg,ld_data_v_r_354_sv2v_reg,
  ld_data_v_r_353_sv2v_reg,ld_data_v_r_352_sv2v_reg,ld_data_v_r_351_sv2v_reg,ld_data_v_r_350_sv2v_reg,
  ld_data_v_r_349_sv2v_reg,ld_data_v_r_348_sv2v_reg,ld_data_v_r_347_sv2v_reg,
  ld_data_v_r_346_sv2v_reg,ld_data_v_r_345_sv2v_reg,ld_data_v_r_344_sv2v_reg,
  ld_data_v_r_343_sv2v_reg,ld_data_v_r_342_sv2v_reg,ld_data_v_r_341_sv2v_reg,
  ld_data_v_r_340_sv2v_reg,ld_data_v_r_339_sv2v_reg,ld_data_v_r_338_sv2v_reg,
  ld_data_v_r_337_sv2v_reg,ld_data_v_r_336_sv2v_reg,ld_data_v_r_335_sv2v_reg,ld_data_v_r_334_sv2v_reg,
  ld_data_v_r_333_sv2v_reg,ld_data_v_r_332_sv2v_reg,ld_data_v_r_331_sv2v_reg,
  ld_data_v_r_330_sv2v_reg,ld_data_v_r_329_sv2v_reg,ld_data_v_r_328_sv2v_reg,
  ld_data_v_r_327_sv2v_reg,ld_data_v_r_326_sv2v_reg,ld_data_v_r_325_sv2v_reg,
  ld_data_v_r_324_sv2v_reg,ld_data_v_r_323_sv2v_reg,ld_data_v_r_322_sv2v_reg,
  ld_data_v_r_321_sv2v_reg,ld_data_v_r_320_sv2v_reg,ld_data_v_r_319_sv2v_reg,ld_data_v_r_318_sv2v_reg,
  ld_data_v_r_317_sv2v_reg,ld_data_v_r_316_sv2v_reg,ld_data_v_r_315_sv2v_reg,
  ld_data_v_r_314_sv2v_reg,ld_data_v_r_313_sv2v_reg,ld_data_v_r_312_sv2v_reg,
  ld_data_v_r_311_sv2v_reg,ld_data_v_r_310_sv2v_reg,ld_data_v_r_309_sv2v_reg,
  ld_data_v_r_308_sv2v_reg,ld_data_v_r_307_sv2v_reg,ld_data_v_r_306_sv2v_reg,
  ld_data_v_r_305_sv2v_reg,ld_data_v_r_304_sv2v_reg,ld_data_v_r_303_sv2v_reg,ld_data_v_r_302_sv2v_reg,
  ld_data_v_r_301_sv2v_reg,ld_data_v_r_300_sv2v_reg,ld_data_v_r_299_sv2v_reg,
  ld_data_v_r_298_sv2v_reg,ld_data_v_r_297_sv2v_reg,ld_data_v_r_296_sv2v_reg,
  ld_data_v_r_295_sv2v_reg,ld_data_v_r_294_sv2v_reg,ld_data_v_r_293_sv2v_reg,
  ld_data_v_r_292_sv2v_reg,ld_data_v_r_291_sv2v_reg,ld_data_v_r_290_sv2v_reg,
  ld_data_v_r_289_sv2v_reg,ld_data_v_r_288_sv2v_reg,ld_data_v_r_287_sv2v_reg,ld_data_v_r_286_sv2v_reg,
  ld_data_v_r_285_sv2v_reg,ld_data_v_r_284_sv2v_reg,ld_data_v_r_283_sv2v_reg,
  ld_data_v_r_282_sv2v_reg,ld_data_v_r_281_sv2v_reg,ld_data_v_r_280_sv2v_reg,
  ld_data_v_r_279_sv2v_reg,ld_data_v_r_278_sv2v_reg,ld_data_v_r_277_sv2v_reg,
  ld_data_v_r_276_sv2v_reg,ld_data_v_r_275_sv2v_reg,ld_data_v_r_274_sv2v_reg,
  ld_data_v_r_273_sv2v_reg,ld_data_v_r_272_sv2v_reg,ld_data_v_r_271_sv2v_reg,ld_data_v_r_270_sv2v_reg,
  ld_data_v_r_269_sv2v_reg,ld_data_v_r_268_sv2v_reg,ld_data_v_r_267_sv2v_reg,
  ld_data_v_r_266_sv2v_reg,ld_data_v_r_265_sv2v_reg,ld_data_v_r_264_sv2v_reg,
  ld_data_v_r_263_sv2v_reg,ld_data_v_r_262_sv2v_reg,ld_data_v_r_261_sv2v_reg,
  ld_data_v_r_260_sv2v_reg,ld_data_v_r_259_sv2v_reg,ld_data_v_r_258_sv2v_reg,
  ld_data_v_r_257_sv2v_reg,ld_data_v_r_256_sv2v_reg,ld_data_v_r_255_sv2v_reg,ld_data_v_r_254_sv2v_reg,
  ld_data_v_r_253_sv2v_reg,ld_data_v_r_252_sv2v_reg,ld_data_v_r_251_sv2v_reg,
  ld_data_v_r_250_sv2v_reg,ld_data_v_r_249_sv2v_reg,ld_data_v_r_248_sv2v_reg,
  ld_data_v_r_247_sv2v_reg,ld_data_v_r_246_sv2v_reg,ld_data_v_r_245_sv2v_reg,
  ld_data_v_r_244_sv2v_reg,ld_data_v_r_243_sv2v_reg,ld_data_v_r_242_sv2v_reg,
  ld_data_v_r_241_sv2v_reg,ld_data_v_r_240_sv2v_reg,ld_data_v_r_239_sv2v_reg,ld_data_v_r_238_sv2v_reg,
  ld_data_v_r_237_sv2v_reg,ld_data_v_r_236_sv2v_reg,ld_data_v_r_235_sv2v_reg,
  ld_data_v_r_234_sv2v_reg,ld_data_v_r_233_sv2v_reg,ld_data_v_r_232_sv2v_reg,
  ld_data_v_r_231_sv2v_reg,ld_data_v_r_230_sv2v_reg,ld_data_v_r_229_sv2v_reg,
  ld_data_v_r_228_sv2v_reg,ld_data_v_r_227_sv2v_reg,ld_data_v_r_226_sv2v_reg,
  ld_data_v_r_225_sv2v_reg,ld_data_v_r_224_sv2v_reg,ld_data_v_r_223_sv2v_reg,ld_data_v_r_222_sv2v_reg,
  ld_data_v_r_221_sv2v_reg,ld_data_v_r_220_sv2v_reg,ld_data_v_r_219_sv2v_reg,
  ld_data_v_r_218_sv2v_reg,ld_data_v_r_217_sv2v_reg,ld_data_v_r_216_sv2v_reg,
  ld_data_v_r_215_sv2v_reg,ld_data_v_r_214_sv2v_reg,ld_data_v_r_213_sv2v_reg,
  ld_data_v_r_212_sv2v_reg,ld_data_v_r_211_sv2v_reg,ld_data_v_r_210_sv2v_reg,
  ld_data_v_r_209_sv2v_reg,ld_data_v_r_208_sv2v_reg,ld_data_v_r_207_sv2v_reg,ld_data_v_r_206_sv2v_reg,
  ld_data_v_r_205_sv2v_reg,ld_data_v_r_204_sv2v_reg,ld_data_v_r_203_sv2v_reg,
  ld_data_v_r_202_sv2v_reg,ld_data_v_r_201_sv2v_reg,ld_data_v_r_200_sv2v_reg,
  ld_data_v_r_199_sv2v_reg,ld_data_v_r_198_sv2v_reg,ld_data_v_r_197_sv2v_reg,
  ld_data_v_r_196_sv2v_reg,ld_data_v_r_195_sv2v_reg,ld_data_v_r_194_sv2v_reg,
  ld_data_v_r_193_sv2v_reg,ld_data_v_r_192_sv2v_reg,ld_data_v_r_191_sv2v_reg,ld_data_v_r_190_sv2v_reg,
  ld_data_v_r_189_sv2v_reg,ld_data_v_r_188_sv2v_reg,ld_data_v_r_187_sv2v_reg,
  ld_data_v_r_186_sv2v_reg,ld_data_v_r_185_sv2v_reg,ld_data_v_r_184_sv2v_reg,
  ld_data_v_r_183_sv2v_reg,ld_data_v_r_182_sv2v_reg,ld_data_v_r_181_sv2v_reg,
  ld_data_v_r_180_sv2v_reg,ld_data_v_r_179_sv2v_reg,ld_data_v_r_178_sv2v_reg,
  ld_data_v_r_177_sv2v_reg,ld_data_v_r_176_sv2v_reg,ld_data_v_r_175_sv2v_reg,ld_data_v_r_174_sv2v_reg,
  ld_data_v_r_173_sv2v_reg,ld_data_v_r_172_sv2v_reg,ld_data_v_r_171_sv2v_reg,
  ld_data_v_r_170_sv2v_reg,ld_data_v_r_169_sv2v_reg,ld_data_v_r_168_sv2v_reg,
  ld_data_v_r_167_sv2v_reg,ld_data_v_r_166_sv2v_reg,ld_data_v_r_165_sv2v_reg,
  ld_data_v_r_164_sv2v_reg,ld_data_v_r_163_sv2v_reg,ld_data_v_r_162_sv2v_reg,
  ld_data_v_r_161_sv2v_reg,ld_data_v_r_160_sv2v_reg,ld_data_v_r_159_sv2v_reg,ld_data_v_r_158_sv2v_reg,
  ld_data_v_r_157_sv2v_reg,ld_data_v_r_156_sv2v_reg,ld_data_v_r_155_sv2v_reg,
  ld_data_v_r_154_sv2v_reg,ld_data_v_r_153_sv2v_reg,ld_data_v_r_152_sv2v_reg,
  ld_data_v_r_151_sv2v_reg,ld_data_v_r_150_sv2v_reg,ld_data_v_r_149_sv2v_reg,
  ld_data_v_r_148_sv2v_reg,ld_data_v_r_147_sv2v_reg,ld_data_v_r_146_sv2v_reg,
  ld_data_v_r_145_sv2v_reg,ld_data_v_r_144_sv2v_reg,ld_data_v_r_143_sv2v_reg,ld_data_v_r_142_sv2v_reg,
  ld_data_v_r_141_sv2v_reg,ld_data_v_r_140_sv2v_reg,ld_data_v_r_139_sv2v_reg,
  ld_data_v_r_138_sv2v_reg,ld_data_v_r_137_sv2v_reg,ld_data_v_r_136_sv2v_reg,
  ld_data_v_r_135_sv2v_reg,ld_data_v_r_134_sv2v_reg,ld_data_v_r_133_sv2v_reg,
  ld_data_v_r_132_sv2v_reg,ld_data_v_r_131_sv2v_reg,ld_data_v_r_130_sv2v_reg,
  ld_data_v_r_129_sv2v_reg,ld_data_v_r_128_sv2v_reg,ld_data_v_r_127_sv2v_reg,ld_data_v_r_126_sv2v_reg,
  ld_data_v_r_125_sv2v_reg,ld_data_v_r_124_sv2v_reg,ld_data_v_r_123_sv2v_reg,
  ld_data_v_r_122_sv2v_reg,ld_data_v_r_121_sv2v_reg,ld_data_v_r_120_sv2v_reg,
  ld_data_v_r_119_sv2v_reg,ld_data_v_r_118_sv2v_reg,ld_data_v_r_117_sv2v_reg,
  ld_data_v_r_116_sv2v_reg,ld_data_v_r_115_sv2v_reg,ld_data_v_r_114_sv2v_reg,
  ld_data_v_r_113_sv2v_reg,ld_data_v_r_112_sv2v_reg,ld_data_v_r_111_sv2v_reg,ld_data_v_r_110_sv2v_reg,
  ld_data_v_r_109_sv2v_reg,ld_data_v_r_108_sv2v_reg,ld_data_v_r_107_sv2v_reg,
  ld_data_v_r_106_sv2v_reg,ld_data_v_r_105_sv2v_reg,ld_data_v_r_104_sv2v_reg,
  ld_data_v_r_103_sv2v_reg,ld_data_v_r_102_sv2v_reg,ld_data_v_r_101_sv2v_reg,
  ld_data_v_r_100_sv2v_reg,ld_data_v_r_99_sv2v_reg,ld_data_v_r_98_sv2v_reg,ld_data_v_r_97_sv2v_reg,
  ld_data_v_r_96_sv2v_reg,ld_data_v_r_95_sv2v_reg,ld_data_v_r_94_sv2v_reg,
  ld_data_v_r_93_sv2v_reg,ld_data_v_r_92_sv2v_reg,ld_data_v_r_91_sv2v_reg,
  ld_data_v_r_90_sv2v_reg,ld_data_v_r_89_sv2v_reg,ld_data_v_r_88_sv2v_reg,ld_data_v_r_87_sv2v_reg,
  ld_data_v_r_86_sv2v_reg,ld_data_v_r_85_sv2v_reg,ld_data_v_r_84_sv2v_reg,
  ld_data_v_r_83_sv2v_reg,ld_data_v_r_82_sv2v_reg,ld_data_v_r_81_sv2v_reg,
  ld_data_v_r_80_sv2v_reg,ld_data_v_r_79_sv2v_reg,ld_data_v_r_78_sv2v_reg,ld_data_v_r_77_sv2v_reg,
  ld_data_v_r_76_sv2v_reg,ld_data_v_r_75_sv2v_reg,ld_data_v_r_74_sv2v_reg,
  ld_data_v_r_73_sv2v_reg,ld_data_v_r_72_sv2v_reg,ld_data_v_r_71_sv2v_reg,
  ld_data_v_r_70_sv2v_reg,ld_data_v_r_69_sv2v_reg,ld_data_v_r_68_sv2v_reg,ld_data_v_r_67_sv2v_reg,
  ld_data_v_r_66_sv2v_reg,ld_data_v_r_65_sv2v_reg,ld_data_v_r_64_sv2v_reg,
  ld_data_v_r_63_sv2v_reg,ld_data_v_r_62_sv2v_reg,ld_data_v_r_61_sv2v_reg,
  ld_data_v_r_60_sv2v_reg,ld_data_v_r_59_sv2v_reg,ld_data_v_r_58_sv2v_reg,ld_data_v_r_57_sv2v_reg,
  ld_data_v_r_56_sv2v_reg,ld_data_v_r_55_sv2v_reg,ld_data_v_r_54_sv2v_reg,
  ld_data_v_r_53_sv2v_reg,ld_data_v_r_52_sv2v_reg,ld_data_v_r_51_sv2v_reg,
  ld_data_v_r_50_sv2v_reg,ld_data_v_r_49_sv2v_reg,ld_data_v_r_48_sv2v_reg,ld_data_v_r_47_sv2v_reg,
  ld_data_v_r_46_sv2v_reg,ld_data_v_r_45_sv2v_reg,ld_data_v_r_44_sv2v_reg,
  ld_data_v_r_43_sv2v_reg,ld_data_v_r_42_sv2v_reg,ld_data_v_r_41_sv2v_reg,
  ld_data_v_r_40_sv2v_reg,ld_data_v_r_39_sv2v_reg,ld_data_v_r_38_sv2v_reg,ld_data_v_r_37_sv2v_reg,
  ld_data_v_r_36_sv2v_reg,ld_data_v_r_35_sv2v_reg,ld_data_v_r_34_sv2v_reg,
  ld_data_v_r_33_sv2v_reg,ld_data_v_r_32_sv2v_reg,ld_data_v_r_31_sv2v_reg,
  ld_data_v_r_30_sv2v_reg,ld_data_v_r_29_sv2v_reg,ld_data_v_r_28_sv2v_reg,ld_data_v_r_27_sv2v_reg,
  ld_data_v_r_26_sv2v_reg,ld_data_v_r_25_sv2v_reg,ld_data_v_r_24_sv2v_reg,
  ld_data_v_r_23_sv2v_reg,ld_data_v_r_22_sv2v_reg,ld_data_v_r_21_sv2v_reg,
  ld_data_v_r_20_sv2v_reg,ld_data_v_r_19_sv2v_reg,ld_data_v_r_18_sv2v_reg,ld_data_v_r_17_sv2v_reg,
  ld_data_v_r_16_sv2v_reg,ld_data_v_r_15_sv2v_reg,ld_data_v_r_14_sv2v_reg,
  ld_data_v_r_13_sv2v_reg,ld_data_v_r_12_sv2v_reg,ld_data_v_r_11_sv2v_reg,
  ld_data_v_r_10_sv2v_reg,ld_data_v_r_9_sv2v_reg,ld_data_v_r_8_sv2v_reg,ld_data_v_r_7_sv2v_reg,
  ld_data_v_r_6_sv2v_reg,ld_data_v_r_5_sv2v_reg,ld_data_v_r_4_sv2v_reg,
  ld_data_v_r_3_sv2v_reg,ld_data_v_r_2_sv2v_reg,ld_data_v_r_1_sv2v_reg,ld_data_v_r_0_sv2v_reg,
  v_v_r_sv2v_reg,track_data_v_r_31_sv2v_reg,track_data_v_r_30_sv2v_reg,
  track_data_v_r_29_sv2v_reg,track_data_v_r_28_sv2v_reg,track_data_v_r_27_sv2v_reg,
  track_data_v_r_26_sv2v_reg,track_data_v_r_25_sv2v_reg,track_data_v_r_24_sv2v_reg,
  track_data_v_r_23_sv2v_reg,track_data_v_r_22_sv2v_reg,track_data_v_r_21_sv2v_reg,
  track_data_v_r_20_sv2v_reg,track_data_v_r_19_sv2v_reg,track_data_v_r_18_sv2v_reg,
  track_data_v_r_17_sv2v_reg,track_data_v_r_16_sv2v_reg,track_data_v_r_15_sv2v_reg,
  track_data_v_r_14_sv2v_reg,track_data_v_r_13_sv2v_reg,track_data_v_r_12_sv2v_reg,
  track_data_v_r_11_sv2v_reg,track_data_v_r_10_sv2v_reg,track_data_v_r_9_sv2v_reg,
  track_data_v_r_8_sv2v_reg,track_data_v_r_7_sv2v_reg,track_data_v_r_6_sv2v_reg,
  track_data_v_r_5_sv2v_reg,track_data_v_r_4_sv2v_reg,track_data_v_r_3_sv2v_reg,
  track_data_v_r_2_sv2v_reg,track_data_v_r_1_sv2v_reg,track_data_v_r_0_sv2v_reg,
  mask_v_r_15_sv2v_reg,mask_v_r_14_sv2v_reg,mask_v_r_13_sv2v_reg,mask_v_r_12_sv2v_reg,
  mask_v_r_11_sv2v_reg,mask_v_r_10_sv2v_reg,mask_v_r_9_sv2v_reg,mask_v_r_8_sv2v_reg,
  mask_v_r_7_sv2v_reg,mask_v_r_6_sv2v_reg,mask_v_r_5_sv2v_reg,mask_v_r_4_sv2v_reg,
  mask_v_r_3_sv2v_reg,mask_v_r_2_sv2v_reg,mask_v_r_1_sv2v_reg,mask_v_r_0_sv2v_reg,
  decode_v_r_20_sv2v_reg,decode_v_r_19_sv2v_reg,decode_v_r_18_sv2v_reg,
  decode_v_r_17_sv2v_reg,decode_v_r_16_sv2v_reg,decode_v_r_15_sv2v_reg,decode_v_r_14_sv2v_reg,
  decode_v_r_13_sv2v_reg,decode_v_r_12_sv2v_reg,decode_v_r_11_sv2v_reg,
  decode_v_r_10_sv2v_reg,decode_v_r_9_sv2v_reg,decode_v_r_8_sv2v_reg,decode_v_r_7_sv2v_reg,
  decode_v_r_6_sv2v_reg,decode_v_r_5_sv2v_reg,decode_v_r_4_sv2v_reg,decode_v_r_3_sv2v_reg,
  decode_v_r_2_sv2v_reg,decode_v_r_1_sv2v_reg,decode_v_r_0_sv2v_reg,
  addr_v_r_32_sv2v_reg,addr_v_r_31_sv2v_reg,addr_v_r_30_sv2v_reg,addr_v_r_29_sv2v_reg,
  addr_v_r_28_sv2v_reg,addr_v_r_27_sv2v_reg,addr_v_r_26_sv2v_reg,addr_v_r_25_sv2v_reg,
  addr_v_r_24_sv2v_reg,addr_v_r_23_sv2v_reg,addr_v_r_22_sv2v_reg,addr_v_r_21_sv2v_reg,
  addr_v_r_20_sv2v_reg,addr_v_r_19_sv2v_reg,addr_v_r_18_sv2v_reg,addr_v_r_17_sv2v_reg,
  addr_v_r_16_sv2v_reg,addr_v_r_15_sv2v_reg,addr_v_r_14_sv2v_reg,
  addr_v_r_13_sv2v_reg,addr_v_r_12_sv2v_reg,addr_v_r_11_sv2v_reg,addr_v_r_10_sv2v_reg,
  addr_v_r_9_sv2v_reg,addr_v_r_8_sv2v_reg,addr_v_r_7_sv2v_reg,addr_v_r_6_sv2v_reg,
  addr_v_r_5_sv2v_reg,addr_v_r_4_sv2v_reg,addr_v_r_3_sv2v_reg,addr_v_r_2_sv2v_reg,
  addr_v_r_1_sv2v_reg,addr_v_r_0_sv2v_reg,data_v_r_127_sv2v_reg,data_v_r_126_sv2v_reg,
  data_v_r_125_sv2v_reg,data_v_r_124_sv2v_reg,data_v_r_123_sv2v_reg,data_v_r_122_sv2v_reg,
  data_v_r_121_sv2v_reg,data_v_r_120_sv2v_reg,data_v_r_119_sv2v_reg,
  data_v_r_118_sv2v_reg,data_v_r_117_sv2v_reg,data_v_r_116_sv2v_reg,data_v_r_115_sv2v_reg,
  data_v_r_114_sv2v_reg,data_v_r_113_sv2v_reg,data_v_r_112_sv2v_reg,
  data_v_r_111_sv2v_reg,data_v_r_110_sv2v_reg,data_v_r_109_sv2v_reg,data_v_r_108_sv2v_reg,
  data_v_r_107_sv2v_reg,data_v_r_106_sv2v_reg,data_v_r_105_sv2v_reg,data_v_r_104_sv2v_reg,
  data_v_r_103_sv2v_reg,data_v_r_102_sv2v_reg,data_v_r_101_sv2v_reg,
  data_v_r_100_sv2v_reg,data_v_r_99_sv2v_reg,data_v_r_98_sv2v_reg,data_v_r_97_sv2v_reg,
  data_v_r_96_sv2v_reg,data_v_r_95_sv2v_reg,data_v_r_94_sv2v_reg,data_v_r_93_sv2v_reg,
  data_v_r_92_sv2v_reg,data_v_r_91_sv2v_reg,data_v_r_90_sv2v_reg,data_v_r_89_sv2v_reg,
  data_v_r_88_sv2v_reg,data_v_r_87_sv2v_reg,data_v_r_86_sv2v_reg,data_v_r_85_sv2v_reg,
  data_v_r_84_sv2v_reg,data_v_r_83_sv2v_reg,data_v_r_82_sv2v_reg,
  data_v_r_81_sv2v_reg,data_v_r_80_sv2v_reg,data_v_r_79_sv2v_reg,data_v_r_78_sv2v_reg,
  data_v_r_77_sv2v_reg,data_v_r_76_sv2v_reg,data_v_r_75_sv2v_reg,data_v_r_74_sv2v_reg,
  data_v_r_73_sv2v_reg,data_v_r_72_sv2v_reg,data_v_r_71_sv2v_reg,data_v_r_70_sv2v_reg,
  data_v_r_69_sv2v_reg,data_v_r_68_sv2v_reg,data_v_r_67_sv2v_reg,data_v_r_66_sv2v_reg,
  data_v_r_65_sv2v_reg,data_v_r_64_sv2v_reg,data_v_r_63_sv2v_reg,
  data_v_r_62_sv2v_reg,data_v_r_61_sv2v_reg,data_v_r_60_sv2v_reg,data_v_r_59_sv2v_reg,
  data_v_r_58_sv2v_reg,data_v_r_57_sv2v_reg,data_v_r_56_sv2v_reg,data_v_r_55_sv2v_reg,
  data_v_r_54_sv2v_reg,data_v_r_53_sv2v_reg,data_v_r_52_sv2v_reg,data_v_r_51_sv2v_reg,
  data_v_r_50_sv2v_reg,data_v_r_49_sv2v_reg,data_v_r_48_sv2v_reg,data_v_r_47_sv2v_reg,
  data_v_r_46_sv2v_reg,data_v_r_45_sv2v_reg,data_v_r_44_sv2v_reg,data_v_r_43_sv2v_reg,
  data_v_r_42_sv2v_reg,data_v_r_41_sv2v_reg,data_v_r_40_sv2v_reg,
  data_v_r_39_sv2v_reg,data_v_r_38_sv2v_reg,data_v_r_37_sv2v_reg,data_v_r_36_sv2v_reg,
  data_v_r_35_sv2v_reg,data_v_r_34_sv2v_reg,data_v_r_33_sv2v_reg,data_v_r_32_sv2v_reg,
  data_v_r_31_sv2v_reg,data_v_r_30_sv2v_reg,data_v_r_29_sv2v_reg,data_v_r_28_sv2v_reg,
  data_v_r_27_sv2v_reg,data_v_r_26_sv2v_reg,data_v_r_25_sv2v_reg,data_v_r_24_sv2v_reg,
  data_v_r_23_sv2v_reg,data_v_r_22_sv2v_reg,data_v_r_21_sv2v_reg,
  data_v_r_20_sv2v_reg,data_v_r_19_sv2v_reg,data_v_r_18_sv2v_reg,data_v_r_17_sv2v_reg,
  data_v_r_16_sv2v_reg,data_v_r_15_sv2v_reg,data_v_r_14_sv2v_reg,data_v_r_13_sv2v_reg,
  data_v_r_12_sv2v_reg,data_v_r_11_sv2v_reg,data_v_r_10_sv2v_reg,data_v_r_9_sv2v_reg,
  data_v_r_8_sv2v_reg,data_v_r_7_sv2v_reg,data_v_r_6_sv2v_reg,data_v_r_5_sv2v_reg,
  data_v_r_4_sv2v_reg,data_v_r_3_sv2v_reg,data_v_r_2_sv2v_reg,data_v_r_1_sv2v_reg,
  data_v_r_0_sv2v_reg,valid_v_r_7_sv2v_reg,valid_v_r_6_sv2v_reg,valid_v_r_5_sv2v_reg,
  valid_v_r_4_sv2v_reg,valid_v_r_3_sv2v_reg,valid_v_r_2_sv2v_reg,valid_v_r_1_sv2v_reg,
  valid_v_r_0_sv2v_reg,lock_v_r_7_sv2v_reg,lock_v_r_6_sv2v_reg,
  lock_v_r_5_sv2v_reg,lock_v_r_4_sv2v_reg,lock_v_r_3_sv2v_reg,lock_v_r_2_sv2v_reg,
  lock_v_r_1_sv2v_reg,lock_v_r_0_sv2v_reg,tag_v_r_159_sv2v_reg,tag_v_r_158_sv2v_reg,
  tag_v_r_157_sv2v_reg,tag_v_r_156_sv2v_reg,tag_v_r_155_sv2v_reg,tag_v_r_154_sv2v_reg,
  tag_v_r_153_sv2v_reg,tag_v_r_152_sv2v_reg,tag_v_r_151_sv2v_reg,tag_v_r_150_sv2v_reg,
  tag_v_r_149_sv2v_reg,tag_v_r_148_sv2v_reg,tag_v_r_147_sv2v_reg,tag_v_r_146_sv2v_reg,
  tag_v_r_145_sv2v_reg,tag_v_r_144_sv2v_reg,tag_v_r_143_sv2v_reg,tag_v_r_142_sv2v_reg,
  tag_v_r_141_sv2v_reg,tag_v_r_140_sv2v_reg,tag_v_r_139_sv2v_reg,
  tag_v_r_138_sv2v_reg,tag_v_r_137_sv2v_reg,tag_v_r_136_sv2v_reg,tag_v_r_135_sv2v_reg,
  tag_v_r_134_sv2v_reg,tag_v_r_133_sv2v_reg,tag_v_r_132_sv2v_reg,tag_v_r_131_sv2v_reg,
  tag_v_r_130_sv2v_reg,tag_v_r_129_sv2v_reg,tag_v_r_128_sv2v_reg,tag_v_r_127_sv2v_reg,
  tag_v_r_126_sv2v_reg,tag_v_r_125_sv2v_reg,tag_v_r_124_sv2v_reg,tag_v_r_123_sv2v_reg,
  tag_v_r_122_sv2v_reg,tag_v_r_121_sv2v_reg,tag_v_r_120_sv2v_reg,
  tag_v_r_119_sv2v_reg,tag_v_r_118_sv2v_reg,tag_v_r_117_sv2v_reg,tag_v_r_116_sv2v_reg,
  tag_v_r_115_sv2v_reg,tag_v_r_114_sv2v_reg,tag_v_r_113_sv2v_reg,tag_v_r_112_sv2v_reg,
  tag_v_r_111_sv2v_reg,tag_v_r_110_sv2v_reg,tag_v_r_109_sv2v_reg,tag_v_r_108_sv2v_reg,
  tag_v_r_107_sv2v_reg,tag_v_r_106_sv2v_reg,tag_v_r_105_sv2v_reg,tag_v_r_104_sv2v_reg,
  tag_v_r_103_sv2v_reg,tag_v_r_102_sv2v_reg,tag_v_r_101_sv2v_reg,
  tag_v_r_100_sv2v_reg,tag_v_r_99_sv2v_reg,tag_v_r_98_sv2v_reg,tag_v_r_97_sv2v_reg,
  tag_v_r_96_sv2v_reg,tag_v_r_95_sv2v_reg,tag_v_r_94_sv2v_reg,tag_v_r_93_sv2v_reg,
  tag_v_r_92_sv2v_reg,tag_v_r_91_sv2v_reg,tag_v_r_90_sv2v_reg,tag_v_r_89_sv2v_reg,
  tag_v_r_88_sv2v_reg,tag_v_r_87_sv2v_reg,tag_v_r_86_sv2v_reg,tag_v_r_85_sv2v_reg,
  tag_v_r_84_sv2v_reg,tag_v_r_83_sv2v_reg,tag_v_r_82_sv2v_reg,tag_v_r_81_sv2v_reg,
  tag_v_r_80_sv2v_reg,tag_v_r_79_sv2v_reg,tag_v_r_78_sv2v_reg,tag_v_r_77_sv2v_reg,
  tag_v_r_76_sv2v_reg,tag_v_r_75_sv2v_reg,tag_v_r_74_sv2v_reg,tag_v_r_73_sv2v_reg,
  tag_v_r_72_sv2v_reg,tag_v_r_71_sv2v_reg,tag_v_r_70_sv2v_reg,tag_v_r_69_sv2v_reg,
  tag_v_r_68_sv2v_reg,tag_v_r_67_sv2v_reg,tag_v_r_66_sv2v_reg,tag_v_r_65_sv2v_reg,
  tag_v_r_64_sv2v_reg,tag_v_r_63_sv2v_reg,tag_v_r_62_sv2v_reg,tag_v_r_61_sv2v_reg,
  tag_v_r_60_sv2v_reg,tag_v_r_59_sv2v_reg,tag_v_r_58_sv2v_reg,tag_v_r_57_sv2v_reg,
  tag_v_r_56_sv2v_reg,tag_v_r_55_sv2v_reg,tag_v_r_54_sv2v_reg,tag_v_r_53_sv2v_reg,
  tag_v_r_52_sv2v_reg,tag_v_r_51_sv2v_reg,tag_v_r_50_sv2v_reg,tag_v_r_49_sv2v_reg,
  tag_v_r_48_sv2v_reg,tag_v_r_47_sv2v_reg,tag_v_r_46_sv2v_reg,tag_v_r_45_sv2v_reg,
  tag_v_r_44_sv2v_reg,tag_v_r_43_sv2v_reg,tag_v_r_42_sv2v_reg,tag_v_r_41_sv2v_reg,
  tag_v_r_40_sv2v_reg,tag_v_r_39_sv2v_reg,tag_v_r_38_sv2v_reg,tag_v_r_37_sv2v_reg,
  tag_v_r_36_sv2v_reg,tag_v_r_35_sv2v_reg,tag_v_r_34_sv2v_reg,tag_v_r_33_sv2v_reg,
  tag_v_r_32_sv2v_reg,tag_v_r_31_sv2v_reg,tag_v_r_30_sv2v_reg,tag_v_r_29_sv2v_reg,
  tag_v_r_28_sv2v_reg,tag_v_r_27_sv2v_reg,tag_v_r_26_sv2v_reg,tag_v_r_25_sv2v_reg,
  tag_v_r_24_sv2v_reg,tag_v_r_23_sv2v_reg,tag_v_r_22_sv2v_reg,tag_v_r_21_sv2v_reg,
  tag_v_r_20_sv2v_reg,tag_v_r_19_sv2v_reg,tag_v_r_18_sv2v_reg,tag_v_r_17_sv2v_reg,
  tag_v_r_16_sv2v_reg,tag_v_r_15_sv2v_reg,tag_v_r_14_sv2v_reg,tag_v_r_13_sv2v_reg,
  tag_v_r_12_sv2v_reg,tag_v_r_11_sv2v_reg,tag_v_r_10_sv2v_reg,tag_v_r_9_sv2v_reg,tag_v_r_8_sv2v_reg,
  tag_v_r_7_sv2v_reg,tag_v_r_6_sv2v_reg,tag_v_r_5_sv2v_reg,tag_v_r_4_sv2v_reg,
  tag_v_r_3_sv2v_reg,tag_v_r_2_sv2v_reg,tag_v_r_1_sv2v_reg,tag_v_r_0_sv2v_reg;
  assign data_tl_r[127] = data_tl_r_127_sv2v_reg;
  assign data_tl_r[126] = data_tl_r_126_sv2v_reg;
  assign data_tl_r[125] = data_tl_r_125_sv2v_reg;
  assign data_tl_r[124] = data_tl_r_124_sv2v_reg;
  assign data_tl_r[123] = data_tl_r_123_sv2v_reg;
  assign data_tl_r[122] = data_tl_r_122_sv2v_reg;
  assign data_tl_r[121] = data_tl_r_121_sv2v_reg;
  assign data_tl_r[120] = data_tl_r_120_sv2v_reg;
  assign data_tl_r[119] = data_tl_r_119_sv2v_reg;
  assign data_tl_r[118] = data_tl_r_118_sv2v_reg;
  assign data_tl_r[117] = data_tl_r_117_sv2v_reg;
  assign data_tl_r[116] = data_tl_r_116_sv2v_reg;
  assign data_tl_r[115] = data_tl_r_115_sv2v_reg;
  assign data_tl_r[114] = data_tl_r_114_sv2v_reg;
  assign data_tl_r[113] = data_tl_r_113_sv2v_reg;
  assign data_tl_r[112] = data_tl_r_112_sv2v_reg;
  assign data_tl_r[111] = data_tl_r_111_sv2v_reg;
  assign data_tl_r[110] = data_tl_r_110_sv2v_reg;
  assign data_tl_r[109] = data_tl_r_109_sv2v_reg;
  assign data_tl_r[108] = data_tl_r_108_sv2v_reg;
  assign data_tl_r[107] = data_tl_r_107_sv2v_reg;
  assign data_tl_r[106] = data_tl_r_106_sv2v_reg;
  assign data_tl_r[105] = data_tl_r_105_sv2v_reg;
  assign data_tl_r[104] = data_tl_r_104_sv2v_reg;
  assign data_tl_r[103] = data_tl_r_103_sv2v_reg;
  assign data_tl_r[102] = data_tl_r_102_sv2v_reg;
  assign data_tl_r[101] = data_tl_r_101_sv2v_reg;
  assign data_tl_r[100] = data_tl_r_100_sv2v_reg;
  assign data_tl_r[99] = data_tl_r_99_sv2v_reg;
  assign data_tl_r[98] = data_tl_r_98_sv2v_reg;
  assign data_tl_r[97] = data_tl_r_97_sv2v_reg;
  assign data_tl_r[96] = data_tl_r_96_sv2v_reg;
  assign data_tl_r[95] = data_tl_r_95_sv2v_reg;
  assign data_tl_r[94] = data_tl_r_94_sv2v_reg;
  assign data_tl_r[93] = data_tl_r_93_sv2v_reg;
  assign data_tl_r[92] = data_tl_r_92_sv2v_reg;
  assign data_tl_r[91] = data_tl_r_91_sv2v_reg;
  assign data_tl_r[90] = data_tl_r_90_sv2v_reg;
  assign data_tl_r[89] = data_tl_r_89_sv2v_reg;
  assign data_tl_r[88] = data_tl_r_88_sv2v_reg;
  assign data_tl_r[87] = data_tl_r_87_sv2v_reg;
  assign data_tl_r[86] = data_tl_r_86_sv2v_reg;
  assign data_tl_r[85] = data_tl_r_85_sv2v_reg;
  assign data_tl_r[84] = data_tl_r_84_sv2v_reg;
  assign data_tl_r[83] = data_tl_r_83_sv2v_reg;
  assign data_tl_r[82] = data_tl_r_82_sv2v_reg;
  assign data_tl_r[81] = data_tl_r_81_sv2v_reg;
  assign data_tl_r[80] = data_tl_r_80_sv2v_reg;
  assign data_tl_r[79] = data_tl_r_79_sv2v_reg;
  assign data_tl_r[78] = data_tl_r_78_sv2v_reg;
  assign data_tl_r[77] = data_tl_r_77_sv2v_reg;
  assign data_tl_r[76] = data_tl_r_76_sv2v_reg;
  assign data_tl_r[75] = data_tl_r_75_sv2v_reg;
  assign data_tl_r[74] = data_tl_r_74_sv2v_reg;
  assign data_tl_r[73] = data_tl_r_73_sv2v_reg;
  assign data_tl_r[72] = data_tl_r_72_sv2v_reg;
  assign data_tl_r[71] = data_tl_r_71_sv2v_reg;
  assign data_tl_r[70] = data_tl_r_70_sv2v_reg;
  assign data_tl_r[69] = data_tl_r_69_sv2v_reg;
  assign data_tl_r[68] = data_tl_r_68_sv2v_reg;
  assign data_tl_r[67] = data_tl_r_67_sv2v_reg;
  assign data_tl_r[66] = data_tl_r_66_sv2v_reg;
  assign data_tl_r[65] = data_tl_r_65_sv2v_reg;
  assign data_tl_r[64] = data_tl_r_64_sv2v_reg;
  assign data_tl_r[63] = data_tl_r_63_sv2v_reg;
  assign data_tl_r[62] = data_tl_r_62_sv2v_reg;
  assign data_tl_r[61] = data_tl_r_61_sv2v_reg;
  assign data_tl_r[60] = data_tl_r_60_sv2v_reg;
  assign data_tl_r[59] = data_tl_r_59_sv2v_reg;
  assign data_tl_r[58] = data_tl_r_58_sv2v_reg;
  assign data_tl_r[57] = data_tl_r_57_sv2v_reg;
  assign data_tl_r[56] = data_tl_r_56_sv2v_reg;
  assign data_tl_r[55] = data_tl_r_55_sv2v_reg;
  assign data_tl_r[54] = data_tl_r_54_sv2v_reg;
  assign data_tl_r[53] = data_tl_r_53_sv2v_reg;
  assign data_tl_r[52] = data_tl_r_52_sv2v_reg;
  assign data_tl_r[51] = data_tl_r_51_sv2v_reg;
  assign data_tl_r[50] = data_tl_r_50_sv2v_reg;
  assign data_tl_r[49] = data_tl_r_49_sv2v_reg;
  assign data_tl_r[48] = data_tl_r_48_sv2v_reg;
  assign data_tl_r[47] = data_tl_r_47_sv2v_reg;
  assign data_tl_r[46] = data_tl_r_46_sv2v_reg;
  assign data_tl_r[45] = data_tl_r_45_sv2v_reg;
  assign data_tl_r[44] = data_tl_r_44_sv2v_reg;
  assign data_tl_r[43] = data_tl_r_43_sv2v_reg;
  assign data_tl_r[42] = data_tl_r_42_sv2v_reg;
  assign data_tl_r[41] = data_tl_r_41_sv2v_reg;
  assign data_tl_r[40] = data_tl_r_40_sv2v_reg;
  assign data_tl_r[39] = data_tl_r_39_sv2v_reg;
  assign data_tl_r[38] = data_tl_r_38_sv2v_reg;
  assign data_tl_r[37] = data_tl_r_37_sv2v_reg;
  assign data_tl_r[36] = data_tl_r_36_sv2v_reg;
  assign data_tl_r[35] = data_tl_r_35_sv2v_reg;
  assign data_tl_r[34] = data_tl_r_34_sv2v_reg;
  assign data_tl_r[33] = data_tl_r_33_sv2v_reg;
  assign data_tl_r[32] = data_tl_r_32_sv2v_reg;
  assign data_tl_r[31] = data_tl_r_31_sv2v_reg;
  assign data_tl_r[30] = data_tl_r_30_sv2v_reg;
  assign data_tl_r[29] = data_tl_r_29_sv2v_reg;
  assign data_tl_r[28] = data_tl_r_28_sv2v_reg;
  assign data_tl_r[27] = data_tl_r_27_sv2v_reg;
  assign data_tl_r[26] = data_tl_r_26_sv2v_reg;
  assign data_tl_r[25] = data_tl_r_25_sv2v_reg;
  assign data_tl_r[24] = data_tl_r_24_sv2v_reg;
  assign data_tl_r[23] = data_tl_r_23_sv2v_reg;
  assign data_tl_r[22] = data_tl_r_22_sv2v_reg;
  assign data_tl_r[21] = data_tl_r_21_sv2v_reg;
  assign data_tl_r[20] = data_tl_r_20_sv2v_reg;
  assign data_tl_r[19] = data_tl_r_19_sv2v_reg;
  assign data_tl_r[18] = data_tl_r_18_sv2v_reg;
  assign data_tl_r[17] = data_tl_r_17_sv2v_reg;
  assign data_tl_r[16] = data_tl_r_16_sv2v_reg;
  assign data_tl_r[15] = data_tl_r_15_sv2v_reg;
  assign data_tl_r[14] = data_tl_r_14_sv2v_reg;
  assign data_tl_r[13] = data_tl_r_13_sv2v_reg;
  assign data_tl_r[12] = data_tl_r_12_sv2v_reg;
  assign data_tl_r[11] = data_tl_r_11_sv2v_reg;
  assign data_tl_r[10] = data_tl_r_10_sv2v_reg;
  assign data_tl_r[9] = data_tl_r_9_sv2v_reg;
  assign data_tl_r[8] = data_tl_r_8_sv2v_reg;
  assign data_tl_r[7] = data_tl_r_7_sv2v_reg;
  assign data_tl_r[6] = data_tl_r_6_sv2v_reg;
  assign data_tl_r[5] = data_tl_r_5_sv2v_reg;
  assign data_tl_r[4] = data_tl_r_4_sv2v_reg;
  assign data_tl_r[3] = data_tl_r_3_sv2v_reg;
  assign data_tl_r[2] = data_tl_r_2_sv2v_reg;
  assign data_tl_r[1] = data_tl_r_1_sv2v_reg;
  assign data_tl_r[0] = data_tl_r_0_sv2v_reg;
  assign v_tl_r = v_tl_r_sv2v_reg;
  assign decode_tl_r[20] = decode_tl_r_20_sv2v_reg;
  assign decode_tl_r[19] = decode_tl_r_19_sv2v_reg;
  assign decode_tl_r[18] = decode_tl_r_18_sv2v_reg;
  assign decode_tl_r[17] = decode_tl_r_17_sv2v_reg;
  assign decode_tl_r[16] = decode_tl_r_16_sv2v_reg;
  assign decode_tl_r[15] = decode_tl_r_15_sv2v_reg;
  assign decode_tl_r[14] = decode_tl_r_14_sv2v_reg;
  assign decode_tl_r[13] = decode_tl_r_13_sv2v_reg;
  assign decode_tl_r[12] = decode_tl_r_12_sv2v_reg;
  assign decode_tl_r[11] = decode_tl_r_11_sv2v_reg;
  assign decode_tl_r[10] = decode_tl_r_10_sv2v_reg;
  assign decode_tl_r[9] = decode_tl_r_9_sv2v_reg;
  assign decode_tl_r[8] = decode_tl_r_8_sv2v_reg;
  assign decode_tl_r[7] = decode_tl_r_7_sv2v_reg;
  assign decode_tl_r[6] = decode_tl_r_6_sv2v_reg;
  assign decode_tl_r[5] = decode_tl_r_5_sv2v_reg;
  assign decode_tl_r[4] = decode_tl_r_4_sv2v_reg;
  assign decode_tl_r[3] = decode_tl_r_3_sv2v_reg;
  assign decode_tl_r[2] = decode_tl_r_2_sv2v_reg;
  assign decode_tl_r[1] = decode_tl_r_1_sv2v_reg;
  assign decode_tl_r[0] = decode_tl_r_0_sv2v_reg;
  assign mask_tl_r[15] = mask_tl_r_15_sv2v_reg;
  assign mask_tl_r[14] = mask_tl_r_14_sv2v_reg;
  assign mask_tl_r[13] = mask_tl_r_13_sv2v_reg;
  assign mask_tl_r[12] = mask_tl_r_12_sv2v_reg;
  assign mask_tl_r[11] = mask_tl_r_11_sv2v_reg;
  assign mask_tl_r[10] = mask_tl_r_10_sv2v_reg;
  assign mask_tl_r[9] = mask_tl_r_9_sv2v_reg;
  assign mask_tl_r[8] = mask_tl_r_8_sv2v_reg;
  assign mask_tl_r[7] = mask_tl_r_7_sv2v_reg;
  assign mask_tl_r[6] = mask_tl_r_6_sv2v_reg;
  assign mask_tl_r[5] = mask_tl_r_5_sv2v_reg;
  assign mask_tl_r[4] = mask_tl_r_4_sv2v_reg;
  assign mask_tl_r[3] = mask_tl_r_3_sv2v_reg;
  assign mask_tl_r[2] = mask_tl_r_2_sv2v_reg;
  assign mask_tl_r[1] = mask_tl_r_1_sv2v_reg;
  assign mask_tl_r[0] = mask_tl_r_0_sv2v_reg;
  assign addr_tl_r[32] = addr_tl_r_32_sv2v_reg;
  assign addr_tl_r[31] = addr_tl_r_31_sv2v_reg;
  assign addr_tl_r[30] = addr_tl_r_30_sv2v_reg;
  assign addr_tl_r[29] = addr_tl_r_29_sv2v_reg;
  assign addr_tl_r[28] = addr_tl_r_28_sv2v_reg;
  assign addr_tl_r[27] = addr_tl_r_27_sv2v_reg;
  assign addr_tl_r[26] = addr_tl_r_26_sv2v_reg;
  assign addr_tl_r[25] = addr_tl_r_25_sv2v_reg;
  assign addr_tl_r[24] = addr_tl_r_24_sv2v_reg;
  assign addr_tl_r[23] = addr_tl_r_23_sv2v_reg;
  assign addr_tl_r[22] = addr_tl_r_22_sv2v_reg;
  assign addr_tl_r[21] = addr_tl_r_21_sv2v_reg;
  assign addr_tl_r[20] = addr_tl_r_20_sv2v_reg;
  assign addr_tl_r[19] = addr_tl_r_19_sv2v_reg;
  assign addr_tl_r[18] = addr_tl_r_18_sv2v_reg;
  assign addr_tl_r[17] = addr_tl_r_17_sv2v_reg;
  assign addr_tl_r[16] = addr_tl_r_16_sv2v_reg;
  assign addr_tl_r[15] = addr_tl_r_15_sv2v_reg;
  assign addr_tl_r[14] = addr_tl_r_14_sv2v_reg;
  assign addr_tl_r[13] = addr_tl_r_13_sv2v_reg;
  assign addr_tl_r[12] = addr_tl_r_12_sv2v_reg;
  assign addr_tl_r[11] = addr_tl_r_11_sv2v_reg;
  assign addr_tl_r[10] = addr_tl_r_10_sv2v_reg;
  assign addr_tl_r[9] = addr_tl_r_9_sv2v_reg;
  assign addr_tl_r[8] = addr_tl_r_8_sv2v_reg;
  assign addr_tl_r[7] = addr_tl_r_7_sv2v_reg;
  assign addr_tl_r[6] = addr_tl_r_6_sv2v_reg;
  assign addr_tl_r[5] = addr_tl_r_5_sv2v_reg;
  assign addr_tl_r[4] = addr_tl_r_4_sv2v_reg;
  assign addr_tl_r[3] = addr_tl_r_3_sv2v_reg;
  assign addr_tl_r[2] = addr_tl_r_2_sv2v_reg;
  assign addr_tl_r[1] = addr_tl_r_1_sv2v_reg;
  assign addr_tl_r[0] = addr_tl_r_0_sv2v_reg;
  assign ld_data_v_r[1023] = ld_data_v_r_1023_sv2v_reg;
  assign ld_data_v_r[1022] = ld_data_v_r_1022_sv2v_reg;
  assign ld_data_v_r[1021] = ld_data_v_r_1021_sv2v_reg;
  assign ld_data_v_r[1020] = ld_data_v_r_1020_sv2v_reg;
  assign ld_data_v_r[1019] = ld_data_v_r_1019_sv2v_reg;
  assign ld_data_v_r[1018] = ld_data_v_r_1018_sv2v_reg;
  assign ld_data_v_r[1017] = ld_data_v_r_1017_sv2v_reg;
  assign ld_data_v_r[1016] = ld_data_v_r_1016_sv2v_reg;
  assign ld_data_v_r[1015] = ld_data_v_r_1015_sv2v_reg;
  assign ld_data_v_r[1014] = ld_data_v_r_1014_sv2v_reg;
  assign ld_data_v_r[1013] = ld_data_v_r_1013_sv2v_reg;
  assign ld_data_v_r[1012] = ld_data_v_r_1012_sv2v_reg;
  assign ld_data_v_r[1011] = ld_data_v_r_1011_sv2v_reg;
  assign ld_data_v_r[1010] = ld_data_v_r_1010_sv2v_reg;
  assign ld_data_v_r[1009] = ld_data_v_r_1009_sv2v_reg;
  assign ld_data_v_r[1008] = ld_data_v_r_1008_sv2v_reg;
  assign ld_data_v_r[1007] = ld_data_v_r_1007_sv2v_reg;
  assign ld_data_v_r[1006] = ld_data_v_r_1006_sv2v_reg;
  assign ld_data_v_r[1005] = ld_data_v_r_1005_sv2v_reg;
  assign ld_data_v_r[1004] = ld_data_v_r_1004_sv2v_reg;
  assign ld_data_v_r[1003] = ld_data_v_r_1003_sv2v_reg;
  assign ld_data_v_r[1002] = ld_data_v_r_1002_sv2v_reg;
  assign ld_data_v_r[1001] = ld_data_v_r_1001_sv2v_reg;
  assign ld_data_v_r[1000] = ld_data_v_r_1000_sv2v_reg;
  assign ld_data_v_r[999] = ld_data_v_r_999_sv2v_reg;
  assign ld_data_v_r[998] = ld_data_v_r_998_sv2v_reg;
  assign ld_data_v_r[997] = ld_data_v_r_997_sv2v_reg;
  assign ld_data_v_r[996] = ld_data_v_r_996_sv2v_reg;
  assign ld_data_v_r[995] = ld_data_v_r_995_sv2v_reg;
  assign ld_data_v_r[994] = ld_data_v_r_994_sv2v_reg;
  assign ld_data_v_r[993] = ld_data_v_r_993_sv2v_reg;
  assign ld_data_v_r[992] = ld_data_v_r_992_sv2v_reg;
  assign ld_data_v_r[991] = ld_data_v_r_991_sv2v_reg;
  assign ld_data_v_r[990] = ld_data_v_r_990_sv2v_reg;
  assign ld_data_v_r[989] = ld_data_v_r_989_sv2v_reg;
  assign ld_data_v_r[988] = ld_data_v_r_988_sv2v_reg;
  assign ld_data_v_r[987] = ld_data_v_r_987_sv2v_reg;
  assign ld_data_v_r[986] = ld_data_v_r_986_sv2v_reg;
  assign ld_data_v_r[985] = ld_data_v_r_985_sv2v_reg;
  assign ld_data_v_r[984] = ld_data_v_r_984_sv2v_reg;
  assign ld_data_v_r[983] = ld_data_v_r_983_sv2v_reg;
  assign ld_data_v_r[982] = ld_data_v_r_982_sv2v_reg;
  assign ld_data_v_r[981] = ld_data_v_r_981_sv2v_reg;
  assign ld_data_v_r[980] = ld_data_v_r_980_sv2v_reg;
  assign ld_data_v_r[979] = ld_data_v_r_979_sv2v_reg;
  assign ld_data_v_r[978] = ld_data_v_r_978_sv2v_reg;
  assign ld_data_v_r[977] = ld_data_v_r_977_sv2v_reg;
  assign ld_data_v_r[976] = ld_data_v_r_976_sv2v_reg;
  assign ld_data_v_r[975] = ld_data_v_r_975_sv2v_reg;
  assign ld_data_v_r[974] = ld_data_v_r_974_sv2v_reg;
  assign ld_data_v_r[973] = ld_data_v_r_973_sv2v_reg;
  assign ld_data_v_r[972] = ld_data_v_r_972_sv2v_reg;
  assign ld_data_v_r[971] = ld_data_v_r_971_sv2v_reg;
  assign ld_data_v_r[970] = ld_data_v_r_970_sv2v_reg;
  assign ld_data_v_r[969] = ld_data_v_r_969_sv2v_reg;
  assign ld_data_v_r[968] = ld_data_v_r_968_sv2v_reg;
  assign ld_data_v_r[967] = ld_data_v_r_967_sv2v_reg;
  assign ld_data_v_r[966] = ld_data_v_r_966_sv2v_reg;
  assign ld_data_v_r[965] = ld_data_v_r_965_sv2v_reg;
  assign ld_data_v_r[964] = ld_data_v_r_964_sv2v_reg;
  assign ld_data_v_r[963] = ld_data_v_r_963_sv2v_reg;
  assign ld_data_v_r[962] = ld_data_v_r_962_sv2v_reg;
  assign ld_data_v_r[961] = ld_data_v_r_961_sv2v_reg;
  assign ld_data_v_r[960] = ld_data_v_r_960_sv2v_reg;
  assign ld_data_v_r[959] = ld_data_v_r_959_sv2v_reg;
  assign ld_data_v_r[958] = ld_data_v_r_958_sv2v_reg;
  assign ld_data_v_r[957] = ld_data_v_r_957_sv2v_reg;
  assign ld_data_v_r[956] = ld_data_v_r_956_sv2v_reg;
  assign ld_data_v_r[955] = ld_data_v_r_955_sv2v_reg;
  assign ld_data_v_r[954] = ld_data_v_r_954_sv2v_reg;
  assign ld_data_v_r[953] = ld_data_v_r_953_sv2v_reg;
  assign ld_data_v_r[952] = ld_data_v_r_952_sv2v_reg;
  assign ld_data_v_r[951] = ld_data_v_r_951_sv2v_reg;
  assign ld_data_v_r[950] = ld_data_v_r_950_sv2v_reg;
  assign ld_data_v_r[949] = ld_data_v_r_949_sv2v_reg;
  assign ld_data_v_r[948] = ld_data_v_r_948_sv2v_reg;
  assign ld_data_v_r[947] = ld_data_v_r_947_sv2v_reg;
  assign ld_data_v_r[946] = ld_data_v_r_946_sv2v_reg;
  assign ld_data_v_r[945] = ld_data_v_r_945_sv2v_reg;
  assign ld_data_v_r[944] = ld_data_v_r_944_sv2v_reg;
  assign ld_data_v_r[943] = ld_data_v_r_943_sv2v_reg;
  assign ld_data_v_r[942] = ld_data_v_r_942_sv2v_reg;
  assign ld_data_v_r[941] = ld_data_v_r_941_sv2v_reg;
  assign ld_data_v_r[940] = ld_data_v_r_940_sv2v_reg;
  assign ld_data_v_r[939] = ld_data_v_r_939_sv2v_reg;
  assign ld_data_v_r[938] = ld_data_v_r_938_sv2v_reg;
  assign ld_data_v_r[937] = ld_data_v_r_937_sv2v_reg;
  assign ld_data_v_r[936] = ld_data_v_r_936_sv2v_reg;
  assign ld_data_v_r[935] = ld_data_v_r_935_sv2v_reg;
  assign ld_data_v_r[934] = ld_data_v_r_934_sv2v_reg;
  assign ld_data_v_r[933] = ld_data_v_r_933_sv2v_reg;
  assign ld_data_v_r[932] = ld_data_v_r_932_sv2v_reg;
  assign ld_data_v_r[931] = ld_data_v_r_931_sv2v_reg;
  assign ld_data_v_r[930] = ld_data_v_r_930_sv2v_reg;
  assign ld_data_v_r[929] = ld_data_v_r_929_sv2v_reg;
  assign ld_data_v_r[928] = ld_data_v_r_928_sv2v_reg;
  assign ld_data_v_r[927] = ld_data_v_r_927_sv2v_reg;
  assign ld_data_v_r[926] = ld_data_v_r_926_sv2v_reg;
  assign ld_data_v_r[925] = ld_data_v_r_925_sv2v_reg;
  assign ld_data_v_r[924] = ld_data_v_r_924_sv2v_reg;
  assign ld_data_v_r[923] = ld_data_v_r_923_sv2v_reg;
  assign ld_data_v_r[922] = ld_data_v_r_922_sv2v_reg;
  assign ld_data_v_r[921] = ld_data_v_r_921_sv2v_reg;
  assign ld_data_v_r[920] = ld_data_v_r_920_sv2v_reg;
  assign ld_data_v_r[919] = ld_data_v_r_919_sv2v_reg;
  assign ld_data_v_r[918] = ld_data_v_r_918_sv2v_reg;
  assign ld_data_v_r[917] = ld_data_v_r_917_sv2v_reg;
  assign ld_data_v_r[916] = ld_data_v_r_916_sv2v_reg;
  assign ld_data_v_r[915] = ld_data_v_r_915_sv2v_reg;
  assign ld_data_v_r[914] = ld_data_v_r_914_sv2v_reg;
  assign ld_data_v_r[913] = ld_data_v_r_913_sv2v_reg;
  assign ld_data_v_r[912] = ld_data_v_r_912_sv2v_reg;
  assign ld_data_v_r[911] = ld_data_v_r_911_sv2v_reg;
  assign ld_data_v_r[910] = ld_data_v_r_910_sv2v_reg;
  assign ld_data_v_r[909] = ld_data_v_r_909_sv2v_reg;
  assign ld_data_v_r[908] = ld_data_v_r_908_sv2v_reg;
  assign ld_data_v_r[907] = ld_data_v_r_907_sv2v_reg;
  assign ld_data_v_r[906] = ld_data_v_r_906_sv2v_reg;
  assign ld_data_v_r[905] = ld_data_v_r_905_sv2v_reg;
  assign ld_data_v_r[904] = ld_data_v_r_904_sv2v_reg;
  assign ld_data_v_r[903] = ld_data_v_r_903_sv2v_reg;
  assign ld_data_v_r[902] = ld_data_v_r_902_sv2v_reg;
  assign ld_data_v_r[901] = ld_data_v_r_901_sv2v_reg;
  assign ld_data_v_r[900] = ld_data_v_r_900_sv2v_reg;
  assign ld_data_v_r[899] = ld_data_v_r_899_sv2v_reg;
  assign ld_data_v_r[898] = ld_data_v_r_898_sv2v_reg;
  assign ld_data_v_r[897] = ld_data_v_r_897_sv2v_reg;
  assign ld_data_v_r[896] = ld_data_v_r_896_sv2v_reg;
  assign ld_data_v_r[895] = ld_data_v_r_895_sv2v_reg;
  assign ld_data_v_r[894] = ld_data_v_r_894_sv2v_reg;
  assign ld_data_v_r[893] = ld_data_v_r_893_sv2v_reg;
  assign ld_data_v_r[892] = ld_data_v_r_892_sv2v_reg;
  assign ld_data_v_r[891] = ld_data_v_r_891_sv2v_reg;
  assign ld_data_v_r[890] = ld_data_v_r_890_sv2v_reg;
  assign ld_data_v_r[889] = ld_data_v_r_889_sv2v_reg;
  assign ld_data_v_r[888] = ld_data_v_r_888_sv2v_reg;
  assign ld_data_v_r[887] = ld_data_v_r_887_sv2v_reg;
  assign ld_data_v_r[886] = ld_data_v_r_886_sv2v_reg;
  assign ld_data_v_r[885] = ld_data_v_r_885_sv2v_reg;
  assign ld_data_v_r[884] = ld_data_v_r_884_sv2v_reg;
  assign ld_data_v_r[883] = ld_data_v_r_883_sv2v_reg;
  assign ld_data_v_r[882] = ld_data_v_r_882_sv2v_reg;
  assign ld_data_v_r[881] = ld_data_v_r_881_sv2v_reg;
  assign ld_data_v_r[880] = ld_data_v_r_880_sv2v_reg;
  assign ld_data_v_r[879] = ld_data_v_r_879_sv2v_reg;
  assign ld_data_v_r[878] = ld_data_v_r_878_sv2v_reg;
  assign ld_data_v_r[877] = ld_data_v_r_877_sv2v_reg;
  assign ld_data_v_r[876] = ld_data_v_r_876_sv2v_reg;
  assign ld_data_v_r[875] = ld_data_v_r_875_sv2v_reg;
  assign ld_data_v_r[874] = ld_data_v_r_874_sv2v_reg;
  assign ld_data_v_r[873] = ld_data_v_r_873_sv2v_reg;
  assign ld_data_v_r[872] = ld_data_v_r_872_sv2v_reg;
  assign ld_data_v_r[871] = ld_data_v_r_871_sv2v_reg;
  assign ld_data_v_r[870] = ld_data_v_r_870_sv2v_reg;
  assign ld_data_v_r[869] = ld_data_v_r_869_sv2v_reg;
  assign ld_data_v_r[868] = ld_data_v_r_868_sv2v_reg;
  assign ld_data_v_r[867] = ld_data_v_r_867_sv2v_reg;
  assign ld_data_v_r[866] = ld_data_v_r_866_sv2v_reg;
  assign ld_data_v_r[865] = ld_data_v_r_865_sv2v_reg;
  assign ld_data_v_r[864] = ld_data_v_r_864_sv2v_reg;
  assign ld_data_v_r[863] = ld_data_v_r_863_sv2v_reg;
  assign ld_data_v_r[862] = ld_data_v_r_862_sv2v_reg;
  assign ld_data_v_r[861] = ld_data_v_r_861_sv2v_reg;
  assign ld_data_v_r[860] = ld_data_v_r_860_sv2v_reg;
  assign ld_data_v_r[859] = ld_data_v_r_859_sv2v_reg;
  assign ld_data_v_r[858] = ld_data_v_r_858_sv2v_reg;
  assign ld_data_v_r[857] = ld_data_v_r_857_sv2v_reg;
  assign ld_data_v_r[856] = ld_data_v_r_856_sv2v_reg;
  assign ld_data_v_r[855] = ld_data_v_r_855_sv2v_reg;
  assign ld_data_v_r[854] = ld_data_v_r_854_sv2v_reg;
  assign ld_data_v_r[853] = ld_data_v_r_853_sv2v_reg;
  assign ld_data_v_r[852] = ld_data_v_r_852_sv2v_reg;
  assign ld_data_v_r[851] = ld_data_v_r_851_sv2v_reg;
  assign ld_data_v_r[850] = ld_data_v_r_850_sv2v_reg;
  assign ld_data_v_r[849] = ld_data_v_r_849_sv2v_reg;
  assign ld_data_v_r[848] = ld_data_v_r_848_sv2v_reg;
  assign ld_data_v_r[847] = ld_data_v_r_847_sv2v_reg;
  assign ld_data_v_r[846] = ld_data_v_r_846_sv2v_reg;
  assign ld_data_v_r[845] = ld_data_v_r_845_sv2v_reg;
  assign ld_data_v_r[844] = ld_data_v_r_844_sv2v_reg;
  assign ld_data_v_r[843] = ld_data_v_r_843_sv2v_reg;
  assign ld_data_v_r[842] = ld_data_v_r_842_sv2v_reg;
  assign ld_data_v_r[841] = ld_data_v_r_841_sv2v_reg;
  assign ld_data_v_r[840] = ld_data_v_r_840_sv2v_reg;
  assign ld_data_v_r[839] = ld_data_v_r_839_sv2v_reg;
  assign ld_data_v_r[838] = ld_data_v_r_838_sv2v_reg;
  assign ld_data_v_r[837] = ld_data_v_r_837_sv2v_reg;
  assign ld_data_v_r[836] = ld_data_v_r_836_sv2v_reg;
  assign ld_data_v_r[835] = ld_data_v_r_835_sv2v_reg;
  assign ld_data_v_r[834] = ld_data_v_r_834_sv2v_reg;
  assign ld_data_v_r[833] = ld_data_v_r_833_sv2v_reg;
  assign ld_data_v_r[832] = ld_data_v_r_832_sv2v_reg;
  assign ld_data_v_r[831] = ld_data_v_r_831_sv2v_reg;
  assign ld_data_v_r[830] = ld_data_v_r_830_sv2v_reg;
  assign ld_data_v_r[829] = ld_data_v_r_829_sv2v_reg;
  assign ld_data_v_r[828] = ld_data_v_r_828_sv2v_reg;
  assign ld_data_v_r[827] = ld_data_v_r_827_sv2v_reg;
  assign ld_data_v_r[826] = ld_data_v_r_826_sv2v_reg;
  assign ld_data_v_r[825] = ld_data_v_r_825_sv2v_reg;
  assign ld_data_v_r[824] = ld_data_v_r_824_sv2v_reg;
  assign ld_data_v_r[823] = ld_data_v_r_823_sv2v_reg;
  assign ld_data_v_r[822] = ld_data_v_r_822_sv2v_reg;
  assign ld_data_v_r[821] = ld_data_v_r_821_sv2v_reg;
  assign ld_data_v_r[820] = ld_data_v_r_820_sv2v_reg;
  assign ld_data_v_r[819] = ld_data_v_r_819_sv2v_reg;
  assign ld_data_v_r[818] = ld_data_v_r_818_sv2v_reg;
  assign ld_data_v_r[817] = ld_data_v_r_817_sv2v_reg;
  assign ld_data_v_r[816] = ld_data_v_r_816_sv2v_reg;
  assign ld_data_v_r[815] = ld_data_v_r_815_sv2v_reg;
  assign ld_data_v_r[814] = ld_data_v_r_814_sv2v_reg;
  assign ld_data_v_r[813] = ld_data_v_r_813_sv2v_reg;
  assign ld_data_v_r[812] = ld_data_v_r_812_sv2v_reg;
  assign ld_data_v_r[811] = ld_data_v_r_811_sv2v_reg;
  assign ld_data_v_r[810] = ld_data_v_r_810_sv2v_reg;
  assign ld_data_v_r[809] = ld_data_v_r_809_sv2v_reg;
  assign ld_data_v_r[808] = ld_data_v_r_808_sv2v_reg;
  assign ld_data_v_r[807] = ld_data_v_r_807_sv2v_reg;
  assign ld_data_v_r[806] = ld_data_v_r_806_sv2v_reg;
  assign ld_data_v_r[805] = ld_data_v_r_805_sv2v_reg;
  assign ld_data_v_r[804] = ld_data_v_r_804_sv2v_reg;
  assign ld_data_v_r[803] = ld_data_v_r_803_sv2v_reg;
  assign ld_data_v_r[802] = ld_data_v_r_802_sv2v_reg;
  assign ld_data_v_r[801] = ld_data_v_r_801_sv2v_reg;
  assign ld_data_v_r[800] = ld_data_v_r_800_sv2v_reg;
  assign ld_data_v_r[799] = ld_data_v_r_799_sv2v_reg;
  assign ld_data_v_r[798] = ld_data_v_r_798_sv2v_reg;
  assign ld_data_v_r[797] = ld_data_v_r_797_sv2v_reg;
  assign ld_data_v_r[796] = ld_data_v_r_796_sv2v_reg;
  assign ld_data_v_r[795] = ld_data_v_r_795_sv2v_reg;
  assign ld_data_v_r[794] = ld_data_v_r_794_sv2v_reg;
  assign ld_data_v_r[793] = ld_data_v_r_793_sv2v_reg;
  assign ld_data_v_r[792] = ld_data_v_r_792_sv2v_reg;
  assign ld_data_v_r[791] = ld_data_v_r_791_sv2v_reg;
  assign ld_data_v_r[790] = ld_data_v_r_790_sv2v_reg;
  assign ld_data_v_r[789] = ld_data_v_r_789_sv2v_reg;
  assign ld_data_v_r[788] = ld_data_v_r_788_sv2v_reg;
  assign ld_data_v_r[787] = ld_data_v_r_787_sv2v_reg;
  assign ld_data_v_r[786] = ld_data_v_r_786_sv2v_reg;
  assign ld_data_v_r[785] = ld_data_v_r_785_sv2v_reg;
  assign ld_data_v_r[784] = ld_data_v_r_784_sv2v_reg;
  assign ld_data_v_r[783] = ld_data_v_r_783_sv2v_reg;
  assign ld_data_v_r[782] = ld_data_v_r_782_sv2v_reg;
  assign ld_data_v_r[781] = ld_data_v_r_781_sv2v_reg;
  assign ld_data_v_r[780] = ld_data_v_r_780_sv2v_reg;
  assign ld_data_v_r[779] = ld_data_v_r_779_sv2v_reg;
  assign ld_data_v_r[778] = ld_data_v_r_778_sv2v_reg;
  assign ld_data_v_r[777] = ld_data_v_r_777_sv2v_reg;
  assign ld_data_v_r[776] = ld_data_v_r_776_sv2v_reg;
  assign ld_data_v_r[775] = ld_data_v_r_775_sv2v_reg;
  assign ld_data_v_r[774] = ld_data_v_r_774_sv2v_reg;
  assign ld_data_v_r[773] = ld_data_v_r_773_sv2v_reg;
  assign ld_data_v_r[772] = ld_data_v_r_772_sv2v_reg;
  assign ld_data_v_r[771] = ld_data_v_r_771_sv2v_reg;
  assign ld_data_v_r[770] = ld_data_v_r_770_sv2v_reg;
  assign ld_data_v_r[769] = ld_data_v_r_769_sv2v_reg;
  assign ld_data_v_r[768] = ld_data_v_r_768_sv2v_reg;
  assign ld_data_v_r[767] = ld_data_v_r_767_sv2v_reg;
  assign ld_data_v_r[766] = ld_data_v_r_766_sv2v_reg;
  assign ld_data_v_r[765] = ld_data_v_r_765_sv2v_reg;
  assign ld_data_v_r[764] = ld_data_v_r_764_sv2v_reg;
  assign ld_data_v_r[763] = ld_data_v_r_763_sv2v_reg;
  assign ld_data_v_r[762] = ld_data_v_r_762_sv2v_reg;
  assign ld_data_v_r[761] = ld_data_v_r_761_sv2v_reg;
  assign ld_data_v_r[760] = ld_data_v_r_760_sv2v_reg;
  assign ld_data_v_r[759] = ld_data_v_r_759_sv2v_reg;
  assign ld_data_v_r[758] = ld_data_v_r_758_sv2v_reg;
  assign ld_data_v_r[757] = ld_data_v_r_757_sv2v_reg;
  assign ld_data_v_r[756] = ld_data_v_r_756_sv2v_reg;
  assign ld_data_v_r[755] = ld_data_v_r_755_sv2v_reg;
  assign ld_data_v_r[754] = ld_data_v_r_754_sv2v_reg;
  assign ld_data_v_r[753] = ld_data_v_r_753_sv2v_reg;
  assign ld_data_v_r[752] = ld_data_v_r_752_sv2v_reg;
  assign ld_data_v_r[751] = ld_data_v_r_751_sv2v_reg;
  assign ld_data_v_r[750] = ld_data_v_r_750_sv2v_reg;
  assign ld_data_v_r[749] = ld_data_v_r_749_sv2v_reg;
  assign ld_data_v_r[748] = ld_data_v_r_748_sv2v_reg;
  assign ld_data_v_r[747] = ld_data_v_r_747_sv2v_reg;
  assign ld_data_v_r[746] = ld_data_v_r_746_sv2v_reg;
  assign ld_data_v_r[745] = ld_data_v_r_745_sv2v_reg;
  assign ld_data_v_r[744] = ld_data_v_r_744_sv2v_reg;
  assign ld_data_v_r[743] = ld_data_v_r_743_sv2v_reg;
  assign ld_data_v_r[742] = ld_data_v_r_742_sv2v_reg;
  assign ld_data_v_r[741] = ld_data_v_r_741_sv2v_reg;
  assign ld_data_v_r[740] = ld_data_v_r_740_sv2v_reg;
  assign ld_data_v_r[739] = ld_data_v_r_739_sv2v_reg;
  assign ld_data_v_r[738] = ld_data_v_r_738_sv2v_reg;
  assign ld_data_v_r[737] = ld_data_v_r_737_sv2v_reg;
  assign ld_data_v_r[736] = ld_data_v_r_736_sv2v_reg;
  assign ld_data_v_r[735] = ld_data_v_r_735_sv2v_reg;
  assign ld_data_v_r[734] = ld_data_v_r_734_sv2v_reg;
  assign ld_data_v_r[733] = ld_data_v_r_733_sv2v_reg;
  assign ld_data_v_r[732] = ld_data_v_r_732_sv2v_reg;
  assign ld_data_v_r[731] = ld_data_v_r_731_sv2v_reg;
  assign ld_data_v_r[730] = ld_data_v_r_730_sv2v_reg;
  assign ld_data_v_r[729] = ld_data_v_r_729_sv2v_reg;
  assign ld_data_v_r[728] = ld_data_v_r_728_sv2v_reg;
  assign ld_data_v_r[727] = ld_data_v_r_727_sv2v_reg;
  assign ld_data_v_r[726] = ld_data_v_r_726_sv2v_reg;
  assign ld_data_v_r[725] = ld_data_v_r_725_sv2v_reg;
  assign ld_data_v_r[724] = ld_data_v_r_724_sv2v_reg;
  assign ld_data_v_r[723] = ld_data_v_r_723_sv2v_reg;
  assign ld_data_v_r[722] = ld_data_v_r_722_sv2v_reg;
  assign ld_data_v_r[721] = ld_data_v_r_721_sv2v_reg;
  assign ld_data_v_r[720] = ld_data_v_r_720_sv2v_reg;
  assign ld_data_v_r[719] = ld_data_v_r_719_sv2v_reg;
  assign ld_data_v_r[718] = ld_data_v_r_718_sv2v_reg;
  assign ld_data_v_r[717] = ld_data_v_r_717_sv2v_reg;
  assign ld_data_v_r[716] = ld_data_v_r_716_sv2v_reg;
  assign ld_data_v_r[715] = ld_data_v_r_715_sv2v_reg;
  assign ld_data_v_r[714] = ld_data_v_r_714_sv2v_reg;
  assign ld_data_v_r[713] = ld_data_v_r_713_sv2v_reg;
  assign ld_data_v_r[712] = ld_data_v_r_712_sv2v_reg;
  assign ld_data_v_r[711] = ld_data_v_r_711_sv2v_reg;
  assign ld_data_v_r[710] = ld_data_v_r_710_sv2v_reg;
  assign ld_data_v_r[709] = ld_data_v_r_709_sv2v_reg;
  assign ld_data_v_r[708] = ld_data_v_r_708_sv2v_reg;
  assign ld_data_v_r[707] = ld_data_v_r_707_sv2v_reg;
  assign ld_data_v_r[706] = ld_data_v_r_706_sv2v_reg;
  assign ld_data_v_r[705] = ld_data_v_r_705_sv2v_reg;
  assign ld_data_v_r[704] = ld_data_v_r_704_sv2v_reg;
  assign ld_data_v_r[703] = ld_data_v_r_703_sv2v_reg;
  assign ld_data_v_r[702] = ld_data_v_r_702_sv2v_reg;
  assign ld_data_v_r[701] = ld_data_v_r_701_sv2v_reg;
  assign ld_data_v_r[700] = ld_data_v_r_700_sv2v_reg;
  assign ld_data_v_r[699] = ld_data_v_r_699_sv2v_reg;
  assign ld_data_v_r[698] = ld_data_v_r_698_sv2v_reg;
  assign ld_data_v_r[697] = ld_data_v_r_697_sv2v_reg;
  assign ld_data_v_r[696] = ld_data_v_r_696_sv2v_reg;
  assign ld_data_v_r[695] = ld_data_v_r_695_sv2v_reg;
  assign ld_data_v_r[694] = ld_data_v_r_694_sv2v_reg;
  assign ld_data_v_r[693] = ld_data_v_r_693_sv2v_reg;
  assign ld_data_v_r[692] = ld_data_v_r_692_sv2v_reg;
  assign ld_data_v_r[691] = ld_data_v_r_691_sv2v_reg;
  assign ld_data_v_r[690] = ld_data_v_r_690_sv2v_reg;
  assign ld_data_v_r[689] = ld_data_v_r_689_sv2v_reg;
  assign ld_data_v_r[688] = ld_data_v_r_688_sv2v_reg;
  assign ld_data_v_r[687] = ld_data_v_r_687_sv2v_reg;
  assign ld_data_v_r[686] = ld_data_v_r_686_sv2v_reg;
  assign ld_data_v_r[685] = ld_data_v_r_685_sv2v_reg;
  assign ld_data_v_r[684] = ld_data_v_r_684_sv2v_reg;
  assign ld_data_v_r[683] = ld_data_v_r_683_sv2v_reg;
  assign ld_data_v_r[682] = ld_data_v_r_682_sv2v_reg;
  assign ld_data_v_r[681] = ld_data_v_r_681_sv2v_reg;
  assign ld_data_v_r[680] = ld_data_v_r_680_sv2v_reg;
  assign ld_data_v_r[679] = ld_data_v_r_679_sv2v_reg;
  assign ld_data_v_r[678] = ld_data_v_r_678_sv2v_reg;
  assign ld_data_v_r[677] = ld_data_v_r_677_sv2v_reg;
  assign ld_data_v_r[676] = ld_data_v_r_676_sv2v_reg;
  assign ld_data_v_r[675] = ld_data_v_r_675_sv2v_reg;
  assign ld_data_v_r[674] = ld_data_v_r_674_sv2v_reg;
  assign ld_data_v_r[673] = ld_data_v_r_673_sv2v_reg;
  assign ld_data_v_r[672] = ld_data_v_r_672_sv2v_reg;
  assign ld_data_v_r[671] = ld_data_v_r_671_sv2v_reg;
  assign ld_data_v_r[670] = ld_data_v_r_670_sv2v_reg;
  assign ld_data_v_r[669] = ld_data_v_r_669_sv2v_reg;
  assign ld_data_v_r[668] = ld_data_v_r_668_sv2v_reg;
  assign ld_data_v_r[667] = ld_data_v_r_667_sv2v_reg;
  assign ld_data_v_r[666] = ld_data_v_r_666_sv2v_reg;
  assign ld_data_v_r[665] = ld_data_v_r_665_sv2v_reg;
  assign ld_data_v_r[664] = ld_data_v_r_664_sv2v_reg;
  assign ld_data_v_r[663] = ld_data_v_r_663_sv2v_reg;
  assign ld_data_v_r[662] = ld_data_v_r_662_sv2v_reg;
  assign ld_data_v_r[661] = ld_data_v_r_661_sv2v_reg;
  assign ld_data_v_r[660] = ld_data_v_r_660_sv2v_reg;
  assign ld_data_v_r[659] = ld_data_v_r_659_sv2v_reg;
  assign ld_data_v_r[658] = ld_data_v_r_658_sv2v_reg;
  assign ld_data_v_r[657] = ld_data_v_r_657_sv2v_reg;
  assign ld_data_v_r[656] = ld_data_v_r_656_sv2v_reg;
  assign ld_data_v_r[655] = ld_data_v_r_655_sv2v_reg;
  assign ld_data_v_r[654] = ld_data_v_r_654_sv2v_reg;
  assign ld_data_v_r[653] = ld_data_v_r_653_sv2v_reg;
  assign ld_data_v_r[652] = ld_data_v_r_652_sv2v_reg;
  assign ld_data_v_r[651] = ld_data_v_r_651_sv2v_reg;
  assign ld_data_v_r[650] = ld_data_v_r_650_sv2v_reg;
  assign ld_data_v_r[649] = ld_data_v_r_649_sv2v_reg;
  assign ld_data_v_r[648] = ld_data_v_r_648_sv2v_reg;
  assign ld_data_v_r[647] = ld_data_v_r_647_sv2v_reg;
  assign ld_data_v_r[646] = ld_data_v_r_646_sv2v_reg;
  assign ld_data_v_r[645] = ld_data_v_r_645_sv2v_reg;
  assign ld_data_v_r[644] = ld_data_v_r_644_sv2v_reg;
  assign ld_data_v_r[643] = ld_data_v_r_643_sv2v_reg;
  assign ld_data_v_r[642] = ld_data_v_r_642_sv2v_reg;
  assign ld_data_v_r[641] = ld_data_v_r_641_sv2v_reg;
  assign ld_data_v_r[640] = ld_data_v_r_640_sv2v_reg;
  assign ld_data_v_r[639] = ld_data_v_r_639_sv2v_reg;
  assign ld_data_v_r[638] = ld_data_v_r_638_sv2v_reg;
  assign ld_data_v_r[637] = ld_data_v_r_637_sv2v_reg;
  assign ld_data_v_r[636] = ld_data_v_r_636_sv2v_reg;
  assign ld_data_v_r[635] = ld_data_v_r_635_sv2v_reg;
  assign ld_data_v_r[634] = ld_data_v_r_634_sv2v_reg;
  assign ld_data_v_r[633] = ld_data_v_r_633_sv2v_reg;
  assign ld_data_v_r[632] = ld_data_v_r_632_sv2v_reg;
  assign ld_data_v_r[631] = ld_data_v_r_631_sv2v_reg;
  assign ld_data_v_r[630] = ld_data_v_r_630_sv2v_reg;
  assign ld_data_v_r[629] = ld_data_v_r_629_sv2v_reg;
  assign ld_data_v_r[628] = ld_data_v_r_628_sv2v_reg;
  assign ld_data_v_r[627] = ld_data_v_r_627_sv2v_reg;
  assign ld_data_v_r[626] = ld_data_v_r_626_sv2v_reg;
  assign ld_data_v_r[625] = ld_data_v_r_625_sv2v_reg;
  assign ld_data_v_r[624] = ld_data_v_r_624_sv2v_reg;
  assign ld_data_v_r[623] = ld_data_v_r_623_sv2v_reg;
  assign ld_data_v_r[622] = ld_data_v_r_622_sv2v_reg;
  assign ld_data_v_r[621] = ld_data_v_r_621_sv2v_reg;
  assign ld_data_v_r[620] = ld_data_v_r_620_sv2v_reg;
  assign ld_data_v_r[619] = ld_data_v_r_619_sv2v_reg;
  assign ld_data_v_r[618] = ld_data_v_r_618_sv2v_reg;
  assign ld_data_v_r[617] = ld_data_v_r_617_sv2v_reg;
  assign ld_data_v_r[616] = ld_data_v_r_616_sv2v_reg;
  assign ld_data_v_r[615] = ld_data_v_r_615_sv2v_reg;
  assign ld_data_v_r[614] = ld_data_v_r_614_sv2v_reg;
  assign ld_data_v_r[613] = ld_data_v_r_613_sv2v_reg;
  assign ld_data_v_r[612] = ld_data_v_r_612_sv2v_reg;
  assign ld_data_v_r[611] = ld_data_v_r_611_sv2v_reg;
  assign ld_data_v_r[610] = ld_data_v_r_610_sv2v_reg;
  assign ld_data_v_r[609] = ld_data_v_r_609_sv2v_reg;
  assign ld_data_v_r[608] = ld_data_v_r_608_sv2v_reg;
  assign ld_data_v_r[607] = ld_data_v_r_607_sv2v_reg;
  assign ld_data_v_r[606] = ld_data_v_r_606_sv2v_reg;
  assign ld_data_v_r[605] = ld_data_v_r_605_sv2v_reg;
  assign ld_data_v_r[604] = ld_data_v_r_604_sv2v_reg;
  assign ld_data_v_r[603] = ld_data_v_r_603_sv2v_reg;
  assign ld_data_v_r[602] = ld_data_v_r_602_sv2v_reg;
  assign ld_data_v_r[601] = ld_data_v_r_601_sv2v_reg;
  assign ld_data_v_r[600] = ld_data_v_r_600_sv2v_reg;
  assign ld_data_v_r[599] = ld_data_v_r_599_sv2v_reg;
  assign ld_data_v_r[598] = ld_data_v_r_598_sv2v_reg;
  assign ld_data_v_r[597] = ld_data_v_r_597_sv2v_reg;
  assign ld_data_v_r[596] = ld_data_v_r_596_sv2v_reg;
  assign ld_data_v_r[595] = ld_data_v_r_595_sv2v_reg;
  assign ld_data_v_r[594] = ld_data_v_r_594_sv2v_reg;
  assign ld_data_v_r[593] = ld_data_v_r_593_sv2v_reg;
  assign ld_data_v_r[592] = ld_data_v_r_592_sv2v_reg;
  assign ld_data_v_r[591] = ld_data_v_r_591_sv2v_reg;
  assign ld_data_v_r[590] = ld_data_v_r_590_sv2v_reg;
  assign ld_data_v_r[589] = ld_data_v_r_589_sv2v_reg;
  assign ld_data_v_r[588] = ld_data_v_r_588_sv2v_reg;
  assign ld_data_v_r[587] = ld_data_v_r_587_sv2v_reg;
  assign ld_data_v_r[586] = ld_data_v_r_586_sv2v_reg;
  assign ld_data_v_r[585] = ld_data_v_r_585_sv2v_reg;
  assign ld_data_v_r[584] = ld_data_v_r_584_sv2v_reg;
  assign ld_data_v_r[583] = ld_data_v_r_583_sv2v_reg;
  assign ld_data_v_r[582] = ld_data_v_r_582_sv2v_reg;
  assign ld_data_v_r[581] = ld_data_v_r_581_sv2v_reg;
  assign ld_data_v_r[580] = ld_data_v_r_580_sv2v_reg;
  assign ld_data_v_r[579] = ld_data_v_r_579_sv2v_reg;
  assign ld_data_v_r[578] = ld_data_v_r_578_sv2v_reg;
  assign ld_data_v_r[577] = ld_data_v_r_577_sv2v_reg;
  assign ld_data_v_r[576] = ld_data_v_r_576_sv2v_reg;
  assign ld_data_v_r[575] = ld_data_v_r_575_sv2v_reg;
  assign ld_data_v_r[574] = ld_data_v_r_574_sv2v_reg;
  assign ld_data_v_r[573] = ld_data_v_r_573_sv2v_reg;
  assign ld_data_v_r[572] = ld_data_v_r_572_sv2v_reg;
  assign ld_data_v_r[571] = ld_data_v_r_571_sv2v_reg;
  assign ld_data_v_r[570] = ld_data_v_r_570_sv2v_reg;
  assign ld_data_v_r[569] = ld_data_v_r_569_sv2v_reg;
  assign ld_data_v_r[568] = ld_data_v_r_568_sv2v_reg;
  assign ld_data_v_r[567] = ld_data_v_r_567_sv2v_reg;
  assign ld_data_v_r[566] = ld_data_v_r_566_sv2v_reg;
  assign ld_data_v_r[565] = ld_data_v_r_565_sv2v_reg;
  assign ld_data_v_r[564] = ld_data_v_r_564_sv2v_reg;
  assign ld_data_v_r[563] = ld_data_v_r_563_sv2v_reg;
  assign ld_data_v_r[562] = ld_data_v_r_562_sv2v_reg;
  assign ld_data_v_r[561] = ld_data_v_r_561_sv2v_reg;
  assign ld_data_v_r[560] = ld_data_v_r_560_sv2v_reg;
  assign ld_data_v_r[559] = ld_data_v_r_559_sv2v_reg;
  assign ld_data_v_r[558] = ld_data_v_r_558_sv2v_reg;
  assign ld_data_v_r[557] = ld_data_v_r_557_sv2v_reg;
  assign ld_data_v_r[556] = ld_data_v_r_556_sv2v_reg;
  assign ld_data_v_r[555] = ld_data_v_r_555_sv2v_reg;
  assign ld_data_v_r[554] = ld_data_v_r_554_sv2v_reg;
  assign ld_data_v_r[553] = ld_data_v_r_553_sv2v_reg;
  assign ld_data_v_r[552] = ld_data_v_r_552_sv2v_reg;
  assign ld_data_v_r[551] = ld_data_v_r_551_sv2v_reg;
  assign ld_data_v_r[550] = ld_data_v_r_550_sv2v_reg;
  assign ld_data_v_r[549] = ld_data_v_r_549_sv2v_reg;
  assign ld_data_v_r[548] = ld_data_v_r_548_sv2v_reg;
  assign ld_data_v_r[547] = ld_data_v_r_547_sv2v_reg;
  assign ld_data_v_r[546] = ld_data_v_r_546_sv2v_reg;
  assign ld_data_v_r[545] = ld_data_v_r_545_sv2v_reg;
  assign ld_data_v_r[544] = ld_data_v_r_544_sv2v_reg;
  assign ld_data_v_r[543] = ld_data_v_r_543_sv2v_reg;
  assign ld_data_v_r[542] = ld_data_v_r_542_sv2v_reg;
  assign ld_data_v_r[541] = ld_data_v_r_541_sv2v_reg;
  assign ld_data_v_r[540] = ld_data_v_r_540_sv2v_reg;
  assign ld_data_v_r[539] = ld_data_v_r_539_sv2v_reg;
  assign ld_data_v_r[538] = ld_data_v_r_538_sv2v_reg;
  assign ld_data_v_r[537] = ld_data_v_r_537_sv2v_reg;
  assign ld_data_v_r[536] = ld_data_v_r_536_sv2v_reg;
  assign ld_data_v_r[535] = ld_data_v_r_535_sv2v_reg;
  assign ld_data_v_r[534] = ld_data_v_r_534_sv2v_reg;
  assign ld_data_v_r[533] = ld_data_v_r_533_sv2v_reg;
  assign ld_data_v_r[532] = ld_data_v_r_532_sv2v_reg;
  assign ld_data_v_r[531] = ld_data_v_r_531_sv2v_reg;
  assign ld_data_v_r[530] = ld_data_v_r_530_sv2v_reg;
  assign ld_data_v_r[529] = ld_data_v_r_529_sv2v_reg;
  assign ld_data_v_r[528] = ld_data_v_r_528_sv2v_reg;
  assign ld_data_v_r[527] = ld_data_v_r_527_sv2v_reg;
  assign ld_data_v_r[526] = ld_data_v_r_526_sv2v_reg;
  assign ld_data_v_r[525] = ld_data_v_r_525_sv2v_reg;
  assign ld_data_v_r[524] = ld_data_v_r_524_sv2v_reg;
  assign ld_data_v_r[523] = ld_data_v_r_523_sv2v_reg;
  assign ld_data_v_r[522] = ld_data_v_r_522_sv2v_reg;
  assign ld_data_v_r[521] = ld_data_v_r_521_sv2v_reg;
  assign ld_data_v_r[520] = ld_data_v_r_520_sv2v_reg;
  assign ld_data_v_r[519] = ld_data_v_r_519_sv2v_reg;
  assign ld_data_v_r[518] = ld_data_v_r_518_sv2v_reg;
  assign ld_data_v_r[517] = ld_data_v_r_517_sv2v_reg;
  assign ld_data_v_r[516] = ld_data_v_r_516_sv2v_reg;
  assign ld_data_v_r[515] = ld_data_v_r_515_sv2v_reg;
  assign ld_data_v_r[514] = ld_data_v_r_514_sv2v_reg;
  assign ld_data_v_r[513] = ld_data_v_r_513_sv2v_reg;
  assign ld_data_v_r[512] = ld_data_v_r_512_sv2v_reg;
  assign ld_data_v_r[511] = ld_data_v_r_511_sv2v_reg;
  assign ld_data_v_r[510] = ld_data_v_r_510_sv2v_reg;
  assign ld_data_v_r[509] = ld_data_v_r_509_sv2v_reg;
  assign ld_data_v_r[508] = ld_data_v_r_508_sv2v_reg;
  assign ld_data_v_r[507] = ld_data_v_r_507_sv2v_reg;
  assign ld_data_v_r[506] = ld_data_v_r_506_sv2v_reg;
  assign ld_data_v_r[505] = ld_data_v_r_505_sv2v_reg;
  assign ld_data_v_r[504] = ld_data_v_r_504_sv2v_reg;
  assign ld_data_v_r[503] = ld_data_v_r_503_sv2v_reg;
  assign ld_data_v_r[502] = ld_data_v_r_502_sv2v_reg;
  assign ld_data_v_r[501] = ld_data_v_r_501_sv2v_reg;
  assign ld_data_v_r[500] = ld_data_v_r_500_sv2v_reg;
  assign ld_data_v_r[499] = ld_data_v_r_499_sv2v_reg;
  assign ld_data_v_r[498] = ld_data_v_r_498_sv2v_reg;
  assign ld_data_v_r[497] = ld_data_v_r_497_sv2v_reg;
  assign ld_data_v_r[496] = ld_data_v_r_496_sv2v_reg;
  assign ld_data_v_r[495] = ld_data_v_r_495_sv2v_reg;
  assign ld_data_v_r[494] = ld_data_v_r_494_sv2v_reg;
  assign ld_data_v_r[493] = ld_data_v_r_493_sv2v_reg;
  assign ld_data_v_r[492] = ld_data_v_r_492_sv2v_reg;
  assign ld_data_v_r[491] = ld_data_v_r_491_sv2v_reg;
  assign ld_data_v_r[490] = ld_data_v_r_490_sv2v_reg;
  assign ld_data_v_r[489] = ld_data_v_r_489_sv2v_reg;
  assign ld_data_v_r[488] = ld_data_v_r_488_sv2v_reg;
  assign ld_data_v_r[487] = ld_data_v_r_487_sv2v_reg;
  assign ld_data_v_r[486] = ld_data_v_r_486_sv2v_reg;
  assign ld_data_v_r[485] = ld_data_v_r_485_sv2v_reg;
  assign ld_data_v_r[484] = ld_data_v_r_484_sv2v_reg;
  assign ld_data_v_r[483] = ld_data_v_r_483_sv2v_reg;
  assign ld_data_v_r[482] = ld_data_v_r_482_sv2v_reg;
  assign ld_data_v_r[481] = ld_data_v_r_481_sv2v_reg;
  assign ld_data_v_r[480] = ld_data_v_r_480_sv2v_reg;
  assign ld_data_v_r[479] = ld_data_v_r_479_sv2v_reg;
  assign ld_data_v_r[478] = ld_data_v_r_478_sv2v_reg;
  assign ld_data_v_r[477] = ld_data_v_r_477_sv2v_reg;
  assign ld_data_v_r[476] = ld_data_v_r_476_sv2v_reg;
  assign ld_data_v_r[475] = ld_data_v_r_475_sv2v_reg;
  assign ld_data_v_r[474] = ld_data_v_r_474_sv2v_reg;
  assign ld_data_v_r[473] = ld_data_v_r_473_sv2v_reg;
  assign ld_data_v_r[472] = ld_data_v_r_472_sv2v_reg;
  assign ld_data_v_r[471] = ld_data_v_r_471_sv2v_reg;
  assign ld_data_v_r[470] = ld_data_v_r_470_sv2v_reg;
  assign ld_data_v_r[469] = ld_data_v_r_469_sv2v_reg;
  assign ld_data_v_r[468] = ld_data_v_r_468_sv2v_reg;
  assign ld_data_v_r[467] = ld_data_v_r_467_sv2v_reg;
  assign ld_data_v_r[466] = ld_data_v_r_466_sv2v_reg;
  assign ld_data_v_r[465] = ld_data_v_r_465_sv2v_reg;
  assign ld_data_v_r[464] = ld_data_v_r_464_sv2v_reg;
  assign ld_data_v_r[463] = ld_data_v_r_463_sv2v_reg;
  assign ld_data_v_r[462] = ld_data_v_r_462_sv2v_reg;
  assign ld_data_v_r[461] = ld_data_v_r_461_sv2v_reg;
  assign ld_data_v_r[460] = ld_data_v_r_460_sv2v_reg;
  assign ld_data_v_r[459] = ld_data_v_r_459_sv2v_reg;
  assign ld_data_v_r[458] = ld_data_v_r_458_sv2v_reg;
  assign ld_data_v_r[457] = ld_data_v_r_457_sv2v_reg;
  assign ld_data_v_r[456] = ld_data_v_r_456_sv2v_reg;
  assign ld_data_v_r[455] = ld_data_v_r_455_sv2v_reg;
  assign ld_data_v_r[454] = ld_data_v_r_454_sv2v_reg;
  assign ld_data_v_r[453] = ld_data_v_r_453_sv2v_reg;
  assign ld_data_v_r[452] = ld_data_v_r_452_sv2v_reg;
  assign ld_data_v_r[451] = ld_data_v_r_451_sv2v_reg;
  assign ld_data_v_r[450] = ld_data_v_r_450_sv2v_reg;
  assign ld_data_v_r[449] = ld_data_v_r_449_sv2v_reg;
  assign ld_data_v_r[448] = ld_data_v_r_448_sv2v_reg;
  assign ld_data_v_r[447] = ld_data_v_r_447_sv2v_reg;
  assign ld_data_v_r[446] = ld_data_v_r_446_sv2v_reg;
  assign ld_data_v_r[445] = ld_data_v_r_445_sv2v_reg;
  assign ld_data_v_r[444] = ld_data_v_r_444_sv2v_reg;
  assign ld_data_v_r[443] = ld_data_v_r_443_sv2v_reg;
  assign ld_data_v_r[442] = ld_data_v_r_442_sv2v_reg;
  assign ld_data_v_r[441] = ld_data_v_r_441_sv2v_reg;
  assign ld_data_v_r[440] = ld_data_v_r_440_sv2v_reg;
  assign ld_data_v_r[439] = ld_data_v_r_439_sv2v_reg;
  assign ld_data_v_r[438] = ld_data_v_r_438_sv2v_reg;
  assign ld_data_v_r[437] = ld_data_v_r_437_sv2v_reg;
  assign ld_data_v_r[436] = ld_data_v_r_436_sv2v_reg;
  assign ld_data_v_r[435] = ld_data_v_r_435_sv2v_reg;
  assign ld_data_v_r[434] = ld_data_v_r_434_sv2v_reg;
  assign ld_data_v_r[433] = ld_data_v_r_433_sv2v_reg;
  assign ld_data_v_r[432] = ld_data_v_r_432_sv2v_reg;
  assign ld_data_v_r[431] = ld_data_v_r_431_sv2v_reg;
  assign ld_data_v_r[430] = ld_data_v_r_430_sv2v_reg;
  assign ld_data_v_r[429] = ld_data_v_r_429_sv2v_reg;
  assign ld_data_v_r[428] = ld_data_v_r_428_sv2v_reg;
  assign ld_data_v_r[427] = ld_data_v_r_427_sv2v_reg;
  assign ld_data_v_r[426] = ld_data_v_r_426_sv2v_reg;
  assign ld_data_v_r[425] = ld_data_v_r_425_sv2v_reg;
  assign ld_data_v_r[424] = ld_data_v_r_424_sv2v_reg;
  assign ld_data_v_r[423] = ld_data_v_r_423_sv2v_reg;
  assign ld_data_v_r[422] = ld_data_v_r_422_sv2v_reg;
  assign ld_data_v_r[421] = ld_data_v_r_421_sv2v_reg;
  assign ld_data_v_r[420] = ld_data_v_r_420_sv2v_reg;
  assign ld_data_v_r[419] = ld_data_v_r_419_sv2v_reg;
  assign ld_data_v_r[418] = ld_data_v_r_418_sv2v_reg;
  assign ld_data_v_r[417] = ld_data_v_r_417_sv2v_reg;
  assign ld_data_v_r[416] = ld_data_v_r_416_sv2v_reg;
  assign ld_data_v_r[415] = ld_data_v_r_415_sv2v_reg;
  assign ld_data_v_r[414] = ld_data_v_r_414_sv2v_reg;
  assign ld_data_v_r[413] = ld_data_v_r_413_sv2v_reg;
  assign ld_data_v_r[412] = ld_data_v_r_412_sv2v_reg;
  assign ld_data_v_r[411] = ld_data_v_r_411_sv2v_reg;
  assign ld_data_v_r[410] = ld_data_v_r_410_sv2v_reg;
  assign ld_data_v_r[409] = ld_data_v_r_409_sv2v_reg;
  assign ld_data_v_r[408] = ld_data_v_r_408_sv2v_reg;
  assign ld_data_v_r[407] = ld_data_v_r_407_sv2v_reg;
  assign ld_data_v_r[406] = ld_data_v_r_406_sv2v_reg;
  assign ld_data_v_r[405] = ld_data_v_r_405_sv2v_reg;
  assign ld_data_v_r[404] = ld_data_v_r_404_sv2v_reg;
  assign ld_data_v_r[403] = ld_data_v_r_403_sv2v_reg;
  assign ld_data_v_r[402] = ld_data_v_r_402_sv2v_reg;
  assign ld_data_v_r[401] = ld_data_v_r_401_sv2v_reg;
  assign ld_data_v_r[400] = ld_data_v_r_400_sv2v_reg;
  assign ld_data_v_r[399] = ld_data_v_r_399_sv2v_reg;
  assign ld_data_v_r[398] = ld_data_v_r_398_sv2v_reg;
  assign ld_data_v_r[397] = ld_data_v_r_397_sv2v_reg;
  assign ld_data_v_r[396] = ld_data_v_r_396_sv2v_reg;
  assign ld_data_v_r[395] = ld_data_v_r_395_sv2v_reg;
  assign ld_data_v_r[394] = ld_data_v_r_394_sv2v_reg;
  assign ld_data_v_r[393] = ld_data_v_r_393_sv2v_reg;
  assign ld_data_v_r[392] = ld_data_v_r_392_sv2v_reg;
  assign ld_data_v_r[391] = ld_data_v_r_391_sv2v_reg;
  assign ld_data_v_r[390] = ld_data_v_r_390_sv2v_reg;
  assign ld_data_v_r[389] = ld_data_v_r_389_sv2v_reg;
  assign ld_data_v_r[388] = ld_data_v_r_388_sv2v_reg;
  assign ld_data_v_r[387] = ld_data_v_r_387_sv2v_reg;
  assign ld_data_v_r[386] = ld_data_v_r_386_sv2v_reg;
  assign ld_data_v_r[385] = ld_data_v_r_385_sv2v_reg;
  assign ld_data_v_r[384] = ld_data_v_r_384_sv2v_reg;
  assign ld_data_v_r[383] = ld_data_v_r_383_sv2v_reg;
  assign ld_data_v_r[382] = ld_data_v_r_382_sv2v_reg;
  assign ld_data_v_r[381] = ld_data_v_r_381_sv2v_reg;
  assign ld_data_v_r[380] = ld_data_v_r_380_sv2v_reg;
  assign ld_data_v_r[379] = ld_data_v_r_379_sv2v_reg;
  assign ld_data_v_r[378] = ld_data_v_r_378_sv2v_reg;
  assign ld_data_v_r[377] = ld_data_v_r_377_sv2v_reg;
  assign ld_data_v_r[376] = ld_data_v_r_376_sv2v_reg;
  assign ld_data_v_r[375] = ld_data_v_r_375_sv2v_reg;
  assign ld_data_v_r[374] = ld_data_v_r_374_sv2v_reg;
  assign ld_data_v_r[373] = ld_data_v_r_373_sv2v_reg;
  assign ld_data_v_r[372] = ld_data_v_r_372_sv2v_reg;
  assign ld_data_v_r[371] = ld_data_v_r_371_sv2v_reg;
  assign ld_data_v_r[370] = ld_data_v_r_370_sv2v_reg;
  assign ld_data_v_r[369] = ld_data_v_r_369_sv2v_reg;
  assign ld_data_v_r[368] = ld_data_v_r_368_sv2v_reg;
  assign ld_data_v_r[367] = ld_data_v_r_367_sv2v_reg;
  assign ld_data_v_r[366] = ld_data_v_r_366_sv2v_reg;
  assign ld_data_v_r[365] = ld_data_v_r_365_sv2v_reg;
  assign ld_data_v_r[364] = ld_data_v_r_364_sv2v_reg;
  assign ld_data_v_r[363] = ld_data_v_r_363_sv2v_reg;
  assign ld_data_v_r[362] = ld_data_v_r_362_sv2v_reg;
  assign ld_data_v_r[361] = ld_data_v_r_361_sv2v_reg;
  assign ld_data_v_r[360] = ld_data_v_r_360_sv2v_reg;
  assign ld_data_v_r[359] = ld_data_v_r_359_sv2v_reg;
  assign ld_data_v_r[358] = ld_data_v_r_358_sv2v_reg;
  assign ld_data_v_r[357] = ld_data_v_r_357_sv2v_reg;
  assign ld_data_v_r[356] = ld_data_v_r_356_sv2v_reg;
  assign ld_data_v_r[355] = ld_data_v_r_355_sv2v_reg;
  assign ld_data_v_r[354] = ld_data_v_r_354_sv2v_reg;
  assign ld_data_v_r[353] = ld_data_v_r_353_sv2v_reg;
  assign ld_data_v_r[352] = ld_data_v_r_352_sv2v_reg;
  assign ld_data_v_r[351] = ld_data_v_r_351_sv2v_reg;
  assign ld_data_v_r[350] = ld_data_v_r_350_sv2v_reg;
  assign ld_data_v_r[349] = ld_data_v_r_349_sv2v_reg;
  assign ld_data_v_r[348] = ld_data_v_r_348_sv2v_reg;
  assign ld_data_v_r[347] = ld_data_v_r_347_sv2v_reg;
  assign ld_data_v_r[346] = ld_data_v_r_346_sv2v_reg;
  assign ld_data_v_r[345] = ld_data_v_r_345_sv2v_reg;
  assign ld_data_v_r[344] = ld_data_v_r_344_sv2v_reg;
  assign ld_data_v_r[343] = ld_data_v_r_343_sv2v_reg;
  assign ld_data_v_r[342] = ld_data_v_r_342_sv2v_reg;
  assign ld_data_v_r[341] = ld_data_v_r_341_sv2v_reg;
  assign ld_data_v_r[340] = ld_data_v_r_340_sv2v_reg;
  assign ld_data_v_r[339] = ld_data_v_r_339_sv2v_reg;
  assign ld_data_v_r[338] = ld_data_v_r_338_sv2v_reg;
  assign ld_data_v_r[337] = ld_data_v_r_337_sv2v_reg;
  assign ld_data_v_r[336] = ld_data_v_r_336_sv2v_reg;
  assign ld_data_v_r[335] = ld_data_v_r_335_sv2v_reg;
  assign ld_data_v_r[334] = ld_data_v_r_334_sv2v_reg;
  assign ld_data_v_r[333] = ld_data_v_r_333_sv2v_reg;
  assign ld_data_v_r[332] = ld_data_v_r_332_sv2v_reg;
  assign ld_data_v_r[331] = ld_data_v_r_331_sv2v_reg;
  assign ld_data_v_r[330] = ld_data_v_r_330_sv2v_reg;
  assign ld_data_v_r[329] = ld_data_v_r_329_sv2v_reg;
  assign ld_data_v_r[328] = ld_data_v_r_328_sv2v_reg;
  assign ld_data_v_r[327] = ld_data_v_r_327_sv2v_reg;
  assign ld_data_v_r[326] = ld_data_v_r_326_sv2v_reg;
  assign ld_data_v_r[325] = ld_data_v_r_325_sv2v_reg;
  assign ld_data_v_r[324] = ld_data_v_r_324_sv2v_reg;
  assign ld_data_v_r[323] = ld_data_v_r_323_sv2v_reg;
  assign ld_data_v_r[322] = ld_data_v_r_322_sv2v_reg;
  assign ld_data_v_r[321] = ld_data_v_r_321_sv2v_reg;
  assign ld_data_v_r[320] = ld_data_v_r_320_sv2v_reg;
  assign ld_data_v_r[319] = ld_data_v_r_319_sv2v_reg;
  assign ld_data_v_r[318] = ld_data_v_r_318_sv2v_reg;
  assign ld_data_v_r[317] = ld_data_v_r_317_sv2v_reg;
  assign ld_data_v_r[316] = ld_data_v_r_316_sv2v_reg;
  assign ld_data_v_r[315] = ld_data_v_r_315_sv2v_reg;
  assign ld_data_v_r[314] = ld_data_v_r_314_sv2v_reg;
  assign ld_data_v_r[313] = ld_data_v_r_313_sv2v_reg;
  assign ld_data_v_r[312] = ld_data_v_r_312_sv2v_reg;
  assign ld_data_v_r[311] = ld_data_v_r_311_sv2v_reg;
  assign ld_data_v_r[310] = ld_data_v_r_310_sv2v_reg;
  assign ld_data_v_r[309] = ld_data_v_r_309_sv2v_reg;
  assign ld_data_v_r[308] = ld_data_v_r_308_sv2v_reg;
  assign ld_data_v_r[307] = ld_data_v_r_307_sv2v_reg;
  assign ld_data_v_r[306] = ld_data_v_r_306_sv2v_reg;
  assign ld_data_v_r[305] = ld_data_v_r_305_sv2v_reg;
  assign ld_data_v_r[304] = ld_data_v_r_304_sv2v_reg;
  assign ld_data_v_r[303] = ld_data_v_r_303_sv2v_reg;
  assign ld_data_v_r[302] = ld_data_v_r_302_sv2v_reg;
  assign ld_data_v_r[301] = ld_data_v_r_301_sv2v_reg;
  assign ld_data_v_r[300] = ld_data_v_r_300_sv2v_reg;
  assign ld_data_v_r[299] = ld_data_v_r_299_sv2v_reg;
  assign ld_data_v_r[298] = ld_data_v_r_298_sv2v_reg;
  assign ld_data_v_r[297] = ld_data_v_r_297_sv2v_reg;
  assign ld_data_v_r[296] = ld_data_v_r_296_sv2v_reg;
  assign ld_data_v_r[295] = ld_data_v_r_295_sv2v_reg;
  assign ld_data_v_r[294] = ld_data_v_r_294_sv2v_reg;
  assign ld_data_v_r[293] = ld_data_v_r_293_sv2v_reg;
  assign ld_data_v_r[292] = ld_data_v_r_292_sv2v_reg;
  assign ld_data_v_r[291] = ld_data_v_r_291_sv2v_reg;
  assign ld_data_v_r[290] = ld_data_v_r_290_sv2v_reg;
  assign ld_data_v_r[289] = ld_data_v_r_289_sv2v_reg;
  assign ld_data_v_r[288] = ld_data_v_r_288_sv2v_reg;
  assign ld_data_v_r[287] = ld_data_v_r_287_sv2v_reg;
  assign ld_data_v_r[286] = ld_data_v_r_286_sv2v_reg;
  assign ld_data_v_r[285] = ld_data_v_r_285_sv2v_reg;
  assign ld_data_v_r[284] = ld_data_v_r_284_sv2v_reg;
  assign ld_data_v_r[283] = ld_data_v_r_283_sv2v_reg;
  assign ld_data_v_r[282] = ld_data_v_r_282_sv2v_reg;
  assign ld_data_v_r[281] = ld_data_v_r_281_sv2v_reg;
  assign ld_data_v_r[280] = ld_data_v_r_280_sv2v_reg;
  assign ld_data_v_r[279] = ld_data_v_r_279_sv2v_reg;
  assign ld_data_v_r[278] = ld_data_v_r_278_sv2v_reg;
  assign ld_data_v_r[277] = ld_data_v_r_277_sv2v_reg;
  assign ld_data_v_r[276] = ld_data_v_r_276_sv2v_reg;
  assign ld_data_v_r[275] = ld_data_v_r_275_sv2v_reg;
  assign ld_data_v_r[274] = ld_data_v_r_274_sv2v_reg;
  assign ld_data_v_r[273] = ld_data_v_r_273_sv2v_reg;
  assign ld_data_v_r[272] = ld_data_v_r_272_sv2v_reg;
  assign ld_data_v_r[271] = ld_data_v_r_271_sv2v_reg;
  assign ld_data_v_r[270] = ld_data_v_r_270_sv2v_reg;
  assign ld_data_v_r[269] = ld_data_v_r_269_sv2v_reg;
  assign ld_data_v_r[268] = ld_data_v_r_268_sv2v_reg;
  assign ld_data_v_r[267] = ld_data_v_r_267_sv2v_reg;
  assign ld_data_v_r[266] = ld_data_v_r_266_sv2v_reg;
  assign ld_data_v_r[265] = ld_data_v_r_265_sv2v_reg;
  assign ld_data_v_r[264] = ld_data_v_r_264_sv2v_reg;
  assign ld_data_v_r[263] = ld_data_v_r_263_sv2v_reg;
  assign ld_data_v_r[262] = ld_data_v_r_262_sv2v_reg;
  assign ld_data_v_r[261] = ld_data_v_r_261_sv2v_reg;
  assign ld_data_v_r[260] = ld_data_v_r_260_sv2v_reg;
  assign ld_data_v_r[259] = ld_data_v_r_259_sv2v_reg;
  assign ld_data_v_r[258] = ld_data_v_r_258_sv2v_reg;
  assign ld_data_v_r[257] = ld_data_v_r_257_sv2v_reg;
  assign ld_data_v_r[256] = ld_data_v_r_256_sv2v_reg;
  assign ld_data_v_r[255] = ld_data_v_r_255_sv2v_reg;
  assign ld_data_v_r[254] = ld_data_v_r_254_sv2v_reg;
  assign ld_data_v_r[253] = ld_data_v_r_253_sv2v_reg;
  assign ld_data_v_r[252] = ld_data_v_r_252_sv2v_reg;
  assign ld_data_v_r[251] = ld_data_v_r_251_sv2v_reg;
  assign ld_data_v_r[250] = ld_data_v_r_250_sv2v_reg;
  assign ld_data_v_r[249] = ld_data_v_r_249_sv2v_reg;
  assign ld_data_v_r[248] = ld_data_v_r_248_sv2v_reg;
  assign ld_data_v_r[247] = ld_data_v_r_247_sv2v_reg;
  assign ld_data_v_r[246] = ld_data_v_r_246_sv2v_reg;
  assign ld_data_v_r[245] = ld_data_v_r_245_sv2v_reg;
  assign ld_data_v_r[244] = ld_data_v_r_244_sv2v_reg;
  assign ld_data_v_r[243] = ld_data_v_r_243_sv2v_reg;
  assign ld_data_v_r[242] = ld_data_v_r_242_sv2v_reg;
  assign ld_data_v_r[241] = ld_data_v_r_241_sv2v_reg;
  assign ld_data_v_r[240] = ld_data_v_r_240_sv2v_reg;
  assign ld_data_v_r[239] = ld_data_v_r_239_sv2v_reg;
  assign ld_data_v_r[238] = ld_data_v_r_238_sv2v_reg;
  assign ld_data_v_r[237] = ld_data_v_r_237_sv2v_reg;
  assign ld_data_v_r[236] = ld_data_v_r_236_sv2v_reg;
  assign ld_data_v_r[235] = ld_data_v_r_235_sv2v_reg;
  assign ld_data_v_r[234] = ld_data_v_r_234_sv2v_reg;
  assign ld_data_v_r[233] = ld_data_v_r_233_sv2v_reg;
  assign ld_data_v_r[232] = ld_data_v_r_232_sv2v_reg;
  assign ld_data_v_r[231] = ld_data_v_r_231_sv2v_reg;
  assign ld_data_v_r[230] = ld_data_v_r_230_sv2v_reg;
  assign ld_data_v_r[229] = ld_data_v_r_229_sv2v_reg;
  assign ld_data_v_r[228] = ld_data_v_r_228_sv2v_reg;
  assign ld_data_v_r[227] = ld_data_v_r_227_sv2v_reg;
  assign ld_data_v_r[226] = ld_data_v_r_226_sv2v_reg;
  assign ld_data_v_r[225] = ld_data_v_r_225_sv2v_reg;
  assign ld_data_v_r[224] = ld_data_v_r_224_sv2v_reg;
  assign ld_data_v_r[223] = ld_data_v_r_223_sv2v_reg;
  assign ld_data_v_r[222] = ld_data_v_r_222_sv2v_reg;
  assign ld_data_v_r[221] = ld_data_v_r_221_sv2v_reg;
  assign ld_data_v_r[220] = ld_data_v_r_220_sv2v_reg;
  assign ld_data_v_r[219] = ld_data_v_r_219_sv2v_reg;
  assign ld_data_v_r[218] = ld_data_v_r_218_sv2v_reg;
  assign ld_data_v_r[217] = ld_data_v_r_217_sv2v_reg;
  assign ld_data_v_r[216] = ld_data_v_r_216_sv2v_reg;
  assign ld_data_v_r[215] = ld_data_v_r_215_sv2v_reg;
  assign ld_data_v_r[214] = ld_data_v_r_214_sv2v_reg;
  assign ld_data_v_r[213] = ld_data_v_r_213_sv2v_reg;
  assign ld_data_v_r[212] = ld_data_v_r_212_sv2v_reg;
  assign ld_data_v_r[211] = ld_data_v_r_211_sv2v_reg;
  assign ld_data_v_r[210] = ld_data_v_r_210_sv2v_reg;
  assign ld_data_v_r[209] = ld_data_v_r_209_sv2v_reg;
  assign ld_data_v_r[208] = ld_data_v_r_208_sv2v_reg;
  assign ld_data_v_r[207] = ld_data_v_r_207_sv2v_reg;
  assign ld_data_v_r[206] = ld_data_v_r_206_sv2v_reg;
  assign ld_data_v_r[205] = ld_data_v_r_205_sv2v_reg;
  assign ld_data_v_r[204] = ld_data_v_r_204_sv2v_reg;
  assign ld_data_v_r[203] = ld_data_v_r_203_sv2v_reg;
  assign ld_data_v_r[202] = ld_data_v_r_202_sv2v_reg;
  assign ld_data_v_r[201] = ld_data_v_r_201_sv2v_reg;
  assign ld_data_v_r[200] = ld_data_v_r_200_sv2v_reg;
  assign ld_data_v_r[199] = ld_data_v_r_199_sv2v_reg;
  assign ld_data_v_r[198] = ld_data_v_r_198_sv2v_reg;
  assign ld_data_v_r[197] = ld_data_v_r_197_sv2v_reg;
  assign ld_data_v_r[196] = ld_data_v_r_196_sv2v_reg;
  assign ld_data_v_r[195] = ld_data_v_r_195_sv2v_reg;
  assign ld_data_v_r[194] = ld_data_v_r_194_sv2v_reg;
  assign ld_data_v_r[193] = ld_data_v_r_193_sv2v_reg;
  assign ld_data_v_r[192] = ld_data_v_r_192_sv2v_reg;
  assign ld_data_v_r[191] = ld_data_v_r_191_sv2v_reg;
  assign ld_data_v_r[190] = ld_data_v_r_190_sv2v_reg;
  assign ld_data_v_r[189] = ld_data_v_r_189_sv2v_reg;
  assign ld_data_v_r[188] = ld_data_v_r_188_sv2v_reg;
  assign ld_data_v_r[187] = ld_data_v_r_187_sv2v_reg;
  assign ld_data_v_r[186] = ld_data_v_r_186_sv2v_reg;
  assign ld_data_v_r[185] = ld_data_v_r_185_sv2v_reg;
  assign ld_data_v_r[184] = ld_data_v_r_184_sv2v_reg;
  assign ld_data_v_r[183] = ld_data_v_r_183_sv2v_reg;
  assign ld_data_v_r[182] = ld_data_v_r_182_sv2v_reg;
  assign ld_data_v_r[181] = ld_data_v_r_181_sv2v_reg;
  assign ld_data_v_r[180] = ld_data_v_r_180_sv2v_reg;
  assign ld_data_v_r[179] = ld_data_v_r_179_sv2v_reg;
  assign ld_data_v_r[178] = ld_data_v_r_178_sv2v_reg;
  assign ld_data_v_r[177] = ld_data_v_r_177_sv2v_reg;
  assign ld_data_v_r[176] = ld_data_v_r_176_sv2v_reg;
  assign ld_data_v_r[175] = ld_data_v_r_175_sv2v_reg;
  assign ld_data_v_r[174] = ld_data_v_r_174_sv2v_reg;
  assign ld_data_v_r[173] = ld_data_v_r_173_sv2v_reg;
  assign ld_data_v_r[172] = ld_data_v_r_172_sv2v_reg;
  assign ld_data_v_r[171] = ld_data_v_r_171_sv2v_reg;
  assign ld_data_v_r[170] = ld_data_v_r_170_sv2v_reg;
  assign ld_data_v_r[169] = ld_data_v_r_169_sv2v_reg;
  assign ld_data_v_r[168] = ld_data_v_r_168_sv2v_reg;
  assign ld_data_v_r[167] = ld_data_v_r_167_sv2v_reg;
  assign ld_data_v_r[166] = ld_data_v_r_166_sv2v_reg;
  assign ld_data_v_r[165] = ld_data_v_r_165_sv2v_reg;
  assign ld_data_v_r[164] = ld_data_v_r_164_sv2v_reg;
  assign ld_data_v_r[163] = ld_data_v_r_163_sv2v_reg;
  assign ld_data_v_r[162] = ld_data_v_r_162_sv2v_reg;
  assign ld_data_v_r[161] = ld_data_v_r_161_sv2v_reg;
  assign ld_data_v_r[160] = ld_data_v_r_160_sv2v_reg;
  assign ld_data_v_r[159] = ld_data_v_r_159_sv2v_reg;
  assign ld_data_v_r[158] = ld_data_v_r_158_sv2v_reg;
  assign ld_data_v_r[157] = ld_data_v_r_157_sv2v_reg;
  assign ld_data_v_r[156] = ld_data_v_r_156_sv2v_reg;
  assign ld_data_v_r[155] = ld_data_v_r_155_sv2v_reg;
  assign ld_data_v_r[154] = ld_data_v_r_154_sv2v_reg;
  assign ld_data_v_r[153] = ld_data_v_r_153_sv2v_reg;
  assign ld_data_v_r[152] = ld_data_v_r_152_sv2v_reg;
  assign ld_data_v_r[151] = ld_data_v_r_151_sv2v_reg;
  assign ld_data_v_r[150] = ld_data_v_r_150_sv2v_reg;
  assign ld_data_v_r[149] = ld_data_v_r_149_sv2v_reg;
  assign ld_data_v_r[148] = ld_data_v_r_148_sv2v_reg;
  assign ld_data_v_r[147] = ld_data_v_r_147_sv2v_reg;
  assign ld_data_v_r[146] = ld_data_v_r_146_sv2v_reg;
  assign ld_data_v_r[145] = ld_data_v_r_145_sv2v_reg;
  assign ld_data_v_r[144] = ld_data_v_r_144_sv2v_reg;
  assign ld_data_v_r[143] = ld_data_v_r_143_sv2v_reg;
  assign ld_data_v_r[142] = ld_data_v_r_142_sv2v_reg;
  assign ld_data_v_r[141] = ld_data_v_r_141_sv2v_reg;
  assign ld_data_v_r[140] = ld_data_v_r_140_sv2v_reg;
  assign ld_data_v_r[139] = ld_data_v_r_139_sv2v_reg;
  assign ld_data_v_r[138] = ld_data_v_r_138_sv2v_reg;
  assign ld_data_v_r[137] = ld_data_v_r_137_sv2v_reg;
  assign ld_data_v_r[136] = ld_data_v_r_136_sv2v_reg;
  assign ld_data_v_r[135] = ld_data_v_r_135_sv2v_reg;
  assign ld_data_v_r[134] = ld_data_v_r_134_sv2v_reg;
  assign ld_data_v_r[133] = ld_data_v_r_133_sv2v_reg;
  assign ld_data_v_r[132] = ld_data_v_r_132_sv2v_reg;
  assign ld_data_v_r[131] = ld_data_v_r_131_sv2v_reg;
  assign ld_data_v_r[130] = ld_data_v_r_130_sv2v_reg;
  assign ld_data_v_r[129] = ld_data_v_r_129_sv2v_reg;
  assign ld_data_v_r[128] = ld_data_v_r_128_sv2v_reg;
  assign ld_data_v_r[127] = ld_data_v_r_127_sv2v_reg;
  assign ld_data_v_r[126] = ld_data_v_r_126_sv2v_reg;
  assign ld_data_v_r[125] = ld_data_v_r_125_sv2v_reg;
  assign ld_data_v_r[124] = ld_data_v_r_124_sv2v_reg;
  assign ld_data_v_r[123] = ld_data_v_r_123_sv2v_reg;
  assign ld_data_v_r[122] = ld_data_v_r_122_sv2v_reg;
  assign ld_data_v_r[121] = ld_data_v_r_121_sv2v_reg;
  assign ld_data_v_r[120] = ld_data_v_r_120_sv2v_reg;
  assign ld_data_v_r[119] = ld_data_v_r_119_sv2v_reg;
  assign ld_data_v_r[118] = ld_data_v_r_118_sv2v_reg;
  assign ld_data_v_r[117] = ld_data_v_r_117_sv2v_reg;
  assign ld_data_v_r[116] = ld_data_v_r_116_sv2v_reg;
  assign ld_data_v_r[115] = ld_data_v_r_115_sv2v_reg;
  assign ld_data_v_r[114] = ld_data_v_r_114_sv2v_reg;
  assign ld_data_v_r[113] = ld_data_v_r_113_sv2v_reg;
  assign ld_data_v_r[112] = ld_data_v_r_112_sv2v_reg;
  assign ld_data_v_r[111] = ld_data_v_r_111_sv2v_reg;
  assign ld_data_v_r[110] = ld_data_v_r_110_sv2v_reg;
  assign ld_data_v_r[109] = ld_data_v_r_109_sv2v_reg;
  assign ld_data_v_r[108] = ld_data_v_r_108_sv2v_reg;
  assign ld_data_v_r[107] = ld_data_v_r_107_sv2v_reg;
  assign ld_data_v_r[106] = ld_data_v_r_106_sv2v_reg;
  assign ld_data_v_r[105] = ld_data_v_r_105_sv2v_reg;
  assign ld_data_v_r[104] = ld_data_v_r_104_sv2v_reg;
  assign ld_data_v_r[103] = ld_data_v_r_103_sv2v_reg;
  assign ld_data_v_r[102] = ld_data_v_r_102_sv2v_reg;
  assign ld_data_v_r[101] = ld_data_v_r_101_sv2v_reg;
  assign ld_data_v_r[100] = ld_data_v_r_100_sv2v_reg;
  assign ld_data_v_r[99] = ld_data_v_r_99_sv2v_reg;
  assign ld_data_v_r[98] = ld_data_v_r_98_sv2v_reg;
  assign ld_data_v_r[97] = ld_data_v_r_97_sv2v_reg;
  assign ld_data_v_r[96] = ld_data_v_r_96_sv2v_reg;
  assign ld_data_v_r[95] = ld_data_v_r_95_sv2v_reg;
  assign ld_data_v_r[94] = ld_data_v_r_94_sv2v_reg;
  assign ld_data_v_r[93] = ld_data_v_r_93_sv2v_reg;
  assign ld_data_v_r[92] = ld_data_v_r_92_sv2v_reg;
  assign ld_data_v_r[91] = ld_data_v_r_91_sv2v_reg;
  assign ld_data_v_r[90] = ld_data_v_r_90_sv2v_reg;
  assign ld_data_v_r[89] = ld_data_v_r_89_sv2v_reg;
  assign ld_data_v_r[88] = ld_data_v_r_88_sv2v_reg;
  assign ld_data_v_r[87] = ld_data_v_r_87_sv2v_reg;
  assign ld_data_v_r[86] = ld_data_v_r_86_sv2v_reg;
  assign ld_data_v_r[85] = ld_data_v_r_85_sv2v_reg;
  assign ld_data_v_r[84] = ld_data_v_r_84_sv2v_reg;
  assign ld_data_v_r[83] = ld_data_v_r_83_sv2v_reg;
  assign ld_data_v_r[82] = ld_data_v_r_82_sv2v_reg;
  assign ld_data_v_r[81] = ld_data_v_r_81_sv2v_reg;
  assign ld_data_v_r[80] = ld_data_v_r_80_sv2v_reg;
  assign ld_data_v_r[79] = ld_data_v_r_79_sv2v_reg;
  assign ld_data_v_r[78] = ld_data_v_r_78_sv2v_reg;
  assign ld_data_v_r[77] = ld_data_v_r_77_sv2v_reg;
  assign ld_data_v_r[76] = ld_data_v_r_76_sv2v_reg;
  assign ld_data_v_r[75] = ld_data_v_r_75_sv2v_reg;
  assign ld_data_v_r[74] = ld_data_v_r_74_sv2v_reg;
  assign ld_data_v_r[73] = ld_data_v_r_73_sv2v_reg;
  assign ld_data_v_r[72] = ld_data_v_r_72_sv2v_reg;
  assign ld_data_v_r[71] = ld_data_v_r_71_sv2v_reg;
  assign ld_data_v_r[70] = ld_data_v_r_70_sv2v_reg;
  assign ld_data_v_r[69] = ld_data_v_r_69_sv2v_reg;
  assign ld_data_v_r[68] = ld_data_v_r_68_sv2v_reg;
  assign ld_data_v_r[67] = ld_data_v_r_67_sv2v_reg;
  assign ld_data_v_r[66] = ld_data_v_r_66_sv2v_reg;
  assign ld_data_v_r[65] = ld_data_v_r_65_sv2v_reg;
  assign ld_data_v_r[64] = ld_data_v_r_64_sv2v_reg;
  assign ld_data_v_r[63] = ld_data_v_r_63_sv2v_reg;
  assign ld_data_v_r[62] = ld_data_v_r_62_sv2v_reg;
  assign ld_data_v_r[61] = ld_data_v_r_61_sv2v_reg;
  assign ld_data_v_r[60] = ld_data_v_r_60_sv2v_reg;
  assign ld_data_v_r[59] = ld_data_v_r_59_sv2v_reg;
  assign ld_data_v_r[58] = ld_data_v_r_58_sv2v_reg;
  assign ld_data_v_r[57] = ld_data_v_r_57_sv2v_reg;
  assign ld_data_v_r[56] = ld_data_v_r_56_sv2v_reg;
  assign ld_data_v_r[55] = ld_data_v_r_55_sv2v_reg;
  assign ld_data_v_r[54] = ld_data_v_r_54_sv2v_reg;
  assign ld_data_v_r[53] = ld_data_v_r_53_sv2v_reg;
  assign ld_data_v_r[52] = ld_data_v_r_52_sv2v_reg;
  assign ld_data_v_r[51] = ld_data_v_r_51_sv2v_reg;
  assign ld_data_v_r[50] = ld_data_v_r_50_sv2v_reg;
  assign ld_data_v_r[49] = ld_data_v_r_49_sv2v_reg;
  assign ld_data_v_r[48] = ld_data_v_r_48_sv2v_reg;
  assign ld_data_v_r[47] = ld_data_v_r_47_sv2v_reg;
  assign ld_data_v_r[46] = ld_data_v_r_46_sv2v_reg;
  assign ld_data_v_r[45] = ld_data_v_r_45_sv2v_reg;
  assign ld_data_v_r[44] = ld_data_v_r_44_sv2v_reg;
  assign ld_data_v_r[43] = ld_data_v_r_43_sv2v_reg;
  assign ld_data_v_r[42] = ld_data_v_r_42_sv2v_reg;
  assign ld_data_v_r[41] = ld_data_v_r_41_sv2v_reg;
  assign ld_data_v_r[40] = ld_data_v_r_40_sv2v_reg;
  assign ld_data_v_r[39] = ld_data_v_r_39_sv2v_reg;
  assign ld_data_v_r[38] = ld_data_v_r_38_sv2v_reg;
  assign ld_data_v_r[37] = ld_data_v_r_37_sv2v_reg;
  assign ld_data_v_r[36] = ld_data_v_r_36_sv2v_reg;
  assign ld_data_v_r[35] = ld_data_v_r_35_sv2v_reg;
  assign ld_data_v_r[34] = ld_data_v_r_34_sv2v_reg;
  assign ld_data_v_r[33] = ld_data_v_r_33_sv2v_reg;
  assign ld_data_v_r[32] = ld_data_v_r_32_sv2v_reg;
  assign ld_data_v_r[31] = ld_data_v_r_31_sv2v_reg;
  assign ld_data_v_r[30] = ld_data_v_r_30_sv2v_reg;
  assign ld_data_v_r[29] = ld_data_v_r_29_sv2v_reg;
  assign ld_data_v_r[28] = ld_data_v_r_28_sv2v_reg;
  assign ld_data_v_r[27] = ld_data_v_r_27_sv2v_reg;
  assign ld_data_v_r[26] = ld_data_v_r_26_sv2v_reg;
  assign ld_data_v_r[25] = ld_data_v_r_25_sv2v_reg;
  assign ld_data_v_r[24] = ld_data_v_r_24_sv2v_reg;
  assign ld_data_v_r[23] = ld_data_v_r_23_sv2v_reg;
  assign ld_data_v_r[22] = ld_data_v_r_22_sv2v_reg;
  assign ld_data_v_r[21] = ld_data_v_r_21_sv2v_reg;
  assign ld_data_v_r[20] = ld_data_v_r_20_sv2v_reg;
  assign ld_data_v_r[19] = ld_data_v_r_19_sv2v_reg;
  assign ld_data_v_r[18] = ld_data_v_r_18_sv2v_reg;
  assign ld_data_v_r[17] = ld_data_v_r_17_sv2v_reg;
  assign ld_data_v_r[16] = ld_data_v_r_16_sv2v_reg;
  assign ld_data_v_r[15] = ld_data_v_r_15_sv2v_reg;
  assign ld_data_v_r[14] = ld_data_v_r_14_sv2v_reg;
  assign ld_data_v_r[13] = ld_data_v_r_13_sv2v_reg;
  assign ld_data_v_r[12] = ld_data_v_r_12_sv2v_reg;
  assign ld_data_v_r[11] = ld_data_v_r_11_sv2v_reg;
  assign ld_data_v_r[10] = ld_data_v_r_10_sv2v_reg;
  assign ld_data_v_r[9] = ld_data_v_r_9_sv2v_reg;
  assign ld_data_v_r[8] = ld_data_v_r_8_sv2v_reg;
  assign ld_data_v_r[7] = ld_data_v_r_7_sv2v_reg;
  assign ld_data_v_r[6] = ld_data_v_r_6_sv2v_reg;
  assign ld_data_v_r[5] = ld_data_v_r_5_sv2v_reg;
  assign ld_data_v_r[4] = ld_data_v_r_4_sv2v_reg;
  assign ld_data_v_r[3] = ld_data_v_r_3_sv2v_reg;
  assign ld_data_v_r[2] = ld_data_v_r_2_sv2v_reg;
  assign ld_data_v_r[1] = ld_data_v_r_1_sv2v_reg;
  assign ld_data_v_r[0] = ld_data_v_r_0_sv2v_reg;
  assign v_v_r = v_v_r_sv2v_reg;
  assign track_data_v_r[31] = track_data_v_r_31_sv2v_reg;
  assign track_data_v_r[30] = track_data_v_r_30_sv2v_reg;
  assign track_data_v_r[29] = track_data_v_r_29_sv2v_reg;
  assign track_data_v_r[28] = track_data_v_r_28_sv2v_reg;
  assign track_data_v_r[27] = track_data_v_r_27_sv2v_reg;
  assign track_data_v_r[26] = track_data_v_r_26_sv2v_reg;
  assign track_data_v_r[25] = track_data_v_r_25_sv2v_reg;
  assign track_data_v_r[24] = track_data_v_r_24_sv2v_reg;
  assign track_data_v_r[23] = track_data_v_r_23_sv2v_reg;
  assign track_data_v_r[22] = track_data_v_r_22_sv2v_reg;
  assign track_data_v_r[21] = track_data_v_r_21_sv2v_reg;
  assign track_data_v_r[20] = track_data_v_r_20_sv2v_reg;
  assign track_data_v_r[19] = track_data_v_r_19_sv2v_reg;
  assign track_data_v_r[18] = track_data_v_r_18_sv2v_reg;
  assign track_data_v_r[17] = track_data_v_r_17_sv2v_reg;
  assign track_data_v_r[16] = track_data_v_r_16_sv2v_reg;
  assign track_data_v_r[15] = track_data_v_r_15_sv2v_reg;
  assign track_data_v_r[14] = track_data_v_r_14_sv2v_reg;
  assign track_data_v_r[13] = track_data_v_r_13_sv2v_reg;
  assign track_data_v_r[12] = track_data_v_r_12_sv2v_reg;
  assign track_data_v_r[11] = track_data_v_r_11_sv2v_reg;
  assign track_data_v_r[10] = track_data_v_r_10_sv2v_reg;
  assign track_data_v_r[9] = track_data_v_r_9_sv2v_reg;
  assign track_data_v_r[8] = track_data_v_r_8_sv2v_reg;
  assign track_data_v_r[7] = track_data_v_r_7_sv2v_reg;
  assign track_data_v_r[6] = track_data_v_r_6_sv2v_reg;
  assign track_data_v_r[5] = track_data_v_r_5_sv2v_reg;
  assign track_data_v_r[4] = track_data_v_r_4_sv2v_reg;
  assign track_data_v_r[3] = track_data_v_r_3_sv2v_reg;
  assign track_data_v_r[2] = track_data_v_r_2_sv2v_reg;
  assign track_data_v_r[1] = track_data_v_r_1_sv2v_reg;
  assign track_data_v_r[0] = track_data_v_r_0_sv2v_reg;
  assign mask_v_r[15] = mask_v_r_15_sv2v_reg;
  assign mask_v_r[14] = mask_v_r_14_sv2v_reg;
  assign mask_v_r[13] = mask_v_r_13_sv2v_reg;
  assign mask_v_r[12] = mask_v_r_12_sv2v_reg;
  assign mask_v_r[11] = mask_v_r_11_sv2v_reg;
  assign mask_v_r[10] = mask_v_r_10_sv2v_reg;
  assign mask_v_r[9] = mask_v_r_9_sv2v_reg;
  assign mask_v_r[8] = mask_v_r_8_sv2v_reg;
  assign mask_v_r[7] = mask_v_r_7_sv2v_reg;
  assign mask_v_r[6] = mask_v_r_6_sv2v_reg;
  assign mask_v_r[5] = mask_v_r_5_sv2v_reg;
  assign mask_v_r[4] = mask_v_r_4_sv2v_reg;
  assign mask_v_r[3] = mask_v_r_3_sv2v_reg;
  assign mask_v_r[2] = mask_v_r_2_sv2v_reg;
  assign mask_v_r[1] = mask_v_r_1_sv2v_reg;
  assign mask_v_r[0] = mask_v_r_0_sv2v_reg;
  assign decode_v_r[20] = decode_v_r_20_sv2v_reg;
  assign decode_v_r[19] = decode_v_r_19_sv2v_reg;
  assign decode_v_r[18] = decode_v_r_18_sv2v_reg;
  assign decode_v_r[17] = decode_v_r_17_sv2v_reg;
  assign decode_v_r[16] = decode_v_r_16_sv2v_reg;
  assign decode_v_r[15] = decode_v_r_15_sv2v_reg;
  assign decode_v_r[14] = decode_v_r_14_sv2v_reg;
  assign decode_v_r[13] = decode_v_r_13_sv2v_reg;
  assign decode_v_r[12] = decode_v_r_12_sv2v_reg;
  assign decode_v_r[11] = decode_v_r_11_sv2v_reg;
  assign decode_v_r[10] = decode_v_r_10_sv2v_reg;
  assign decode_v_r[9] = decode_v_r_9_sv2v_reg;
  assign decode_v_r[8] = decode_v_r_8_sv2v_reg;
  assign decode_v_r[7] = decode_v_r_7_sv2v_reg;
  assign decode_v_r[6] = decode_v_r_6_sv2v_reg;
  assign decode_v_r[5] = decode_v_r_5_sv2v_reg;
  assign decode_v_r[4] = decode_v_r_4_sv2v_reg;
  assign decode_v_r[3] = decode_v_r_3_sv2v_reg;
  assign decode_v_r[2] = decode_v_r_2_sv2v_reg;
  assign decode_v_r[1] = decode_v_r_1_sv2v_reg;
  assign decode_v_r[0] = decode_v_r_0_sv2v_reg;
  assign addr_v_r[32] = addr_v_r_32_sv2v_reg;
  assign addr_v_r[31] = addr_v_r_31_sv2v_reg;
  assign addr_v_r[30] = addr_v_r_30_sv2v_reg;
  assign addr_v_r[29] = addr_v_r_29_sv2v_reg;
  assign addr_v_r[28] = addr_v_r_28_sv2v_reg;
  assign addr_v_r[27] = addr_v_r_27_sv2v_reg;
  assign addr_v_r[26] = addr_v_r_26_sv2v_reg;
  assign addr_v_r[25] = addr_v_r_25_sv2v_reg;
  assign addr_v_r[24] = addr_v_r_24_sv2v_reg;
  assign addr_v_r[23] = addr_v_r_23_sv2v_reg;
  assign addr_v_r[22] = addr_v_r_22_sv2v_reg;
  assign addr_v_r[21] = addr_v_r_21_sv2v_reg;
  assign addr_v_r[20] = addr_v_r_20_sv2v_reg;
  assign addr_v_r[19] = addr_v_r_19_sv2v_reg;
  assign addr_v_r[18] = addr_v_r_18_sv2v_reg;
  assign addr_v_r[17] = addr_v_r_17_sv2v_reg;
  assign addr_v_r[16] = addr_v_r_16_sv2v_reg;
  assign addr_v_r[15] = addr_v_r_15_sv2v_reg;
  assign addr_v_r[14] = addr_v_r_14_sv2v_reg;
  assign addr_v_r[13] = addr_v_r_13_sv2v_reg;
  assign addr_v_r[12] = addr_v_r_12_sv2v_reg;
  assign addr_v_r[11] = addr_v_r_11_sv2v_reg;
  assign addr_v_r[10] = addr_v_r_10_sv2v_reg;
  assign addr_v_r[9] = addr_v_r_9_sv2v_reg;
  assign addr_v_r[8] = addr_v_r_8_sv2v_reg;
  assign addr_v_r[7] = addr_v_r_7_sv2v_reg;
  assign addr_v_r[6] = addr_v_r_6_sv2v_reg;
  assign addr_v_r[5] = addr_v_r_5_sv2v_reg;
  assign addr_v_r[4] = addr_v_r_4_sv2v_reg;
  assign addr_v_r[3] = addr_v_r_3_sv2v_reg;
  assign addr_v_r[2] = addr_v_r_2_sv2v_reg;
  assign addr_v_r[1] = addr_v_r_1_sv2v_reg;
  assign addr_v_r[0] = addr_v_r_0_sv2v_reg;
  assign data_v_r[127] = data_v_r_127_sv2v_reg;
  assign data_v_r[126] = data_v_r_126_sv2v_reg;
  assign data_v_r[125] = data_v_r_125_sv2v_reg;
  assign data_v_r[124] = data_v_r_124_sv2v_reg;
  assign data_v_r[123] = data_v_r_123_sv2v_reg;
  assign data_v_r[122] = data_v_r_122_sv2v_reg;
  assign data_v_r[121] = data_v_r_121_sv2v_reg;
  assign data_v_r[120] = data_v_r_120_sv2v_reg;
  assign data_v_r[119] = data_v_r_119_sv2v_reg;
  assign data_v_r[118] = data_v_r_118_sv2v_reg;
  assign data_v_r[117] = data_v_r_117_sv2v_reg;
  assign data_v_r[116] = data_v_r_116_sv2v_reg;
  assign data_v_r[115] = data_v_r_115_sv2v_reg;
  assign data_v_r[114] = data_v_r_114_sv2v_reg;
  assign data_v_r[113] = data_v_r_113_sv2v_reg;
  assign data_v_r[112] = data_v_r_112_sv2v_reg;
  assign data_v_r[111] = data_v_r_111_sv2v_reg;
  assign data_v_r[110] = data_v_r_110_sv2v_reg;
  assign data_v_r[109] = data_v_r_109_sv2v_reg;
  assign data_v_r[108] = data_v_r_108_sv2v_reg;
  assign data_v_r[107] = data_v_r_107_sv2v_reg;
  assign data_v_r[106] = data_v_r_106_sv2v_reg;
  assign data_v_r[105] = data_v_r_105_sv2v_reg;
  assign data_v_r[104] = data_v_r_104_sv2v_reg;
  assign data_v_r[103] = data_v_r_103_sv2v_reg;
  assign data_v_r[102] = data_v_r_102_sv2v_reg;
  assign data_v_r[101] = data_v_r_101_sv2v_reg;
  assign data_v_r[100] = data_v_r_100_sv2v_reg;
  assign data_v_r[99] = data_v_r_99_sv2v_reg;
  assign data_v_r[98] = data_v_r_98_sv2v_reg;
  assign data_v_r[97] = data_v_r_97_sv2v_reg;
  assign data_v_r[96] = data_v_r_96_sv2v_reg;
  assign data_v_r[95] = data_v_r_95_sv2v_reg;
  assign data_v_r[94] = data_v_r_94_sv2v_reg;
  assign data_v_r[93] = data_v_r_93_sv2v_reg;
  assign data_v_r[92] = data_v_r_92_sv2v_reg;
  assign data_v_r[91] = data_v_r_91_sv2v_reg;
  assign data_v_r[90] = data_v_r_90_sv2v_reg;
  assign data_v_r[89] = data_v_r_89_sv2v_reg;
  assign data_v_r[88] = data_v_r_88_sv2v_reg;
  assign data_v_r[87] = data_v_r_87_sv2v_reg;
  assign data_v_r[86] = data_v_r_86_sv2v_reg;
  assign data_v_r[85] = data_v_r_85_sv2v_reg;
  assign data_v_r[84] = data_v_r_84_sv2v_reg;
  assign data_v_r[83] = data_v_r_83_sv2v_reg;
  assign data_v_r[82] = data_v_r_82_sv2v_reg;
  assign data_v_r[81] = data_v_r_81_sv2v_reg;
  assign data_v_r[80] = data_v_r_80_sv2v_reg;
  assign data_v_r[79] = data_v_r_79_sv2v_reg;
  assign data_v_r[78] = data_v_r_78_sv2v_reg;
  assign data_v_r[77] = data_v_r_77_sv2v_reg;
  assign data_v_r[76] = data_v_r_76_sv2v_reg;
  assign data_v_r[75] = data_v_r_75_sv2v_reg;
  assign data_v_r[74] = data_v_r_74_sv2v_reg;
  assign data_v_r[73] = data_v_r_73_sv2v_reg;
  assign data_v_r[72] = data_v_r_72_sv2v_reg;
  assign data_v_r[71] = data_v_r_71_sv2v_reg;
  assign data_v_r[70] = data_v_r_70_sv2v_reg;
  assign data_v_r[69] = data_v_r_69_sv2v_reg;
  assign data_v_r[68] = data_v_r_68_sv2v_reg;
  assign data_v_r[67] = data_v_r_67_sv2v_reg;
  assign data_v_r[66] = data_v_r_66_sv2v_reg;
  assign data_v_r[65] = data_v_r_65_sv2v_reg;
  assign data_v_r[64] = data_v_r_64_sv2v_reg;
  assign data_v_r[63] = data_v_r_63_sv2v_reg;
  assign data_v_r[62] = data_v_r_62_sv2v_reg;
  assign data_v_r[61] = data_v_r_61_sv2v_reg;
  assign data_v_r[60] = data_v_r_60_sv2v_reg;
  assign data_v_r[59] = data_v_r_59_sv2v_reg;
  assign data_v_r[58] = data_v_r_58_sv2v_reg;
  assign data_v_r[57] = data_v_r_57_sv2v_reg;
  assign data_v_r[56] = data_v_r_56_sv2v_reg;
  assign data_v_r[55] = data_v_r_55_sv2v_reg;
  assign data_v_r[54] = data_v_r_54_sv2v_reg;
  assign data_v_r[53] = data_v_r_53_sv2v_reg;
  assign data_v_r[52] = data_v_r_52_sv2v_reg;
  assign data_v_r[51] = data_v_r_51_sv2v_reg;
  assign data_v_r[50] = data_v_r_50_sv2v_reg;
  assign data_v_r[49] = data_v_r_49_sv2v_reg;
  assign data_v_r[48] = data_v_r_48_sv2v_reg;
  assign data_v_r[47] = data_v_r_47_sv2v_reg;
  assign data_v_r[46] = data_v_r_46_sv2v_reg;
  assign data_v_r[45] = data_v_r_45_sv2v_reg;
  assign data_v_r[44] = data_v_r_44_sv2v_reg;
  assign data_v_r[43] = data_v_r_43_sv2v_reg;
  assign data_v_r[42] = data_v_r_42_sv2v_reg;
  assign data_v_r[41] = data_v_r_41_sv2v_reg;
  assign data_v_r[40] = data_v_r_40_sv2v_reg;
  assign data_v_r[39] = data_v_r_39_sv2v_reg;
  assign data_v_r[38] = data_v_r_38_sv2v_reg;
  assign data_v_r[37] = data_v_r_37_sv2v_reg;
  assign data_v_r[36] = data_v_r_36_sv2v_reg;
  assign data_v_r[35] = data_v_r_35_sv2v_reg;
  assign data_v_r[34] = data_v_r_34_sv2v_reg;
  assign data_v_r[33] = data_v_r_33_sv2v_reg;
  assign data_v_r[32] = data_v_r_32_sv2v_reg;
  assign data_v_r[31] = data_v_r_31_sv2v_reg;
  assign data_v_r[30] = data_v_r_30_sv2v_reg;
  assign data_v_r[29] = data_v_r_29_sv2v_reg;
  assign data_v_r[28] = data_v_r_28_sv2v_reg;
  assign data_v_r[27] = data_v_r_27_sv2v_reg;
  assign data_v_r[26] = data_v_r_26_sv2v_reg;
  assign data_v_r[25] = data_v_r_25_sv2v_reg;
  assign data_v_r[24] = data_v_r_24_sv2v_reg;
  assign data_v_r[23] = data_v_r_23_sv2v_reg;
  assign data_v_r[22] = data_v_r_22_sv2v_reg;
  assign data_v_r[21] = data_v_r_21_sv2v_reg;
  assign data_v_r[20] = data_v_r_20_sv2v_reg;
  assign data_v_r[19] = data_v_r_19_sv2v_reg;
  assign data_v_r[18] = data_v_r_18_sv2v_reg;
  assign data_v_r[17] = data_v_r_17_sv2v_reg;
  assign data_v_r[16] = data_v_r_16_sv2v_reg;
  assign data_v_r[15] = data_v_r_15_sv2v_reg;
  assign data_v_r[14] = data_v_r_14_sv2v_reg;
  assign data_v_r[13] = data_v_r_13_sv2v_reg;
  assign data_v_r[12] = data_v_r_12_sv2v_reg;
  assign data_v_r[11] = data_v_r_11_sv2v_reg;
  assign data_v_r[10] = data_v_r_10_sv2v_reg;
  assign data_v_r[9] = data_v_r_9_sv2v_reg;
  assign data_v_r[8] = data_v_r_8_sv2v_reg;
  assign data_v_r[7] = data_v_r_7_sv2v_reg;
  assign data_v_r[6] = data_v_r_6_sv2v_reg;
  assign data_v_r[5] = data_v_r_5_sv2v_reg;
  assign data_v_r[4] = data_v_r_4_sv2v_reg;
  assign data_v_r[3] = data_v_r_3_sv2v_reg;
  assign data_v_r[2] = data_v_r_2_sv2v_reg;
  assign data_v_r[1] = data_v_r_1_sv2v_reg;
  assign data_v_r[0] = data_v_r_0_sv2v_reg;
  assign valid_v_r[7] = valid_v_r_7_sv2v_reg;
  assign valid_v_r[6] = valid_v_r_6_sv2v_reg;
  assign valid_v_r[5] = valid_v_r_5_sv2v_reg;
  assign valid_v_r[4] = valid_v_r_4_sv2v_reg;
  assign valid_v_r[3] = valid_v_r_3_sv2v_reg;
  assign valid_v_r[2] = valid_v_r_2_sv2v_reg;
  assign valid_v_r[1] = valid_v_r_1_sv2v_reg;
  assign valid_v_r[0] = valid_v_r_0_sv2v_reg;
  assign lock_v_r[7] = lock_v_r_7_sv2v_reg;
  assign lock_v_r[6] = lock_v_r_6_sv2v_reg;
  assign lock_v_r[5] = lock_v_r_5_sv2v_reg;
  assign lock_v_r[4] = lock_v_r_4_sv2v_reg;
  assign lock_v_r[3] = lock_v_r_3_sv2v_reg;
  assign lock_v_r[2] = lock_v_r_2_sv2v_reg;
  assign lock_v_r[1] = lock_v_r_1_sv2v_reg;
  assign lock_v_r[0] = lock_v_r_0_sv2v_reg;
  assign tag_v_r[159] = tag_v_r_159_sv2v_reg;
  assign tag_v_r[158] = tag_v_r_158_sv2v_reg;
  assign tag_v_r[157] = tag_v_r_157_sv2v_reg;
  assign tag_v_r[156] = tag_v_r_156_sv2v_reg;
  assign tag_v_r[155] = tag_v_r_155_sv2v_reg;
  assign tag_v_r[154] = tag_v_r_154_sv2v_reg;
  assign tag_v_r[153] = tag_v_r_153_sv2v_reg;
  assign tag_v_r[152] = tag_v_r_152_sv2v_reg;
  assign tag_v_r[151] = tag_v_r_151_sv2v_reg;
  assign tag_v_r[150] = tag_v_r_150_sv2v_reg;
  assign tag_v_r[149] = tag_v_r_149_sv2v_reg;
  assign tag_v_r[148] = tag_v_r_148_sv2v_reg;
  assign tag_v_r[147] = tag_v_r_147_sv2v_reg;
  assign tag_v_r[146] = tag_v_r_146_sv2v_reg;
  assign tag_v_r[145] = tag_v_r_145_sv2v_reg;
  assign tag_v_r[144] = tag_v_r_144_sv2v_reg;
  assign tag_v_r[143] = tag_v_r_143_sv2v_reg;
  assign tag_v_r[142] = tag_v_r_142_sv2v_reg;
  assign tag_v_r[141] = tag_v_r_141_sv2v_reg;
  assign tag_v_r[140] = tag_v_r_140_sv2v_reg;
  assign tag_v_r[139] = tag_v_r_139_sv2v_reg;
  assign tag_v_r[138] = tag_v_r_138_sv2v_reg;
  assign tag_v_r[137] = tag_v_r_137_sv2v_reg;
  assign tag_v_r[136] = tag_v_r_136_sv2v_reg;
  assign tag_v_r[135] = tag_v_r_135_sv2v_reg;
  assign tag_v_r[134] = tag_v_r_134_sv2v_reg;
  assign tag_v_r[133] = tag_v_r_133_sv2v_reg;
  assign tag_v_r[132] = tag_v_r_132_sv2v_reg;
  assign tag_v_r[131] = tag_v_r_131_sv2v_reg;
  assign tag_v_r[130] = tag_v_r_130_sv2v_reg;
  assign tag_v_r[129] = tag_v_r_129_sv2v_reg;
  assign tag_v_r[128] = tag_v_r_128_sv2v_reg;
  assign tag_v_r[127] = tag_v_r_127_sv2v_reg;
  assign tag_v_r[126] = tag_v_r_126_sv2v_reg;
  assign tag_v_r[125] = tag_v_r_125_sv2v_reg;
  assign tag_v_r[124] = tag_v_r_124_sv2v_reg;
  assign tag_v_r[123] = tag_v_r_123_sv2v_reg;
  assign tag_v_r[122] = tag_v_r_122_sv2v_reg;
  assign tag_v_r[121] = tag_v_r_121_sv2v_reg;
  assign tag_v_r[120] = tag_v_r_120_sv2v_reg;
  assign tag_v_r[119] = tag_v_r_119_sv2v_reg;
  assign tag_v_r[118] = tag_v_r_118_sv2v_reg;
  assign tag_v_r[117] = tag_v_r_117_sv2v_reg;
  assign tag_v_r[116] = tag_v_r_116_sv2v_reg;
  assign tag_v_r[115] = tag_v_r_115_sv2v_reg;
  assign tag_v_r[114] = tag_v_r_114_sv2v_reg;
  assign tag_v_r[113] = tag_v_r_113_sv2v_reg;
  assign tag_v_r[112] = tag_v_r_112_sv2v_reg;
  assign tag_v_r[111] = tag_v_r_111_sv2v_reg;
  assign tag_v_r[110] = tag_v_r_110_sv2v_reg;
  assign tag_v_r[109] = tag_v_r_109_sv2v_reg;
  assign tag_v_r[108] = tag_v_r_108_sv2v_reg;
  assign tag_v_r[107] = tag_v_r_107_sv2v_reg;
  assign tag_v_r[106] = tag_v_r_106_sv2v_reg;
  assign tag_v_r[105] = tag_v_r_105_sv2v_reg;
  assign tag_v_r[104] = tag_v_r_104_sv2v_reg;
  assign tag_v_r[103] = tag_v_r_103_sv2v_reg;
  assign tag_v_r[102] = tag_v_r_102_sv2v_reg;
  assign tag_v_r[101] = tag_v_r_101_sv2v_reg;
  assign tag_v_r[100] = tag_v_r_100_sv2v_reg;
  assign tag_v_r[99] = tag_v_r_99_sv2v_reg;
  assign tag_v_r[98] = tag_v_r_98_sv2v_reg;
  assign tag_v_r[97] = tag_v_r_97_sv2v_reg;
  assign tag_v_r[96] = tag_v_r_96_sv2v_reg;
  assign tag_v_r[95] = tag_v_r_95_sv2v_reg;
  assign tag_v_r[94] = tag_v_r_94_sv2v_reg;
  assign tag_v_r[93] = tag_v_r_93_sv2v_reg;
  assign tag_v_r[92] = tag_v_r_92_sv2v_reg;
  assign tag_v_r[91] = tag_v_r_91_sv2v_reg;
  assign tag_v_r[90] = tag_v_r_90_sv2v_reg;
  assign tag_v_r[89] = tag_v_r_89_sv2v_reg;
  assign tag_v_r[88] = tag_v_r_88_sv2v_reg;
  assign tag_v_r[87] = tag_v_r_87_sv2v_reg;
  assign tag_v_r[86] = tag_v_r_86_sv2v_reg;
  assign tag_v_r[85] = tag_v_r_85_sv2v_reg;
  assign tag_v_r[84] = tag_v_r_84_sv2v_reg;
  assign tag_v_r[83] = tag_v_r_83_sv2v_reg;
  assign tag_v_r[82] = tag_v_r_82_sv2v_reg;
  assign tag_v_r[81] = tag_v_r_81_sv2v_reg;
  assign tag_v_r[80] = tag_v_r_80_sv2v_reg;
  assign tag_v_r[79] = tag_v_r_79_sv2v_reg;
  assign tag_v_r[78] = tag_v_r_78_sv2v_reg;
  assign tag_v_r[77] = tag_v_r_77_sv2v_reg;
  assign tag_v_r[76] = tag_v_r_76_sv2v_reg;
  assign tag_v_r[75] = tag_v_r_75_sv2v_reg;
  assign tag_v_r[74] = tag_v_r_74_sv2v_reg;
  assign tag_v_r[73] = tag_v_r_73_sv2v_reg;
  assign tag_v_r[72] = tag_v_r_72_sv2v_reg;
  assign tag_v_r[71] = tag_v_r_71_sv2v_reg;
  assign tag_v_r[70] = tag_v_r_70_sv2v_reg;
  assign tag_v_r[69] = tag_v_r_69_sv2v_reg;
  assign tag_v_r[68] = tag_v_r_68_sv2v_reg;
  assign tag_v_r[67] = tag_v_r_67_sv2v_reg;
  assign tag_v_r[66] = tag_v_r_66_sv2v_reg;
  assign tag_v_r[65] = tag_v_r_65_sv2v_reg;
  assign tag_v_r[64] = tag_v_r_64_sv2v_reg;
  assign tag_v_r[63] = tag_v_r_63_sv2v_reg;
  assign tag_v_r[62] = tag_v_r_62_sv2v_reg;
  assign tag_v_r[61] = tag_v_r_61_sv2v_reg;
  assign tag_v_r[60] = tag_v_r_60_sv2v_reg;
  assign tag_v_r[59] = tag_v_r_59_sv2v_reg;
  assign tag_v_r[58] = tag_v_r_58_sv2v_reg;
  assign tag_v_r[57] = tag_v_r_57_sv2v_reg;
  assign tag_v_r[56] = tag_v_r_56_sv2v_reg;
  assign tag_v_r[55] = tag_v_r_55_sv2v_reg;
  assign tag_v_r[54] = tag_v_r_54_sv2v_reg;
  assign tag_v_r[53] = tag_v_r_53_sv2v_reg;
  assign tag_v_r[52] = tag_v_r_52_sv2v_reg;
  assign tag_v_r[51] = tag_v_r_51_sv2v_reg;
  assign tag_v_r[50] = tag_v_r_50_sv2v_reg;
  assign tag_v_r[49] = tag_v_r_49_sv2v_reg;
  assign tag_v_r[48] = tag_v_r_48_sv2v_reg;
  assign tag_v_r[47] = tag_v_r_47_sv2v_reg;
  assign tag_v_r[46] = tag_v_r_46_sv2v_reg;
  assign tag_v_r[45] = tag_v_r_45_sv2v_reg;
  assign tag_v_r[44] = tag_v_r_44_sv2v_reg;
  assign tag_v_r[43] = tag_v_r_43_sv2v_reg;
  assign tag_v_r[42] = tag_v_r_42_sv2v_reg;
  assign tag_v_r[41] = tag_v_r_41_sv2v_reg;
  assign tag_v_r[40] = tag_v_r_40_sv2v_reg;
  assign tag_v_r[39] = tag_v_r_39_sv2v_reg;
  assign tag_v_r[38] = tag_v_r_38_sv2v_reg;
  assign tag_v_r[37] = tag_v_r_37_sv2v_reg;
  assign tag_v_r[36] = tag_v_r_36_sv2v_reg;
  assign tag_v_r[35] = tag_v_r_35_sv2v_reg;
  assign tag_v_r[34] = tag_v_r_34_sv2v_reg;
  assign tag_v_r[33] = tag_v_r_33_sv2v_reg;
  assign tag_v_r[32] = tag_v_r_32_sv2v_reg;
  assign tag_v_r[31] = tag_v_r_31_sv2v_reg;
  assign tag_v_r[30] = tag_v_r_30_sv2v_reg;
  assign tag_v_r[29] = tag_v_r_29_sv2v_reg;
  assign tag_v_r[28] = tag_v_r_28_sv2v_reg;
  assign tag_v_r[27] = tag_v_r_27_sv2v_reg;
  assign tag_v_r[26] = tag_v_r_26_sv2v_reg;
  assign tag_v_r[25] = tag_v_r_25_sv2v_reg;
  assign tag_v_r[24] = tag_v_r_24_sv2v_reg;
  assign tag_v_r[23] = tag_v_r_23_sv2v_reg;
  assign tag_v_r[22] = tag_v_r_22_sv2v_reg;
  assign tag_v_r[21] = tag_v_r_21_sv2v_reg;
  assign tag_v_r[20] = tag_v_r_20_sv2v_reg;
  assign tag_v_r[19] = tag_v_r_19_sv2v_reg;
  assign tag_v_r[18] = tag_v_r_18_sv2v_reg;
  assign tag_v_r[17] = tag_v_r_17_sv2v_reg;
  assign tag_v_r[16] = tag_v_r_16_sv2v_reg;
  assign tag_v_r[15] = tag_v_r_15_sv2v_reg;
  assign tag_v_r[14] = tag_v_r_14_sv2v_reg;
  assign tag_v_r[13] = tag_v_r_13_sv2v_reg;
  assign tag_v_r[12] = tag_v_r_12_sv2v_reg;
  assign tag_v_r[11] = tag_v_r_11_sv2v_reg;
  assign tag_v_r[10] = tag_v_r_10_sv2v_reg;
  assign tag_v_r[9] = tag_v_r_9_sv2v_reg;
  assign tag_v_r[8] = tag_v_r_8_sv2v_reg;
  assign tag_v_r[7] = tag_v_r_7_sv2v_reg;
  assign tag_v_r[6] = tag_v_r_6_sv2v_reg;
  assign tag_v_r[5] = tag_v_r_5_sv2v_reg;
  assign tag_v_r[4] = tag_v_r_4_sv2v_reg;
  assign tag_v_r[3] = tag_v_r_3_sv2v_reg;
  assign tag_v_r[2] = tag_v_r_2_sv2v_reg;
  assign tag_v_r[1] = tag_v_r_1_sv2v_reg;
  assign tag_v_r[0] = tag_v_r_0_sv2v_reg;

  bsg_cache_decode
  decode0
  (
    .opcode_i(cache_pkt_i[182:177]),
    .decode_o(decode)
  );


  bsg_mem_1rw_sync_mask_write_bit_000000b0_00000080_1
  tag_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(tag_mem_data_li),
    .addr_i(tag_mem_addr_li),
    .v_i(tag_mem_v_li),
    .w_mask_i(tag_mem_w_mask_li),
    .w_i(tag_mem_w_li),
    .data_o(tag_mem_data_lo)
  );


  bsg_mem_1rw_sync_mask_write_byte_00000200_00000400_1
  data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li),
    .data_i(data_mem_data_li),
    .write_mask_i(data_mem_w_mask_li),
    .data_o(data_mem_data_lo)
  );


  bsg_mem_1rw_sync_mask_write_bit_00000020_00000080_1
  \track_mem_gen.track_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(track_mem_data_li),
    .addr_i(track_mem_addr_li),
    .v_i(track_mem_v_li),
    .w_mask_i(track_mem_w_mask_li),
    .w_i(track_mem_w_li),
    .data_o(track_mem_data_lo)
  );

  assign N117 = addr_v_r[32:13] == tag_v_r[19:0];
  assign N118 = addr_v_r[32:13] == tag_v_r[39:20];
  assign N119 = addr_v_r[32:13] == tag_v_r[59:40];
  assign N120 = addr_v_r[32:13] == tag_v_r[79:60];
  assign N121 = addr_v_r[32:13] == tag_v_r[99:80];
  assign N122 = addr_v_r[32:13] == tag_v_r[119:100];
  assign N123 = addr_v_r[32:13] == tag_v_r[139:120];
  assign N124 = addr_v_r[32:13] == tag_v_r[159:140];

  bsg_priority_encode_00000008_1
  tag_hit_pe
  (
    .i(tag_hit_v),
    .addr_o(tag_hit_way_id),
    .v_o(tag_hit_found)
  );

  assign N150 = (N142)? track_data_v_r[3] : 
                (N144)? track_data_v_r[7] : 
                (N146)? track_data_v_r[11] : 
                (N148)? track_data_v_r[15] : 
                (N143)? track_data_v_r[19] : 
                (N145)? track_data_v_r[23] : 
                (N147)? track_data_v_r[27] : 
                (N149)? track_data_v_r[31] : 1'b0;
  assign N151 = (N142)? track_data_v_r[2] : 
                (N144)? track_data_v_r[6] : 
                (N146)? track_data_v_r[10] : 
                (N148)? track_data_v_r[14] : 
                (N143)? track_data_v_r[18] : 
                (N145)? track_data_v_r[22] : 
                (N147)? track_data_v_r[26] : 
                (N149)? track_data_v_r[30] : 1'b0;
  assign N152 = (N142)? track_data_v_r[1] : 
                (N144)? track_data_v_r[5] : 
                (N146)? track_data_v_r[9] : 
                (N148)? track_data_v_r[13] : 
                (N143)? track_data_v_r[17] : 
                (N145)? track_data_v_r[21] : 
                (N147)? track_data_v_r[25] : 
                (N149)? track_data_v_r[29] : 1'b0;
  assign N153 = (N142)? track_data_v_r[0] : 
                (N144)? track_data_v_r[4] : 
                (N146)? track_data_v_r[8] : 
                (N148)? track_data_v_r[12] : 
                (N143)? track_data_v_r[16] : 
                (N145)? track_data_v_r[20] : 
                (N147)? track_data_v_r[24] : 
                (N149)? track_data_v_r[28] : 1'b0;
  assign N160 = (N156)? N153 : 
                (N158)? N152 : 
                (N157)? N151 : 
                (N159)? N150 : 1'b0;
  assign N176 = (N168)? valid_v_r[0] : 
                (N170)? valid_v_r[1] : 
                (N172)? valid_v_r[2] : 
                (N174)? valid_v_r[3] : 
                (N169)? valid_v_r[4] : 
                (N171)? valid_v_r[5] : 
                (N173)? valid_v_r[6] : 
                (N175)? valid_v_r[7] : 1'b0;
  assign N194 = (N186)? lock_v_r[0] : 
                (N188)? lock_v_r[1] : 
                (N190)? lock_v_r[2] : 
                (N192)? lock_v_r[3] : 
                (N187)? lock_v_r[4] : 
                (N189)? lock_v_r[5] : 
                (N191)? lock_v_r[6] : 
                (N193)? lock_v_r[7] : 1'b0;
  assign N214 = (N206)? lock_v_r[0] : 
                (N208)? lock_v_r[1] : 
                (N210)? lock_v_r[2] : 
                (N212)? lock_v_r[3] : 
                (N207)? lock_v_r[4] : 
                (N209)? lock_v_r[5] : 
                (N211)? lock_v_r[6] : 
                (N213)? lock_v_r[7] : 1'b0;

  bsg_mem_1rw_sync_mask_write_bit_0000000f_00000080_1
  stat_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(stat_mem_data_li),
    .addr_i(stat_mem_addr_li),
    .v_i(stat_mem_v_li),
    .w_mask_i(stat_mem_w_mask_li),
    .w_i(stat_mem_w_li),
    .data_o(stat_mem_data_lo)
  );


  bsg_cache_miss_00000021_00000080_00000004_00000080_00000008_1
  miss
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .miss_v_i(miss_v),
    .track_miss_i(track_miss),
    .decode_v_i(decode_v_r),
    .addr_v_i(addr_v_r),
    .mask_v_i(mask_v_r),
    .tag_v_i(tag_v_r),
    .valid_v_i(valid_v_r),
    .lock_v_i(lock_v_r),
    .tag_hit_v_i(tag_hit_v),
    .tag_hit_way_id_i(tag_hit_way_id),
    .tag_hit_found_i(tag_hit_found),
    .sbuf_empty_i(sbuf_empty_lo),
    .tbuf_empty_i(tbuf_empty_lo),
    .dma_cmd_o(dma_cmd_lo),
    .dma_way_o(dma_way_lo),
    .dma_addr_o(dma_addr_lo),
    .dma_done_i(dma_done_li),
    .track_data_we_o(miss_track_data_we_lo),
    .stat_info_i(stat_mem_data_lo),
    .stat_mem_v_o(miss_stat_mem_v_lo),
    .stat_mem_w_o(miss_stat_mem_w_lo),
    .stat_mem_addr_o(miss_stat_mem_addr_lo),
    .stat_mem_data_o(miss_stat_mem_data_lo),
    .stat_mem_w_mask_o(miss_stat_mem_w_mask_lo),
    .tag_mem_v_o(miss_tag_mem_v_lo),
    .tag_mem_w_o(miss_tag_mem_w_lo),
    .tag_mem_addr_o(miss_tag_mem_addr_lo),
    .tag_mem_data_o(miss_tag_mem_data_lo),
    .tag_mem_w_mask_o(miss_tag_mem_w_mask_lo),
    .track_mem_v_o(miss_track_mem_v_lo),
    .track_mem_w_o(miss_track_mem_w_lo),
    .track_mem_addr_o(miss_track_mem_addr_lo),
    .track_mem_w_mask_o(miss_track_mem_w_mask_lo),
    .track_mem_data_o(miss_track_mem_data_lo),
    .done_o(miss_done_lo),
    .recover_o(recover_lo),
    .chosen_way_o(chosen_way_lo),
    .select_snoop_data_r_o(select_snoop_data_r_lo),
    .ack_i(_1_net_)
  );


  bsg_cache_dma_00000021_00000080_00000004_00000080_00000008_1_00000080_0
  dma
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .dma_cmd_i(dma_cmd_lo),
    .dma_way_i(dma_way_lo),
    .dma_addr_i(dma_addr_lo),
    .done_o(dma_done_li),
    .track_data_we_i(miss_track_data_we_lo),
    .snoop_word_o(snoop_word_lo),
    .dma_pkt_o(dma_pkt_o),
    .dma_pkt_v_o(dma_pkt_v_o),
    .dma_pkt_yumi_i(dma_pkt_yumi_i),
    .dma_data_i(dma_data_i),
    .dma_data_v_i(dma_data_v_i),
    .dma_data_ready_and_o(dma_data_ready_and_o),
    .dma_data_o(dma_data_o),
    .dma_data_v_o(dma_data_v_o),
    .dma_data_yumi_i(dma_data_yumi_i),
    .data_mem_v_o(dma_data_mem_v_lo),
    .data_mem_w_o(dma_data_mem_w_lo),
    .data_mem_addr_o(dma_data_mem_addr_lo),
    .data_mem_w_mask_o(dma_data_mem_w_mask_lo),
    .data_mem_data_o(dma_data_mem_data_lo),
    .data_mem_data_i(data_mem_data_lo),
    .track_miss_i(track_miss),
    .track_mem_data_i(track_mem_data_lo),
    .dma_evict_o(dma_evict_lo)
  );


  bsg_cache_sbuf_00000080_00000021_00000008
  sbuf
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .sbuf_entry_i({ addr_v_r, sbuf_entry_li_data__127_, sbuf_entry_li_data__126_, sbuf_entry_li_data__125_, sbuf_entry_li_data__124_, sbuf_entry_li_data__123_, sbuf_entry_li_data__122_, sbuf_entry_li_data__121_, sbuf_entry_li_data__120_, sbuf_entry_li_data__119_, sbuf_entry_li_data__118_, sbuf_entry_li_data__117_, sbuf_entry_li_data__116_, sbuf_entry_li_data__115_, sbuf_entry_li_data__114_, sbuf_entry_li_data__113_, sbuf_entry_li_data__112_, sbuf_entry_li_data__111_, sbuf_entry_li_data__110_, sbuf_entry_li_data__109_, sbuf_entry_li_data__108_, sbuf_entry_li_data__107_, sbuf_entry_li_data__106_, sbuf_entry_li_data__105_, sbuf_entry_li_data__104_, sbuf_entry_li_data__103_, sbuf_entry_li_data__102_, sbuf_entry_li_data__101_, sbuf_entry_li_data__100_, sbuf_entry_li_data__99_, sbuf_entry_li_data__98_, sbuf_entry_li_data__97_, sbuf_entry_li_data__96_, sbuf_entry_li_data__95_, sbuf_entry_li_data__94_, sbuf_entry_li_data__93_, sbuf_entry_li_data__92_, sbuf_entry_li_data__91_, sbuf_entry_li_data__90_, sbuf_entry_li_data__89_, sbuf_entry_li_data__88_, sbuf_entry_li_data__87_, sbuf_entry_li_data__86_, sbuf_entry_li_data__85_, sbuf_entry_li_data__84_, sbuf_entry_li_data__83_, sbuf_entry_li_data__82_, sbuf_entry_li_data__81_, sbuf_entry_li_data__80_, sbuf_entry_li_data__79_, sbuf_entry_li_data__78_, sbuf_entry_li_data__77_, sbuf_entry_li_data__76_, sbuf_entry_li_data__75_, sbuf_entry_li_data__74_, sbuf_entry_li_data__73_, sbuf_entry_li_data__72_, sbuf_entry_li_data__71_, sbuf_entry_li_data__70_, sbuf_entry_li_data__69_, sbuf_entry_li_data__68_, sbuf_entry_li_data__67_, sbuf_entry_li_data__66_, sbuf_entry_li_data__65_, sbuf_entry_li_data__64_, sbuf_entry_li_data__63_, sbuf_entry_li_data__62_, sbuf_entry_li_data__61_, sbuf_entry_li_data__60_, sbuf_entry_li_data__59_, sbuf_entry_li_data__58_, sbuf_entry_li_data__57_, sbuf_entry_li_data__56_, sbuf_entry_li_data__55_, sbuf_entry_li_data__54_, sbuf_entry_li_data__53_, sbuf_entry_li_data__52_, sbuf_entry_li_data__51_, sbuf_entry_li_data__50_, sbuf_entry_li_data__49_, sbuf_entry_li_data__48_, sbuf_entry_li_data__47_, sbuf_entry_li_data__46_, sbuf_entry_li_data__45_, sbuf_entry_li_data__44_, sbuf_entry_li_data__43_, sbuf_entry_li_data__42_, sbuf_entry_li_data__41_, sbuf_entry_li_data__40_, sbuf_entry_li_data__39_, sbuf_entry_li_data__38_, sbuf_entry_li_data__37_, sbuf_entry_li_data__36_, sbuf_entry_li_data__35_, sbuf_entry_li_data__34_, sbuf_entry_li_data__33_, sbuf_entry_li_data__32_, sbuf_entry_li_data__31_, sbuf_entry_li_data__30_, sbuf_entry_li_data__29_, sbuf_entry_li_data__28_, sbuf_entry_li_data__27_, sbuf_entry_li_data__26_, sbuf_entry_li_data__25_, sbuf_entry_li_data__24_, sbuf_entry_li_data__23_, sbuf_entry_li_data__22_, sbuf_entry_li_data__21_, sbuf_entry_li_data__20_, sbuf_entry_li_data__19_, sbuf_entry_li_data__18_, sbuf_entry_li_data__17_, sbuf_entry_li_data__16_, sbuf_entry_li_data__15_, sbuf_entry_li_data__14_, sbuf_entry_li_data__13_, sbuf_entry_li_data__12_, sbuf_entry_li_data__11_, sbuf_entry_li_data__10_, sbuf_entry_li_data__9_, sbuf_entry_li_data__8_, sbuf_entry_li_data__7_, sbuf_entry_li_data__6_, sbuf_entry_li_data__5_, sbuf_entry_li_data__4_, sbuf_entry_li_data__3_, sbuf_entry_li_data__2_, sbuf_entry_li_data__1_, sbuf_entry_li_data__0_, sbuf_entry_li_mask__15_, sbuf_entry_li_mask__14_, sbuf_entry_li_mask__13_, sbuf_entry_li_mask__12_, sbuf_entry_li_mask__11_, sbuf_entry_li_mask__10_, sbuf_entry_li_mask__9_, sbuf_entry_li_mask__8_, sbuf_entry_li_mask__7_, sbuf_entry_li_mask__6_, sbuf_entry_li_mask__5_, sbuf_entry_li_mask__4_, sbuf_entry_li_mask__3_, sbuf_entry_li_mask__2_, sbuf_entry_li_mask__1_, sbuf_entry_li_mask__0_, sbuf_entry_li_way_id__2_, sbuf_entry_li_way_id__1_, sbuf_entry_li_way_id__0_ }),
    .v_i(sbuf_v_li),
    .sbuf_entry_o(sbuf_entry_lo),
    .v_o(sbuf_v_lo),
    .yumi_i(sbuf_yumi_li),
    .empty_o(sbuf_empty_lo),
    .full_o(sbuf_full_lo),
    .bypass_addr_i(addr_tl_r),
    .bypass_v_i(sbuf_bypass_v_li),
    .bypass_data_o(bypass_data_lo),
    .bypass_mask_o(bypass_mask_lo)
  );


  bsg_decode_00000008
  sbuf_way_demux
  (
    .i(sbuf_entry_lo[2:0]),
    .o(sbuf_way_decode)
  );


  bsg_decode_00000001
  sbuf_bo_demux
  (
    .i(sbuf_entry_lo[151]),
    .o(sbuf_burst_offset_decode[0])
  );


  bsg_expand_bitmask_00000001_00000010
  expand0
  (
    .i(sbuf_burst_offset_decode[0]),
    .o(sbuf_expand_mask)
  );


  bsg_mux_00000080_00000004
  sbuf_data_in_mux
  (
    .data_i({ \sbuf_in_sel_3_.slice_data , \sbuf_in_sel_3_.slice_data , \sbuf_in_sel_2_.slice_data , \sbuf_in_sel_2_.slice_data , \sbuf_in_sel_2_.slice_data , \sbuf_in_sel_2_.slice_data , data_v_r[15:0], data_v_r[15:0], data_v_r[15:0], data_v_r[15:0], data_v_r[15:0], data_v_r[15:0], data_v_r[15:0], data_v_r[15:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0] }),
    .sel_i(decode_v_r[20:19]),
    .data_o(sbuf_data_in)
  );


  bsg_mux_00000010_00000004
  sbuf_mask_in_mux
  (
    .data_i(sbuf_mask_in_mux_li),
    .sel_i(decode_v_r[20:19]),
    .data_o(sbuf_mask_in)
  );

  assign N358 = N357 | decode_v_r[3];
  assign N359 = decode_v_r[2] | decode_v_r[1];
  assign N360 = N358 | N359;
  assign N361 = N360 | decode_v_r[0];
  assign N365 = N357 | decode_v_r[3];
  assign N366 = decode_v_r[2] | N363;
  assign N367 = N365 | N366;
  assign N368 = N367 | N364;
  assign N371 = N357 | decode_v_r[3];
  assign N372 = N370 | decode_v_r[1];
  assign N373 = N371 | N372;
  assign N374 = N373 | decode_v_r[0];
  assign N377 = N357 | decode_v_r[3];
  assign N378 = decode_v_r[2] | N376;
  assign N379 = N377 | N378;
  assign N380 = N379 | decode_v_r[0];
  assign N383 = N357 | decode_v_r[3];
  assign N384 = decode_v_r[2] | decode_v_r[1];
  assign N385 = N383 | N384;
  assign N386 = N385 | N382;
  assign N390 = N357 | decode_v_r[3];
  assign N391 = N388 | decode_v_r[1];
  assign N392 = N390 | N391;
  assign N393 = N392 | N389;
  assign N397 = N357 | decode_v_r[3];
  assign N398 = N395 | N396;
  assign N399 = N397 | N398;
  assign N400 = N399 | decode_v_r[0];
  assign N405 = N357 | decode_v_r[3];
  assign N406 = N402 | N403;
  assign N407 = N405 | N406;
  assign N408 = N407 | N404;
  assign N411 = N357 | N410;
  assign N412 = decode_v_r[2] | decode_v_r[1];
  assign N413 = N411 | N412;
  assign N414 = N413 | decode_v_r[0];
  assign N416 = N356 & decode_v_r[3];
  assign N417 = N416 & decode_v_r[0];
  assign N418 = N356 & decode_v_r[3];
  assign N419 = N418 & decode_v_r[1];
  assign N420 = N356 & decode_v_r[3];
  assign N421 = N420 & decode_v_r[2];
  assign N679 = $signed(atomic_reg_data) < $signed(atomic_mem_data);
  assign N745 = $signed(atomic_reg_data) > $signed(atomic_mem_data);
  assign N811 = atomic_reg_data < atomic_mem_data;
  assign N877 = atomic_reg_data > atomic_mem_data;

  bsg_decode_00000010
  \sbuf_in_sel_0_.dec 
  (
    .i(addr_v_r[3:0]),
    .o(\sbuf_in_sel_0_.decode_lo )
  );


  bsg_expand_bitmask_00000010_1
  \sbuf_in_sel_0_.exp 
  (
    .i(\sbuf_in_sel_0_.decode_lo ),
    .o(sbuf_mask_in_mux_li[15:0])
  );


  bsg_decode_00000008
  \sbuf_in_sel_1_.dec 
  (
    .i(addr_v_r[3:1]),
    .o(\sbuf_in_sel_1_.decode_lo )
  );


  bsg_expand_bitmask_00000008_2
  \sbuf_in_sel_1_.exp 
  (
    .i(\sbuf_in_sel_1_.decode_lo ),
    .o(sbuf_mask_in_mux_li[31:16])
  );


  bsg_decode_00000004
  \sbuf_in_sel_2_.dec 
  (
    .i(addr_v_r[3:2]),
    .o(\sbuf_in_sel_2_.decode_lo )
  );


  bsg_expand_bitmask_00000004_4
  \sbuf_in_sel_2_.exp 
  (
    .i(\sbuf_in_sel_2_.decode_lo ),
    .o(sbuf_mask_in_mux_li[47:32])
  );


  bsg_decode_00000002
  \sbuf_in_sel_3_.dec 
  (
    .i(addr_v_r[3]),
    .o(\sbuf_in_sel_3_.decode_lo )
  );


  bsg_expand_bitmask_00000002_8
  \sbuf_in_sel_3_.exp 
  (
    .i(\sbuf_in_sel_3_.decode_lo ),
    .o(sbuf_mask_in_mux_li[63:48])
  );


  bsg_cache_tbuf_00000080_00000021_00000008
  \tbuf_gen.tbuf 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .addr_i(addr_v_r),
    .way_i(tbuf_way_li),
    .v_i(tbuf_v_li),
    .addr_o(tbuf_addr_lo),
    .way_o(tbuf_way_lo),
    .v_o(tbuf_v_lo),
    .yumi_i(tbuf_yumi_li),
    .empty_o(tbuf_empty_lo),
    .full_o(tbuf_full_lo),
    .bypass_addr_i(addr_tl_r),
    .bypass_v_i(tbuf_bypass_v_li),
    .bypass_track_o(bypass_track_lo)
  );


  bsg_decode_00000008
  tbuf_way_demux
  (
    .i(tbuf_way_lo),
    .o(tbuf_way_decode)
  );


  bsg_decode_00000004
  tbuf_wo_demux
  (
    .i(tbuf_addr_lo[5:4]),
    .o(tbuf_word_offset_decode)
  );


  bsg_mux_00000080_00000008
  ld_data_mux
  (
    .data_i(ld_data_v_r),
    .sel_i(tag_hit_way_id),
    .data_o(ld_data_way_picked)
  );


  bsg_mux_00000080_00000001
  mux00
  (
    .data_i(ld_data_way_picked),
    .sel_i(addr_v_r[4]),
    .data_o(ld_data_offset_picked)
  );


  bsg_mux_segmented_00000010_8
  bypass_mux_segmented
  (
    .data0_i(ld_data_offset_picked),
    .data1_i(bypass_data_lo),
    .sel_i(bypass_mask_lo),
    .data_o(bypass_data_masked)
  );


  bsg_expand_bitmask_00000010_8
  mask_v_expand
  (
    .i(mask_v_r),
    .o(expanded_mask_v)
  );


  bsg_mux_8_00000010
  \ld_data_sel_0_.byte_mux 
  (
    .data_i(snoop_or_ld_data),
    .sel_i(addr_v_r[3:0]),
    .data_o(\ld_data_sel_0_.byte_sel )
  );


  bsg_mux_16_00000008
  \ld_data_sel_1_.byte_mux 
  (
    .data_i(snoop_or_ld_data),
    .sel_i(addr_v_r[3:1]),
    .data_o(\ld_data_sel_1_.byte_sel )
  );


  bsg_mux_32_00000004
  \ld_data_sel_2_.byte_mux 
  (
    .data_i(snoop_or_ld_data),
    .sel_i(addr_v_r[3:2]),
    .data_o(\atomic_64.amo32_mem_in )
  );


  bsg_mux_64_00000002
  \ld_data_sel_3_.byte_mux 
  (
    .data_i(snoop_or_ld_data),
    .sel_i(addr_v_r[3]),
    .data_o(\atomic_64.amo64_mem_in )
  );


  bsg_mux_00000080_00000004
  ld_data_size_mux
  (
    .data_i({ ld_data_final_li_3__127_, ld_data_final_li_3__126_, ld_data_final_li_3__125_, ld_data_final_li_3__124_, ld_data_final_li_3__123_, ld_data_final_li_3__122_, ld_data_final_li_3__121_, ld_data_final_li_3__120_, ld_data_final_li_3__119_, ld_data_final_li_3__118_, ld_data_final_li_3__117_, ld_data_final_li_3__116_, ld_data_final_li_3__115_, ld_data_final_li_3__114_, ld_data_final_li_3__113_, ld_data_final_li_3__112_, ld_data_final_li_3__111_, ld_data_final_li_3__110_, ld_data_final_li_3__109_, ld_data_final_li_3__108_, ld_data_final_li_3__107_, ld_data_final_li_3__106_, ld_data_final_li_3__105_, ld_data_final_li_3__104_, ld_data_final_li_3__103_, ld_data_final_li_3__102_, ld_data_final_li_3__101_, ld_data_final_li_3__100_, ld_data_final_li_3__99_, ld_data_final_li_3__98_, ld_data_final_li_3__97_, ld_data_final_li_3__96_, ld_data_final_li_3__95_, ld_data_final_li_3__94_, ld_data_final_li_3__93_, ld_data_final_li_3__92_, ld_data_final_li_3__91_, ld_data_final_li_3__90_, ld_data_final_li_3__89_, ld_data_final_li_3__88_, ld_data_final_li_3__87_, ld_data_final_li_3__86_, ld_data_final_li_3__85_, ld_data_final_li_3__84_, ld_data_final_li_3__83_, ld_data_final_li_3__82_, ld_data_final_li_3__81_, ld_data_final_li_3__80_, ld_data_final_li_3__79_, ld_data_final_li_3__78_, ld_data_final_li_3__77_, ld_data_final_li_3__76_, ld_data_final_li_3__75_, ld_data_final_li_3__74_, ld_data_final_li_3__73_, ld_data_final_li_3__72_, ld_data_final_li_3__71_, ld_data_final_li_3__70_, ld_data_final_li_3__69_, ld_data_final_li_3__68_, ld_data_final_li_3__67_, ld_data_final_li_3__66_, ld_data_final_li_3__65_, ld_data_final_li_3__64_, \atomic_64.amo64_mem_in , ld_data_final_li_2__127_, ld_data_final_li_2__126_, ld_data_final_li_2__125_, ld_data_final_li_2__124_, ld_data_final_li_2__123_, ld_data_final_li_2__122_, ld_data_final_li_2__121_, ld_data_final_li_2__120_, ld_data_final_li_2__119_, ld_data_final_li_2__118_, ld_data_final_li_2__117_, ld_data_final_li_2__116_, ld_data_final_li_2__115_, ld_data_final_li_2__114_, ld_data_final_li_2__113_, ld_data_final_li_2__112_, ld_data_final_li_2__111_, ld_data_final_li_2__110_, ld_data_final_li_2__109_, ld_data_final_li_2__108_, ld_data_final_li_2__107_, ld_data_final_li_2__106_, ld_data_final_li_2__105_, ld_data_final_li_2__104_, ld_data_final_li_2__103_, ld_data_final_li_2__102_, ld_data_final_li_2__101_, ld_data_final_li_2__100_, ld_data_final_li_2__99_, ld_data_final_li_2__98_, ld_data_final_li_2__97_, ld_data_final_li_2__96_, ld_data_final_li_2__95_, ld_data_final_li_2__94_, ld_data_final_li_2__93_, ld_data_final_li_2__92_, ld_data_final_li_2__91_, ld_data_final_li_2__90_, ld_data_final_li_2__89_, ld_data_final_li_2__88_, ld_data_final_li_2__87_, ld_data_final_li_2__86_, ld_data_final_li_2__85_, ld_data_final_li_2__84_, ld_data_final_li_2__83_, ld_data_final_li_2__82_, ld_data_final_li_2__81_, ld_data_final_li_2__80_, ld_data_final_li_2__79_, ld_data_final_li_2__78_, ld_data_final_li_2__77_, ld_data_final_li_2__76_, ld_data_final_li_2__75_, ld_data_final_li_2__74_, ld_data_final_li_2__73_, ld_data_final_li_2__72_, ld_data_final_li_2__71_, ld_data_final_li_2__70_, ld_data_final_li_2__69_, ld_data_final_li_2__68_, ld_data_final_li_2__67_, ld_data_final_li_2__66_, ld_data_final_li_2__65_, ld_data_final_li_2__64_, ld_data_final_li_2__63_, ld_data_final_li_2__62_, ld_data_final_li_2__61_, ld_data_final_li_2__60_, ld_data_final_li_2__59_, ld_data_final_li_2__58_, ld_data_final_li_2__57_, ld_data_final_li_2__56_, ld_data_final_li_2__55_, ld_data_final_li_2__54_, ld_data_final_li_2__53_, ld_data_final_li_2__52_, ld_data_final_li_2__51_, ld_data_final_li_2__50_, ld_data_final_li_2__49_, ld_data_final_li_2__48_, ld_data_final_li_2__47_, ld_data_final_li_2__46_, ld_data_final_li_2__45_, ld_data_final_li_2__44_, ld_data_final_li_2__43_, ld_data_final_li_2__42_, ld_data_final_li_2__41_, ld_data_final_li_2__40_, ld_data_final_li_2__39_, ld_data_final_li_2__38_, ld_data_final_li_2__37_, ld_data_final_li_2__36_, ld_data_final_li_2__35_, ld_data_final_li_2__34_, ld_data_final_li_2__33_, ld_data_final_li_2__32_, \atomic_64.amo32_mem_in , ld_data_final_li_1__127_, ld_data_final_li_1__126_, ld_data_final_li_1__125_, ld_data_final_li_1__124_, ld_data_final_li_1__123_, ld_data_final_li_1__122_, ld_data_final_li_1__121_, ld_data_final_li_1__120_, ld_data_final_li_1__119_, ld_data_final_li_1__118_, ld_data_final_li_1__117_, ld_data_final_li_1__116_, ld_data_final_li_1__115_, ld_data_final_li_1__114_, ld_data_final_li_1__113_, ld_data_final_li_1__112_, ld_data_final_li_1__111_, ld_data_final_li_1__110_, ld_data_final_li_1__109_, ld_data_final_li_1__108_, ld_data_final_li_1__107_, ld_data_final_li_1__106_, ld_data_final_li_1__105_, ld_data_final_li_1__104_, ld_data_final_li_1__103_, ld_data_final_li_1__102_, ld_data_final_li_1__101_, ld_data_final_li_1__100_, ld_data_final_li_1__99_, ld_data_final_li_1__98_, ld_data_final_li_1__97_, ld_data_final_li_1__96_, ld_data_final_li_1__95_, ld_data_final_li_1__94_, ld_data_final_li_1__93_, ld_data_final_li_1__92_, ld_data_final_li_1__91_, ld_data_final_li_1__90_, ld_data_final_li_1__89_, ld_data_final_li_1__88_, ld_data_final_li_1__87_, ld_data_final_li_1__86_, ld_data_final_li_1__85_, ld_data_final_li_1__84_, ld_data_final_li_1__83_, ld_data_final_li_1__82_, ld_data_final_li_1__81_, ld_data_final_li_1__80_, ld_data_final_li_1__79_, ld_data_final_li_1__78_, ld_data_final_li_1__77_, ld_data_final_li_1__76_, ld_data_final_li_1__75_, ld_data_final_li_1__74_, ld_data_final_li_1__73_, ld_data_final_li_1__72_, ld_data_final_li_1__71_, ld_data_final_li_1__70_, ld_data_final_li_1__69_, ld_data_final_li_1__68_, ld_data_final_li_1__67_, ld_data_final_li_1__66_, ld_data_final_li_1__65_, ld_data_final_li_1__64_, ld_data_final_li_1__63_, ld_data_final_li_1__62_, ld_data_final_li_1__61_, ld_data_final_li_1__60_, ld_data_final_li_1__59_, ld_data_final_li_1__58_, ld_data_final_li_1__57_, ld_data_final_li_1__56_, ld_data_final_li_1__55_, ld_data_final_li_1__54_, ld_data_final_li_1__53_, ld_data_final_li_1__52_, ld_data_final_li_1__51_, ld_data_final_li_1__50_, ld_data_final_li_1__49_, ld_data_final_li_1__48_, ld_data_final_li_1__47_, ld_data_final_li_1__46_, ld_data_final_li_1__45_, ld_data_final_li_1__44_, ld_data_final_li_1__43_, ld_data_final_li_1__42_, ld_data_final_li_1__41_, ld_data_final_li_1__40_, ld_data_final_li_1__39_, ld_data_final_li_1__38_, ld_data_final_li_1__37_, ld_data_final_li_1__36_, ld_data_final_li_1__35_, ld_data_final_li_1__34_, ld_data_final_li_1__33_, ld_data_final_li_1__32_, ld_data_final_li_1__31_, ld_data_final_li_1__30_, ld_data_final_li_1__29_, ld_data_final_li_1__28_, ld_data_final_li_1__27_, ld_data_final_li_1__26_, ld_data_final_li_1__25_, ld_data_final_li_1__24_, ld_data_final_li_1__23_, ld_data_final_li_1__22_, ld_data_final_li_1__21_, ld_data_final_li_1__20_, ld_data_final_li_1__19_, ld_data_final_li_1__18_, ld_data_final_li_1__17_, ld_data_final_li_1__16_, \ld_data_sel_1_.byte_sel , ld_data_final_li_0__127_, ld_data_final_li_0__126_, ld_data_final_li_0__125_, ld_data_final_li_0__124_, ld_data_final_li_0__123_, ld_data_final_li_0__122_, ld_data_final_li_0__121_, ld_data_final_li_0__120_, ld_data_final_li_0__119_, ld_data_final_li_0__118_, ld_data_final_li_0__117_, ld_data_final_li_0__116_, ld_data_final_li_0__115_, ld_data_final_li_0__114_, ld_data_final_li_0__113_, ld_data_final_li_0__112_, ld_data_final_li_0__111_, ld_data_final_li_0__110_, ld_data_final_li_0__109_, ld_data_final_li_0__108_, ld_data_final_li_0__107_, ld_data_final_li_0__106_, ld_data_final_li_0__105_, ld_data_final_li_0__104_, ld_data_final_li_0__103_, ld_data_final_li_0__102_, ld_data_final_li_0__101_, ld_data_final_li_0__100_, ld_data_final_li_0__99_, ld_data_final_li_0__98_, ld_data_final_li_0__97_, ld_data_final_li_0__96_, ld_data_final_li_0__95_, ld_data_final_li_0__94_, ld_data_final_li_0__93_, ld_data_final_li_0__92_, ld_data_final_li_0__91_, ld_data_final_li_0__90_, ld_data_final_li_0__89_, ld_data_final_li_0__88_, ld_data_final_li_0__87_, ld_data_final_li_0__86_, ld_data_final_li_0__85_, ld_data_final_li_0__84_, ld_data_final_li_0__83_, ld_data_final_li_0__82_, ld_data_final_li_0__81_, ld_data_final_li_0__80_, ld_data_final_li_0__79_, ld_data_final_li_0__78_, ld_data_final_li_0__77_, ld_data_final_li_0__76_, ld_data_final_li_0__75_, ld_data_final_li_0__74_, ld_data_final_li_0__73_, ld_data_final_li_0__72_, ld_data_final_li_0__71_, ld_data_final_li_0__70_, ld_data_final_li_0__69_, ld_data_final_li_0__68_, ld_data_final_li_0__67_, ld_data_final_li_0__66_, ld_data_final_li_0__65_, ld_data_final_li_0__64_, ld_data_final_li_0__63_, ld_data_final_li_0__62_, ld_data_final_li_0__61_, ld_data_final_li_0__60_, ld_data_final_li_0__59_, ld_data_final_li_0__58_, ld_data_final_li_0__57_, ld_data_final_li_0__56_, ld_data_final_li_0__55_, ld_data_final_li_0__54_, ld_data_final_li_0__53_, ld_data_final_li_0__52_, ld_data_final_li_0__51_, ld_data_final_li_0__50_, ld_data_final_li_0__49_, ld_data_final_li_0__48_, ld_data_final_li_0__47_, ld_data_final_li_0__46_, ld_data_final_li_0__45_, ld_data_final_li_0__44_, ld_data_final_li_0__43_, ld_data_final_li_0__42_, ld_data_final_li_0__41_, ld_data_final_li_0__40_, ld_data_final_li_0__39_, ld_data_final_li_0__38_, ld_data_final_li_0__37_, ld_data_final_li_0__36_, ld_data_final_li_0__35_, ld_data_final_li_0__34_, ld_data_final_li_0__33_, ld_data_final_li_0__32_, ld_data_final_li_0__31_, ld_data_final_li_0__30_, ld_data_final_li_0__29_, ld_data_final_li_0__28_, ld_data_final_li_0__27_, ld_data_final_li_0__26_, ld_data_final_li_0__25_, ld_data_final_li_0__24_, ld_data_final_li_0__23_, ld_data_final_li_0__22_, ld_data_final_li_0__21_, ld_data_final_li_0__20_, ld_data_final_li_0__19_, ld_data_final_li_0__18_, ld_data_final_li_0__17_, ld_data_final_li_0__16_, ld_data_final_li_0__15_, ld_data_final_li_0__14_, ld_data_final_li_0__13_, ld_data_final_li_0__12_, ld_data_final_li_0__11_, ld_data_final_li_0__10_, ld_data_final_li_0__9_, ld_data_final_li_0__8_, \ld_data_sel_0_.byte_sel  }),
    .sel_i(decode_v_r[20:19]),
    .data_o(ld_data_final_lo)
  );

  assign N982 = (N974)? lock_v_r[0] : 
                (N976)? lock_v_r[1] : 
                (N978)? lock_v_r[2] : 
                (N980)? lock_v_r[3] : 
                (N975)? lock_v_r[4] : 
                (N977)? lock_v_r[5] : 
                (N979)? lock_v_r[6] : 
                (N981)? lock_v_r[7] : 1'b0;
  assign N998 = (N990)? valid_v_r[0] : 
                (N992)? valid_v_r[1] : 
                (N994)? valid_v_r[2] : 
                (N996)? valid_v_r[3] : 
                (N991)? valid_v_r[4] : 
                (N993)? valid_v_r[5] : 
                (N995)? valid_v_r[6] : 
                (N997)? valid_v_r[7] : 1'b0;
  assign N1014 = (N1006)? tag_v_r[19] : 
                 (N1008)? tag_v_r[39] : 
                 (N1010)? tag_v_r[59] : 
                 (N1012)? tag_v_r[79] : 
                 (N1007)? tag_v_r[99] : 
                 (N1009)? tag_v_r[119] : 
                 (N1011)? tag_v_r[139] : 
                 (N1013)? tag_v_r[159] : 1'b0;
  assign N1015 = (N1006)? tag_v_r[18] : 
                 (N1008)? tag_v_r[38] : 
                 (N1010)? tag_v_r[58] : 
                 (N1012)? tag_v_r[78] : 
                 (N1007)? tag_v_r[98] : 
                 (N1009)? tag_v_r[118] : 
                 (N1011)? tag_v_r[138] : 
                 (N1013)? tag_v_r[158] : 1'b0;
  assign N1016 = (N1006)? tag_v_r[17] : 
                 (N1008)? tag_v_r[37] : 
                 (N1010)? tag_v_r[57] : 
                 (N1012)? tag_v_r[77] : 
                 (N1007)? tag_v_r[97] : 
                 (N1009)? tag_v_r[117] : 
                 (N1011)? tag_v_r[137] : 
                 (N1013)? tag_v_r[157] : 1'b0;
  assign N1017 = (N1006)? tag_v_r[16] : 
                 (N1008)? tag_v_r[36] : 
                 (N1010)? tag_v_r[56] : 
                 (N1012)? tag_v_r[76] : 
                 (N1007)? tag_v_r[96] : 
                 (N1009)? tag_v_r[116] : 
                 (N1011)? tag_v_r[136] : 
                 (N1013)? tag_v_r[156] : 1'b0;
  assign N1018 = (N1006)? tag_v_r[15] : 
                 (N1008)? tag_v_r[35] : 
                 (N1010)? tag_v_r[55] : 
                 (N1012)? tag_v_r[75] : 
                 (N1007)? tag_v_r[95] : 
                 (N1009)? tag_v_r[115] : 
                 (N1011)? tag_v_r[135] : 
                 (N1013)? tag_v_r[155] : 1'b0;
  assign N1019 = (N1006)? tag_v_r[14] : 
                 (N1008)? tag_v_r[34] : 
                 (N1010)? tag_v_r[54] : 
                 (N1012)? tag_v_r[74] : 
                 (N1007)? tag_v_r[94] : 
                 (N1009)? tag_v_r[114] : 
                 (N1011)? tag_v_r[134] : 
                 (N1013)? tag_v_r[154] : 1'b0;
  assign N1020 = (N1006)? tag_v_r[13] : 
                 (N1008)? tag_v_r[33] : 
                 (N1010)? tag_v_r[53] : 
                 (N1012)? tag_v_r[73] : 
                 (N1007)? tag_v_r[93] : 
                 (N1009)? tag_v_r[113] : 
                 (N1011)? tag_v_r[133] : 
                 (N1013)? tag_v_r[153] : 1'b0;
  assign N1021 = (N1006)? tag_v_r[12] : 
                 (N1008)? tag_v_r[32] : 
                 (N1010)? tag_v_r[52] : 
                 (N1012)? tag_v_r[72] : 
                 (N1007)? tag_v_r[92] : 
                 (N1009)? tag_v_r[112] : 
                 (N1011)? tag_v_r[132] : 
                 (N1013)? tag_v_r[152] : 1'b0;
  assign N1022 = (N1006)? tag_v_r[11] : 
                 (N1008)? tag_v_r[31] : 
                 (N1010)? tag_v_r[51] : 
                 (N1012)? tag_v_r[71] : 
                 (N1007)? tag_v_r[91] : 
                 (N1009)? tag_v_r[111] : 
                 (N1011)? tag_v_r[131] : 
                 (N1013)? tag_v_r[151] : 1'b0;
  assign N1023 = (N1006)? tag_v_r[10] : 
                 (N1008)? tag_v_r[30] : 
                 (N1010)? tag_v_r[50] : 
                 (N1012)? tag_v_r[70] : 
                 (N1007)? tag_v_r[90] : 
                 (N1009)? tag_v_r[110] : 
                 (N1011)? tag_v_r[130] : 
                 (N1013)? tag_v_r[150] : 1'b0;
  assign N1024 = (N1006)? tag_v_r[9] : 
                 (N1008)? tag_v_r[29] : 
                 (N1010)? tag_v_r[49] : 
                 (N1012)? tag_v_r[69] : 
                 (N1007)? tag_v_r[89] : 
                 (N1009)? tag_v_r[109] : 
                 (N1011)? tag_v_r[129] : 
                 (N1013)? tag_v_r[149] : 1'b0;
  assign N1025 = (N1006)? tag_v_r[8] : 
                 (N1008)? tag_v_r[28] : 
                 (N1010)? tag_v_r[48] : 
                 (N1012)? tag_v_r[68] : 
                 (N1007)? tag_v_r[88] : 
                 (N1009)? tag_v_r[108] : 
                 (N1011)? tag_v_r[128] : 
                 (N1013)? tag_v_r[148] : 1'b0;
  assign N1026 = (N1006)? tag_v_r[7] : 
                 (N1008)? tag_v_r[27] : 
                 (N1010)? tag_v_r[47] : 
                 (N1012)? tag_v_r[67] : 
                 (N1007)? tag_v_r[87] : 
                 (N1009)? tag_v_r[107] : 
                 (N1011)? tag_v_r[127] : 
                 (N1013)? tag_v_r[147] : 1'b0;
  assign N1027 = (N1006)? tag_v_r[6] : 
                 (N1008)? tag_v_r[26] : 
                 (N1010)? tag_v_r[46] : 
                 (N1012)? tag_v_r[66] : 
                 (N1007)? tag_v_r[86] : 
                 (N1009)? tag_v_r[106] : 
                 (N1011)? tag_v_r[126] : 
                 (N1013)? tag_v_r[146] : 1'b0;
  assign N1028 = (N1006)? tag_v_r[5] : 
                 (N1008)? tag_v_r[25] : 
                 (N1010)? tag_v_r[45] : 
                 (N1012)? tag_v_r[65] : 
                 (N1007)? tag_v_r[85] : 
                 (N1009)? tag_v_r[105] : 
                 (N1011)? tag_v_r[125] : 
                 (N1013)? tag_v_r[145] : 1'b0;
  assign N1029 = (N1006)? tag_v_r[4] : 
                 (N1008)? tag_v_r[24] : 
                 (N1010)? tag_v_r[44] : 
                 (N1012)? tag_v_r[64] : 
                 (N1007)? tag_v_r[84] : 
                 (N1009)? tag_v_r[104] : 
                 (N1011)? tag_v_r[124] : 
                 (N1013)? tag_v_r[144] : 1'b0;
  assign N1030 = (N1006)? tag_v_r[3] : 
                 (N1008)? tag_v_r[23] : 
                 (N1010)? tag_v_r[43] : 
                 (N1012)? tag_v_r[63] : 
                 (N1007)? tag_v_r[83] : 
                 (N1009)? tag_v_r[103] : 
                 (N1011)? tag_v_r[123] : 
                 (N1013)? tag_v_r[143] : 1'b0;
  assign N1031 = (N1006)? tag_v_r[2] : 
                 (N1008)? tag_v_r[22] : 
                 (N1010)? tag_v_r[42] : 
                 (N1012)? tag_v_r[62] : 
                 (N1007)? tag_v_r[82] : 
                 (N1009)? tag_v_r[102] : 
                 (N1011)? tag_v_r[122] : 
                 (N1013)? tag_v_r[142] : 1'b0;
  assign N1032 = (N1006)? tag_v_r[1] : 
                 (N1008)? tag_v_r[21] : 
                 (N1010)? tag_v_r[41] : 
                 (N1012)? tag_v_r[61] : 
                 (N1007)? tag_v_r[81] : 
                 (N1009)? tag_v_r[101] : 
                 (N1011)? tag_v_r[121] : 
                 (N1013)? tag_v_r[141] : 1'b0;
  assign N1033 = (N1006)? tag_v_r[0] : 
                 (N1008)? tag_v_r[20] : 
                 (N1010)? tag_v_r[40] : 
                 (N1012)? tag_v_r[60] : 
                 (N1007)? tag_v_r[80] : 
                 (N1009)? tag_v_r[100] : 
                 (N1011)? tag_v_r[120] : 
                 (N1013)? tag_v_r[140] : 1'b0;

  bsg_decode_00000008
  addr_way_demux
  (
    .i(cache_pkt_i[159:157]),
    .o(addr_way_decode)
  );


  bsg_lru_pseudo_tree_decode_00000008
  plru_decode
  (
    .way_id_i(tag_hit_way_id),
    .data_o(plru_decode_data_lo),
    .mask_o(plru_decode_mask_lo)
  );

  assign { N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615 } = atomic_reg_data + atomic_mem_data;
  assign N79 = (N0)? 1'b1 : 
               (N84)? 1'b1 : 
               (N78)? 1'b0 : 1'b0;
  assign N0 = tl_we;
  assign N80 = (N0)? v_i : 
               (N84)? 1'b0 : 1'b0;
  assign N81 = (N0)? v_i : 
               (N84)? 1'b0 : 
               (N78)? 1'b0 : 1'b0;
  assign N82 = (N0)? v_i : 
               (N84)? 1'b0 : 
               (N78)? 1'b0 : 1'b0;
  assign N88 = (N1)? 1'b1 : 
               (N2)? 1'b0 : 1'b0;
  assign N1 = v_we_o;
  assign N89 = (N1)? v_tl_r : 
               (N2)? 1'b0 : 1'b0;
  assign { N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90 } = (N1)? { v_tl_r, v_tl_r, v_tl_r, v_tl_r, v_tl_r, v_tl_r, v_tl_r, v_tl_r, v_tl_r, v_tl_r, v_tl_r, v_tl_r, v_tl_r, v_tl_r } : 
                                                                                        (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104 } = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                (N116)? { v_tl_r, v_tl_r, v_tl_r, v_tl_r, v_tl_r, v_tl_r, v_tl_r, v_tl_r, v_tl_r, v_tl_r, v_tl_r } : 
                                                                                (N87)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N3 = N85;
  assign N127 = (N4)? N126 : 
                (N125)? 1'b1 : 1'b0;
  assign N4 = decode[17];
  assign N130 = (N5)? N129 : 
                (N128)? 1'b1 : 1'b0;
  assign N5 = decode_tl_r[17];
  assign N134 = (N6)? N133 : 
                (N132)? 1'b1 : 1'b0;
  assign N6 = N131;
  assign N196 = (N7)? N195 : 
                (N8)? 1'b1 : 1'b0;
  assign N7 = N178;
  assign N8 = N177;
  assign N215 = (N9)? N214 : 
                (N10)? 1'b0 : 1'b0;
  assign N9 = N198;
  assign N10 = N197;
  assign sbuf_data_mem_w_mask[15:0] = (N11)? { N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232 } : 
                                      (N216)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = sbuf_way_decode[0];
  assign sbuf_data_mem_w_mask[31:16] = (N12)? { N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249 } : 
                                       (N233)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = sbuf_way_decode[1];
  assign sbuf_data_mem_w_mask[47:32] = (N13)? { N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266 } : 
                                       (N250)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = sbuf_way_decode[2];
  assign sbuf_data_mem_w_mask[63:48] = (N14)? { N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283 } : 
                                       (N267)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N14 = sbuf_way_decode[3];
  assign sbuf_data_mem_w_mask[79:64] = (N15)? { N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300 } : 
                                       (N284)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = sbuf_way_decode[4];
  assign sbuf_data_mem_w_mask[95:80] = (N16)? { N302, N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317 } : 
                                       (N301)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = sbuf_way_decode[5];
  assign sbuf_data_mem_w_mask[111:96] = (N17)? { N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334 } : 
                                        (N318)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N17 = sbuf_way_decode[6];
  assign sbuf_data_mem_w_mask[127:112] = (N18)? { N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351 } : 
                                         (N335)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N18 = sbuf_way_decode[7];
  assign atomic_reg_data = (N19)? data_v_r[63:0] : 
                           (N353)? { data_v_r[31:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N19 = N352;
  assign atomic_mem_data = (N20)? \atomic_64.amo64_mem_in  : 
                           (N355)? { \atomic_64.amo32_mem_in , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N20 = N354;
  assign { N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681 } = (N21)? atomic_reg_data : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N680)? atomic_mem_data : 1'b0;
  assign N21 = N679;
  assign { N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747 } = (N22)? atomic_reg_data : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N746)? atomic_mem_data : 1'b0;
  assign N22 = N745;
  assign { N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813 } = (N23)? atomic_reg_data : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N812)? atomic_mem_data : 1'b0;
  assign N23 = N811;
  assign { N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879 } = (N24)? atomic_reg_data : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N878)? atomic_mem_data : 1'b0;
  assign N24 = N877;
  assign atomic_alu_result = (N25)? atomic_reg_data : 
                             (N26)? { N423, N424, N425, N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486 } : 
                             (N27)? { N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546, N547, N548, N549, N550 } : 
                             (N28)? { N551, N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595, N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606, N607, N608, N609, N610, N611, N612, N613, N614 } : 
                             (N29)? { N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615 } : 
                             (N30)? { N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681 } : 
                             (N31)? { N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747 } : 
                             (N32)? { N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813 } : 
                             (N33)? { N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879 } : 
                             (N34)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N25 = N362;
  assign N26 = N369;
  assign N27 = N375;
  assign N28 = N381;
  assign N29 = N387;
  assign N30 = N394;
  assign N31 = N401;
  assign N32 = N409;
  assign N33 = N415;
  assign N34 = N357;
  assign N35 = N422;
  assign atomic_result = (N36)? atomic_alu_result : 
                         (N944)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, atomic_alu_result[63:32] } : 1'b0;
  assign N36 = N943;
  assign \sbuf_in_sel_2_.slice_data  = (N37)? atomic_result[31:0] : 
                                       (N946)? data_v_r[31:0] : 1'b0;
  assign N37 = N945;
  assign \sbuf_in_sel_3_.slice_data  = (N38)? atomic_result : 
                                       (N948)? data_v_r[63:0] : 1'b0;
  assign N38 = N947;
  assign { sbuf_entry_li_data__127_, sbuf_entry_li_data__126_, sbuf_entry_li_data__125_, sbuf_entry_li_data__124_, sbuf_entry_li_data__123_, sbuf_entry_li_data__122_, sbuf_entry_li_data__121_, sbuf_entry_li_data__120_, sbuf_entry_li_data__119_, sbuf_entry_li_data__118_, sbuf_entry_li_data__117_, sbuf_entry_li_data__116_, sbuf_entry_li_data__115_, sbuf_entry_li_data__114_, sbuf_entry_li_data__113_, sbuf_entry_li_data__112_, sbuf_entry_li_data__111_, sbuf_entry_li_data__110_, sbuf_entry_li_data__109_, sbuf_entry_li_data__108_, sbuf_entry_li_data__107_, sbuf_entry_li_data__106_, sbuf_entry_li_data__105_, sbuf_entry_li_data__104_, sbuf_entry_li_data__103_, sbuf_entry_li_data__102_, sbuf_entry_li_data__101_, sbuf_entry_li_data__100_, sbuf_entry_li_data__99_, sbuf_entry_li_data__98_, sbuf_entry_li_data__97_, sbuf_entry_li_data__96_, sbuf_entry_li_data__95_, sbuf_entry_li_data__94_, sbuf_entry_li_data__93_, sbuf_entry_li_data__92_, sbuf_entry_li_data__91_, sbuf_entry_li_data__90_, sbuf_entry_li_data__89_, sbuf_entry_li_data__88_, sbuf_entry_li_data__87_, sbuf_entry_li_data__86_, sbuf_entry_li_data__85_, sbuf_entry_li_data__84_, sbuf_entry_li_data__83_, sbuf_entry_li_data__82_, sbuf_entry_li_data__81_, sbuf_entry_li_data__80_, sbuf_entry_li_data__79_, sbuf_entry_li_data__78_, sbuf_entry_li_data__77_, sbuf_entry_li_data__76_, sbuf_entry_li_data__75_, sbuf_entry_li_data__74_, sbuf_entry_li_data__73_, sbuf_entry_li_data__72_, sbuf_entry_li_data__71_, sbuf_entry_li_data__70_, sbuf_entry_li_data__69_, sbuf_entry_li_data__68_, sbuf_entry_li_data__67_, sbuf_entry_li_data__66_, sbuf_entry_li_data__65_, sbuf_entry_li_data__64_, sbuf_entry_li_data__63_, sbuf_entry_li_data__62_, sbuf_entry_li_data__61_, sbuf_entry_li_data__60_, sbuf_entry_li_data__59_, sbuf_entry_li_data__58_, sbuf_entry_li_data__57_, sbuf_entry_li_data__56_, sbuf_entry_li_data__55_, sbuf_entry_li_data__54_, sbuf_entry_li_data__53_, sbuf_entry_li_data__52_, sbuf_entry_li_data__51_, sbuf_entry_li_data__50_, sbuf_entry_li_data__49_, sbuf_entry_li_data__48_, sbuf_entry_li_data__47_, sbuf_entry_li_data__46_, sbuf_entry_li_data__45_, sbuf_entry_li_data__44_, sbuf_entry_li_data__43_, sbuf_entry_li_data__42_, sbuf_entry_li_data__41_, sbuf_entry_li_data__40_, sbuf_entry_li_data__39_, sbuf_entry_li_data__38_, sbuf_entry_li_data__37_, sbuf_entry_li_data__36_, sbuf_entry_li_data__35_, sbuf_entry_li_data__34_, sbuf_entry_li_data__33_, sbuf_entry_li_data__32_, sbuf_entry_li_data__31_, sbuf_entry_li_data__30_, sbuf_entry_li_data__29_, sbuf_entry_li_data__28_, sbuf_entry_li_data__27_, sbuf_entry_li_data__26_, sbuf_entry_li_data__25_, sbuf_entry_li_data__24_, sbuf_entry_li_data__23_, sbuf_entry_li_data__22_, sbuf_entry_li_data__21_, sbuf_entry_li_data__20_, sbuf_entry_li_data__19_, sbuf_entry_li_data__18_, sbuf_entry_li_data__17_, sbuf_entry_li_data__16_, sbuf_entry_li_data__15_, sbuf_entry_li_data__14_, sbuf_entry_li_data__13_, sbuf_entry_li_data__12_, sbuf_entry_li_data__11_, sbuf_entry_li_data__10_, sbuf_entry_li_data__9_, sbuf_entry_li_data__8_, sbuf_entry_li_data__7_, sbuf_entry_li_data__6_, sbuf_entry_li_data__5_, sbuf_entry_li_data__4_, sbuf_entry_li_data__3_, sbuf_entry_li_data__2_, sbuf_entry_li_data__1_, sbuf_entry_li_data__0_, sbuf_entry_li_mask__15_, sbuf_entry_li_mask__14_, sbuf_entry_li_mask__13_, sbuf_entry_li_mask__12_, sbuf_entry_li_mask__11_, sbuf_entry_li_mask__10_, sbuf_entry_li_mask__9_, sbuf_entry_li_mask__8_, sbuf_entry_li_mask__7_, sbuf_entry_li_mask__6_, sbuf_entry_li_mask__5_, sbuf_entry_li_mask__4_, sbuf_entry_li_mask__3_, sbuf_entry_li_mask__2_, sbuf_entry_li_mask__1_, sbuf_entry_li_mask__0_ } = (N39)? { data_v_r, mask_v_r } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N950)? { sbuf_data_in, sbuf_mask_in } : 1'b0;
  assign N39 = N949;
  assign tbuf_track_mem_w_mask[3:0] = (N40)? tbuf_word_offset_decode : 
                                      (N951)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N40 = tbuf_way_decode[0];
  assign tbuf_track_mem_w_mask[7:4] = (N41)? tbuf_word_offset_decode : 
                                      (N952)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N41 = tbuf_way_decode[1];
  assign tbuf_track_mem_w_mask[11:8] = (N42)? tbuf_word_offset_decode : 
                                       (N953)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N42 = tbuf_way_decode[2];
  assign tbuf_track_mem_w_mask[15:12] = (N43)? tbuf_word_offset_decode : 
                                        (N954)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N43 = tbuf_way_decode[3];
  assign tbuf_track_mem_w_mask[19:16] = (N44)? tbuf_word_offset_decode : 
                                        (N955)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N44 = tbuf_way_decode[4];
  assign tbuf_track_mem_w_mask[23:20] = (N45)? tbuf_word_offset_decode : 
                                        (N956)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N45 = tbuf_way_decode[5];
  assign tbuf_track_mem_w_mask[27:24] = (N46)? tbuf_word_offset_decode : 
                                        (N957)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N46 = tbuf_way_decode[6];
  assign tbuf_track_mem_w_mask[31:28] = (N47)? tbuf_word_offset_decode : 
                                        (N958)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N47 = tbuf_way_decode[7];
  assign snoop_or_ld_data = (N48)? snoop_word_lo : 
                            (N49)? bypass_data_masked : 1'b0;
  assign N48 = select_snoop_data_r_lo;
  assign N49 = N959;
  assign { N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034 } = (N50)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N982, N998 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1163)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033, addr_v_r[12:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1166)? ld_data_masked : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N966)? ld_data_final_lo : 1'b0;
  assign N50 = N961;
  assign data_o = (N51)? { N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034 } : 
                  (N52)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N51 = retval_op_v;
  assign N52 = N960;
  assign N1169 = (N53)? miss_done_lo : 
                 (N54)? 1'b1 : 1'b0;
  assign N53 = N1168;
  assign N54 = N1167;
  assign v_we_o = (N55)? N1171 : 
                  (N56)? 1'b1 : 1'b0;
  assign N55 = v_v_r;
  assign N56 = N1170;
  assign N1175 = (N57)? N1174 : 
                 (N58)? 1'b1 : 1'b0;
  assign N57 = N1173;
  assign N58 = N1172;
  assign N1177 = (N59)? v_we_o : 
                 (N60)? 1'b1 : 1'b0;
  assign N59 = v_tl_r;
  assign N60 = N1176;
  assign tag_mem_w_li = (N61)? N1180 : 
                        (N62)? tagst_write_en : 1'b0;
  assign N61 = N1179;
  assign N62 = N1178;
  assign { N1191, N1190, N1189, N1188, N1187, N1186, N1185 } = (N63)? addr_tl_r[12:6] : 
                                                               (N1193)? miss_tag_mem_addr_lo : 
                                                               (N1184)? cache_pkt_i[156:150] : 1'b0;
  assign N63 = recover_lo;
  assign tag_mem_addr_li = (N64)? { N1191, N1190, N1189, N1188, N1187, N1186, N1185 } : 
                           (N65)? cache_pkt_i[156:150] : 1'b0;
  assign N64 = N1182;
  assign N65 = N1181;
  assign tag_mem_data_li = (N64)? miss_tag_mem_data_lo : 
                           (N65)? { cache_pkt_i[143:142], cache_pkt_i[35:16], cache_pkt_i[143:142], cache_pkt_i[35:16], cache_pkt_i[143:142], cache_pkt_i[35:16], cache_pkt_i[143:142], cache_pkt_i[35:16], cache_pkt_i[143:142], cache_pkt_i[35:16], cache_pkt_i[143:142], cache_pkt_i[35:16], cache_pkt_i[143:142], cache_pkt_i[35:16], cache_pkt_i[143:142], cache_pkt_i[35:16] } : 1'b0;
  assign tag_mem_w_mask_li = (N64)? miss_tag_mem_w_mask_lo : 
                             (N65)? { addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:7], addr_way_decode[7:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:6], addr_way_decode[6:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:5], addr_way_decode[5:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:4], addr_way_decode[4:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0] } : 1'b0;
  assign data_mem_data_li = (N66)? dma_data_mem_data_lo : 
                            (N67)? { sbuf_entry_lo[146:19], sbuf_entry_lo[146:19], sbuf_entry_lo[146:19], sbuf_entry_lo[146:19], sbuf_entry_lo[146:19], sbuf_entry_lo[146:19], sbuf_entry_lo[146:19], sbuf_entry_lo[146:19] } : 1'b0;
  assign N66 = dma_data_mem_w_lo;
  assign N67 = N1194;
  assign data_mem_addr_li = (N63)? addr_tl_r[12:4] : 
                            (N1199)? dma_data_mem_addr_lo : 
                            (N1202)? cache_pkt_i[156:148] : 
                            (N1198)? sbuf_entry_lo[159:151] : 1'b0;
  assign data_mem_w_mask_li = (N66)? dma_data_mem_w_mask_lo : 
                              (N67)? sbuf_data_mem_w_mask : 1'b0;
  assign track_mem_w_li = (N68)? miss_track_mem_w_lo : 
                          (N69)? N1203 : 1'b0;
  assign N68 = miss_track_mem_v_lo;
  assign N69 = N1375;
  assign track_mem_data_li = (N68)? miss_track_mem_data_lo : 
                             (N69)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign track_mem_w_mask_li = (N68)? miss_track_mem_w_mask_lo : 
                               (N69)? tbuf_track_mem_w_mask : 1'b0;
  assign track_mem_addr_li = (N63)? addr_tl_r[12:6] : 
                             (N1208)? miss_track_mem_addr_lo : 
                             (N1211)? cache_pkt_i[156:150] : 
                             (N1207)? tbuf_addr_lo[12:6] : 1'b0;
  assign { N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234 } = (N70)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                       (N1217)? { N1218, N1219, N1220, N1221, N1222, N1223, N1224, N1225, plru_decode_data_lo } : 1'b0;
  assign N70 = N1216;
  assign { N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249 } = (N70)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                       (N1217)? { N1226, N1227, N1228, N1229, N1230, N1231, N1232, N1233, plru_decode_mask_lo } : 1'b0;
  assign stat_mem_v_li = (N71)? miss_stat_mem_v_lo : 
                         (N72)? N1214 : 1'b0;
  assign N71 = N1213;
  assign N72 = N1212;
  assign stat_mem_w_li = (N71)? miss_stat_mem_w_lo : 
                         (N72)? N1215 : 1'b0;
  assign stat_mem_addr_li = (N71)? miss_stat_mem_addr_lo : 
                            (N72)? addr_v_r[12:6] : 1'b0;
  assign stat_mem_data_li = (N71)? miss_stat_mem_data_lo : 
                            (N72)? { N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234 } : 1'b0;
  assign stat_mem_w_mask_li = (N71)? miss_stat_mem_w_mask_lo : 
                              (N72)? { N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249 } : 1'b0;
  assign { sbuf_entry_li_way_id__2_, sbuf_entry_li_way_id__1_, sbuf_entry_li_way_id__0_ } = (N73)? chosen_way_lo : 
                                                                                            (N74)? tag_hit_way_id : 1'b0;
  assign N73 = N1265;
  assign N74 = N1264;
  assign tbuf_way_li = (N75)? chosen_way_lo : 
                       (N76)? tag_hit_way_id : 1'b0;
  assign N75 = N1267;
  assign N76 = N1266;
  assign N356 = (N1284)? 1'b1 : 
                (N1286)? 1'b0 : 
                (N1288)? 1'b0 : 
                (N1290)? 1'b0 : 
                (N1292)? 1'b0 : 
                (N1294)? 1'b0 : 
                (N1296)? 1'b0 : 
                (N1298)? 1'b0 : 
                (N1285)? 1'b0 : 
                (N1287)? 1'b0 : 
                (N1289)? 1'b0 : 
                (N1291)? 1'b0 : 
                (N1293)? 1'b0 : 
                (N1295)? 1'b0 : 
                (N1297)? 1'b0 : 
                (N1299)? 1'b0 : 1'b0;
  assign N77 = sbuf_hazard | tl_we;
  assign N78 = ~N77;
  assign N83 = ~tl_we;
  assign N84 = sbuf_hazard & N83;
  assign N85 = reset_i;
  assign N86 = v_we_o | N85;
  assign N87 = ~N86;
  assign N115 = ~N85;
  assign N116 = v_we_o & N115;
  assign tag_hit_v[0] = N117 & valid_v_r[0];
  assign tag_hit_v[1] = N118 & valid_v_r[1];
  assign tag_hit_v[2] = N119 & valid_v_r[2];
  assign tag_hit_v[3] = N120 & valid_v_r[3];
  assign tag_hit_v[4] = N121 & valid_v_r[4];
  assign tag_hit_v[5] = N122 & valid_v_r[5];
  assign tag_hit_v[6] = N123 & valid_v_r[6];
  assign tag_hit_v[7] = N124 & valid_v_r[7];
  assign N125 = ~decode[17];
  assign N126 = ~N1314;
  assign N1314 = N1313 & cache_pkt_i[0];
  assign N1313 = N1312 & cache_pkt_i[1];
  assign N1312 = N1311 & cache_pkt_i[2];
  assign N1311 = N1310 & cache_pkt_i[3];
  assign N1310 = N1309 & cache_pkt_i[4];
  assign N1309 = N1308 & cache_pkt_i[5];
  assign N1308 = N1307 & cache_pkt_i[6];
  assign N1307 = N1306 & cache_pkt_i[7];
  assign N1306 = N1305 & cache_pkt_i[8];
  assign N1305 = N1304 & cache_pkt_i[9];
  assign N1304 = N1303 & cache_pkt_i[10];
  assign N1303 = N1302 & cache_pkt_i[11];
  assign N1302 = N1301 & cache_pkt_i[12];
  assign N1301 = N1300 & cache_pkt_i[13];
  assign N1300 = cache_pkt_i[15] & cache_pkt_i[14];
  assign partial_st = decode[15] & N127;
  assign N128 = ~decode_tl_r[17];
  assign N129 = ~N1329;
  assign N1329 = N1328 & mask_tl_r[0];
  assign N1328 = N1327 & mask_tl_r[1];
  assign N1327 = N1326 & mask_tl_r[2];
  assign N1326 = N1325 & mask_tl_r[3];
  assign N1325 = N1324 & mask_tl_r[4];
  assign N1324 = N1323 & mask_tl_r[5];
  assign N1323 = N1322 & mask_tl_r[6];
  assign N1322 = N1321 & mask_tl_r[7];
  assign N1321 = N1320 & mask_tl_r[8];
  assign N1320 = N1319 & mask_tl_r[9];
  assign N1319 = N1318 & mask_tl_r[10];
  assign N1318 = N1317 & mask_tl_r[11];
  assign N1317 = N1316 & mask_tl_r[12];
  assign N1316 = N1315 & mask_tl_r[13];
  assign N1315 = mask_tl_r[15] & mask_tl_r[14];
  assign partial_st_tl = decode_tl_r[15] & N130;
  assign N131 = decode_v_r[17];
  assign N132 = ~N131;
  assign N133 = ~N1344;
  assign N1344 = N1343 & mask_v_r[0];
  assign N1343 = N1342 & mask_v_r[1];
  assign N1342 = N1341 & mask_v_r[2];
  assign N1341 = N1340 & mask_v_r[3];
  assign N1340 = N1339 & mask_v_r[4];
  assign N1339 = N1338 & mask_v_r[5];
  assign N1338 = N1337 & mask_v_r[6];
  assign N1337 = N1336 & mask_v_r[7];
  assign N1336 = N1335 & mask_v_r[8];
  assign N1335 = N1334 & mask_v_r[9];
  assign N1334 = N1333 & mask_v_r[10];
  assign N1333 = N1332 & mask_v_r[11];
  assign N1332 = N1331 & mask_v_r[12];
  assign N1331 = N1330 & mask_v_r[13];
  assign N1330 = mask_v_r[15] & mask_v_r[14];
  assign partial_st_v = decode_v_r[15] & N134;
  assign ld_st_amo_tag_miss = N1346 & N1347;
  assign N1346 = N1345 | decode_v_r[4];
  assign N1345 = decode_v_r[16] | decode_v_r[15];
  assign N1347 = ~tag_hit_found;
  assign N135 = ~tag_hit_way_id[0];
  assign N136 = ~tag_hit_way_id[1];
  assign N137 = N135 & N136;
  assign N138 = N135 & tag_hit_way_id[1];
  assign N139 = tag_hit_way_id[0] & N136;
  assign N140 = tag_hit_way_id[0] & tag_hit_way_id[1];
  assign N141 = ~tag_hit_way_id[2];
  assign N142 = N137 & N141;
  assign N143 = N137 & tag_hit_way_id[2];
  assign N144 = N139 & N141;
  assign N145 = N139 & tag_hit_way_id[2];
  assign N146 = N138 & N141;
  assign N147 = N138 & tag_hit_way_id[2];
  assign N148 = N140 & N141;
  assign N149 = N140 & tag_hit_way_id[2];
  assign N154 = ~addr_v_r[4];
  assign N155 = ~addr_v_r[5];
  assign N156 = N154 & N155;
  assign N157 = N154 & addr_v_r[5];
  assign N158 = addr_v_r[4] & N155;
  assign N159 = addr_v_r[4] & addr_v_r[5];
  assign track_miss = N1350 & N1352;
  assign N1350 = N1349 & tag_hit_found;
  assign N1349 = N1348 | partial_st_v;
  assign N1348 = decode_v_r[16] | decode_v_r[4];
  assign N1352 = ~N1351;
  assign N1351 = N160 | bypass_track_lo;
  assign N161 = ~addr_v_r[13];
  assign N162 = ~addr_v_r[14];
  assign N163 = N161 & N162;
  assign N164 = N161 & addr_v_r[14];
  assign N165 = addr_v_r[13] & N162;
  assign N166 = addr_v_r[13] & addr_v_r[14];
  assign N167 = ~addr_v_r[15];
  assign N168 = N163 & N167;
  assign N169 = N163 & addr_v_r[15];
  assign N170 = N165 & N167;
  assign N171 = N165 & addr_v_r[15];
  assign N172 = N164 & N167;
  assign N173 = N164 & addr_v_r[15];
  assign N174 = N166 & N167;
  assign N175 = N166 & addr_v_r[15];
  assign tagfl_hit = decode_v_r[13] & N176;
  assign aflinv_hit = N1354 & tag_hit_found;
  assign N1354 = N1353 | decode_v_r[8];
  assign N1353 = decode_v_r[10] | decode_v_r[9];
  assign N177 = ~tag_hit_found;
  assign N178 = tag_hit_found;
  assign N179 = ~tag_hit_way_id[0];
  assign N180 = ~tag_hit_way_id[1];
  assign N181 = N179 & N180;
  assign N182 = N179 & tag_hit_way_id[1];
  assign N183 = tag_hit_way_id[0] & N180;
  assign N184 = tag_hit_way_id[0] & tag_hit_way_id[1];
  assign N185 = ~tag_hit_way_id[2];
  assign N186 = N181 & N185;
  assign N187 = N181 & tag_hit_way_id[2];
  assign N188 = N183 & N185;
  assign N189 = N183 & tag_hit_way_id[2];
  assign N190 = N182 & N185;
  assign N191 = N182 & tag_hit_way_id[2];
  assign N192 = N184 & N185;
  assign N193 = N184 & tag_hit_way_id[2];
  assign N195 = ~N194;
  assign alock_miss = decode_v_r[7] & N196;
  assign N197 = ~tag_hit_found;
  assign N198 = tag_hit_found;
  assign N199 = ~tag_hit_way_id[0];
  assign N200 = ~tag_hit_way_id[1];
  assign N201 = N199 & N200;
  assign N202 = N199 & tag_hit_way_id[1];
  assign N203 = tag_hit_way_id[0] & N200;
  assign N204 = tag_hit_way_id[0] & tag_hit_way_id[1];
  assign N205 = ~tag_hit_way_id[2];
  assign N206 = N201 & N205;
  assign N207 = N201 & tag_hit_way_id[2];
  assign N208 = N203 & N205;
  assign N209 = N203 & tag_hit_way_id[2];
  assign N210 = N202 & N205;
  assign N211 = N202 & tag_hit_way_id[2];
  assign N212 = N204 & N205;
  assign N213 = N204 & tag_hit_way_id[2];
  assign aunlock_hit = decode_v_r[6] & N215;
  assign miss_v = N1356 & N1361;
  assign N1356 = N1355 & v_v_r;
  assign N1355 = ~decode_v_r[14];
  assign N1361 = N1360 | aunlock_hit;
  assign N1360 = N1359 | alock_miss;
  assign N1359 = N1358 | aflinv_hit;
  assign N1358 = N1357 | tagfl_hit;
  assign N1357 = ld_st_amo_tag_miss | track_miss;
  assign retval_op_v = N1363 | decode_v_r[4];
  assign N1363 = N1362 | decode_v_r[11];
  assign N1362 = decode_v_r[16] | decode_v_r[12];
  assign _1_net_ = v_o & yumi_i;
  assign N216 = ~sbuf_way_decode[0];
  assign N217 = sbuf_expand_mask[15] & sbuf_entry_lo[18];
  assign N218 = sbuf_expand_mask[14] & sbuf_entry_lo[17];
  assign N219 = sbuf_expand_mask[13] & sbuf_entry_lo[16];
  assign N220 = sbuf_expand_mask[12] & sbuf_entry_lo[15];
  assign N221 = sbuf_expand_mask[11] & sbuf_entry_lo[14];
  assign N222 = sbuf_expand_mask[10] & sbuf_entry_lo[13];
  assign N223 = sbuf_expand_mask[9] & sbuf_entry_lo[12];
  assign N224 = sbuf_expand_mask[8] & sbuf_entry_lo[11];
  assign N225 = sbuf_expand_mask[7] & sbuf_entry_lo[10];
  assign N226 = sbuf_expand_mask[6] & sbuf_entry_lo[9];
  assign N227 = sbuf_expand_mask[5] & sbuf_entry_lo[8];
  assign N228 = sbuf_expand_mask[4] & sbuf_entry_lo[7];
  assign N229 = sbuf_expand_mask[3] & sbuf_entry_lo[6];
  assign N230 = sbuf_expand_mask[2] & sbuf_entry_lo[5];
  assign N231 = sbuf_expand_mask[1] & sbuf_entry_lo[4];
  assign N232 = sbuf_expand_mask[0] & sbuf_entry_lo[3];
  assign N233 = ~sbuf_way_decode[1];
  assign N234 = sbuf_expand_mask[15] & sbuf_entry_lo[18];
  assign N235 = sbuf_expand_mask[14] & sbuf_entry_lo[17];
  assign N236 = sbuf_expand_mask[13] & sbuf_entry_lo[16];
  assign N237 = sbuf_expand_mask[12] & sbuf_entry_lo[15];
  assign N238 = sbuf_expand_mask[11] & sbuf_entry_lo[14];
  assign N239 = sbuf_expand_mask[10] & sbuf_entry_lo[13];
  assign N240 = sbuf_expand_mask[9] & sbuf_entry_lo[12];
  assign N241 = sbuf_expand_mask[8] & sbuf_entry_lo[11];
  assign N242 = sbuf_expand_mask[7] & sbuf_entry_lo[10];
  assign N243 = sbuf_expand_mask[6] & sbuf_entry_lo[9];
  assign N244 = sbuf_expand_mask[5] & sbuf_entry_lo[8];
  assign N245 = sbuf_expand_mask[4] & sbuf_entry_lo[7];
  assign N246 = sbuf_expand_mask[3] & sbuf_entry_lo[6];
  assign N247 = sbuf_expand_mask[2] & sbuf_entry_lo[5];
  assign N248 = sbuf_expand_mask[1] & sbuf_entry_lo[4];
  assign N249 = sbuf_expand_mask[0] & sbuf_entry_lo[3];
  assign N250 = ~sbuf_way_decode[2];
  assign N251 = sbuf_expand_mask[15] & sbuf_entry_lo[18];
  assign N252 = sbuf_expand_mask[14] & sbuf_entry_lo[17];
  assign N253 = sbuf_expand_mask[13] & sbuf_entry_lo[16];
  assign N254 = sbuf_expand_mask[12] & sbuf_entry_lo[15];
  assign N255 = sbuf_expand_mask[11] & sbuf_entry_lo[14];
  assign N256 = sbuf_expand_mask[10] & sbuf_entry_lo[13];
  assign N257 = sbuf_expand_mask[9] & sbuf_entry_lo[12];
  assign N258 = sbuf_expand_mask[8] & sbuf_entry_lo[11];
  assign N259 = sbuf_expand_mask[7] & sbuf_entry_lo[10];
  assign N260 = sbuf_expand_mask[6] & sbuf_entry_lo[9];
  assign N261 = sbuf_expand_mask[5] & sbuf_entry_lo[8];
  assign N262 = sbuf_expand_mask[4] & sbuf_entry_lo[7];
  assign N263 = sbuf_expand_mask[3] & sbuf_entry_lo[6];
  assign N264 = sbuf_expand_mask[2] & sbuf_entry_lo[5];
  assign N265 = sbuf_expand_mask[1] & sbuf_entry_lo[4];
  assign N266 = sbuf_expand_mask[0] & sbuf_entry_lo[3];
  assign N267 = ~sbuf_way_decode[3];
  assign N268 = sbuf_expand_mask[15] & sbuf_entry_lo[18];
  assign N269 = sbuf_expand_mask[14] & sbuf_entry_lo[17];
  assign N270 = sbuf_expand_mask[13] & sbuf_entry_lo[16];
  assign N271 = sbuf_expand_mask[12] & sbuf_entry_lo[15];
  assign N272 = sbuf_expand_mask[11] & sbuf_entry_lo[14];
  assign N273 = sbuf_expand_mask[10] & sbuf_entry_lo[13];
  assign N274 = sbuf_expand_mask[9] & sbuf_entry_lo[12];
  assign N275 = sbuf_expand_mask[8] & sbuf_entry_lo[11];
  assign N276 = sbuf_expand_mask[7] & sbuf_entry_lo[10];
  assign N277 = sbuf_expand_mask[6] & sbuf_entry_lo[9];
  assign N278 = sbuf_expand_mask[5] & sbuf_entry_lo[8];
  assign N279 = sbuf_expand_mask[4] & sbuf_entry_lo[7];
  assign N280 = sbuf_expand_mask[3] & sbuf_entry_lo[6];
  assign N281 = sbuf_expand_mask[2] & sbuf_entry_lo[5];
  assign N282 = sbuf_expand_mask[1] & sbuf_entry_lo[4];
  assign N283 = sbuf_expand_mask[0] & sbuf_entry_lo[3];
  assign N284 = ~sbuf_way_decode[4];
  assign N285 = sbuf_expand_mask[15] & sbuf_entry_lo[18];
  assign N286 = sbuf_expand_mask[14] & sbuf_entry_lo[17];
  assign N287 = sbuf_expand_mask[13] & sbuf_entry_lo[16];
  assign N288 = sbuf_expand_mask[12] & sbuf_entry_lo[15];
  assign N289 = sbuf_expand_mask[11] & sbuf_entry_lo[14];
  assign N290 = sbuf_expand_mask[10] & sbuf_entry_lo[13];
  assign N291 = sbuf_expand_mask[9] & sbuf_entry_lo[12];
  assign N292 = sbuf_expand_mask[8] & sbuf_entry_lo[11];
  assign N293 = sbuf_expand_mask[7] & sbuf_entry_lo[10];
  assign N294 = sbuf_expand_mask[6] & sbuf_entry_lo[9];
  assign N295 = sbuf_expand_mask[5] & sbuf_entry_lo[8];
  assign N296 = sbuf_expand_mask[4] & sbuf_entry_lo[7];
  assign N297 = sbuf_expand_mask[3] & sbuf_entry_lo[6];
  assign N298 = sbuf_expand_mask[2] & sbuf_entry_lo[5];
  assign N299 = sbuf_expand_mask[1] & sbuf_entry_lo[4];
  assign N300 = sbuf_expand_mask[0] & sbuf_entry_lo[3];
  assign N301 = ~sbuf_way_decode[5];
  assign N302 = sbuf_expand_mask[15] & sbuf_entry_lo[18];
  assign N303 = sbuf_expand_mask[14] & sbuf_entry_lo[17];
  assign N304 = sbuf_expand_mask[13] & sbuf_entry_lo[16];
  assign N305 = sbuf_expand_mask[12] & sbuf_entry_lo[15];
  assign N306 = sbuf_expand_mask[11] & sbuf_entry_lo[14];
  assign N307 = sbuf_expand_mask[10] & sbuf_entry_lo[13];
  assign N308 = sbuf_expand_mask[9] & sbuf_entry_lo[12];
  assign N309 = sbuf_expand_mask[8] & sbuf_entry_lo[11];
  assign N310 = sbuf_expand_mask[7] & sbuf_entry_lo[10];
  assign N311 = sbuf_expand_mask[6] & sbuf_entry_lo[9];
  assign N312 = sbuf_expand_mask[5] & sbuf_entry_lo[8];
  assign N313 = sbuf_expand_mask[4] & sbuf_entry_lo[7];
  assign N314 = sbuf_expand_mask[3] & sbuf_entry_lo[6];
  assign N315 = sbuf_expand_mask[2] & sbuf_entry_lo[5];
  assign N316 = sbuf_expand_mask[1] & sbuf_entry_lo[4];
  assign N317 = sbuf_expand_mask[0] & sbuf_entry_lo[3];
  assign N318 = ~sbuf_way_decode[6];
  assign N319 = sbuf_expand_mask[15] & sbuf_entry_lo[18];
  assign N320 = sbuf_expand_mask[14] & sbuf_entry_lo[17];
  assign N321 = sbuf_expand_mask[13] & sbuf_entry_lo[16];
  assign N322 = sbuf_expand_mask[12] & sbuf_entry_lo[15];
  assign N323 = sbuf_expand_mask[11] & sbuf_entry_lo[14];
  assign N324 = sbuf_expand_mask[10] & sbuf_entry_lo[13];
  assign N325 = sbuf_expand_mask[9] & sbuf_entry_lo[12];
  assign N326 = sbuf_expand_mask[8] & sbuf_entry_lo[11];
  assign N327 = sbuf_expand_mask[7] & sbuf_entry_lo[10];
  assign N328 = sbuf_expand_mask[6] & sbuf_entry_lo[9];
  assign N329 = sbuf_expand_mask[5] & sbuf_entry_lo[8];
  assign N330 = sbuf_expand_mask[4] & sbuf_entry_lo[7];
  assign N331 = sbuf_expand_mask[3] & sbuf_entry_lo[6];
  assign N332 = sbuf_expand_mask[2] & sbuf_entry_lo[5];
  assign N333 = sbuf_expand_mask[1] & sbuf_entry_lo[4];
  assign N334 = sbuf_expand_mask[0] & sbuf_entry_lo[3];
  assign N335 = ~sbuf_way_decode[7];
  assign N336 = sbuf_expand_mask[15] & sbuf_entry_lo[18];
  assign N337 = sbuf_expand_mask[14] & sbuf_entry_lo[17];
  assign N338 = sbuf_expand_mask[13] & sbuf_entry_lo[16];
  assign N339 = sbuf_expand_mask[12] & sbuf_entry_lo[15];
  assign N340 = sbuf_expand_mask[11] & sbuf_entry_lo[14];
  assign N341 = sbuf_expand_mask[10] & sbuf_entry_lo[13];
  assign N342 = sbuf_expand_mask[9] & sbuf_entry_lo[12];
  assign N343 = sbuf_expand_mask[8] & sbuf_entry_lo[11];
  assign N344 = sbuf_expand_mask[7] & sbuf_entry_lo[10];
  assign N345 = sbuf_expand_mask[6] & sbuf_entry_lo[9];
  assign N346 = sbuf_expand_mask[5] & sbuf_entry_lo[8];
  assign N347 = sbuf_expand_mask[4] & sbuf_entry_lo[7];
  assign N348 = sbuf_expand_mask[3] & sbuf_entry_lo[6];
  assign N349 = sbuf_expand_mask[2] & sbuf_entry_lo[5];
  assign N350 = sbuf_expand_mask[1] & sbuf_entry_lo[4];
  assign N351 = sbuf_expand_mask[0] & sbuf_entry_lo[3];
  assign N352 = decode_v_r[19];
  assign N353 = ~N352;
  assign N354 = decode_v_r[19];
  assign N355 = ~N354;
  assign N357 = ~N356;
  assign N362 = ~N361;
  assign N363 = ~decode_v_r[1];
  assign N364 = ~decode_v_r[0];
  assign N369 = ~N368;
  assign N370 = ~decode_v_r[2];
  assign N375 = ~N374;
  assign N376 = ~decode_v_r[1];
  assign N381 = ~N380;
  assign N382 = ~decode_v_r[0];
  assign N387 = ~N386;
  assign N388 = ~decode_v_r[2];
  assign N389 = ~decode_v_r[0];
  assign N394 = ~N393;
  assign N395 = ~decode_v_r[2];
  assign N396 = ~decode_v_r[1];
  assign N401 = ~N400;
  assign N402 = ~decode_v_r[2];
  assign N403 = ~decode_v_r[1];
  assign N404 = ~decode_v_r[0];
  assign N409 = ~N408;
  assign N410 = ~decode_v_r[3];
  assign N415 = ~N414;
  assign N422 = N417 | N1364;
  assign N1364 = N419 | N421;
  assign N423 = atomic_reg_data[63] & atomic_mem_data[63];
  assign N424 = atomic_reg_data[62] & atomic_mem_data[62];
  assign N425 = atomic_reg_data[61] & atomic_mem_data[61];
  assign N426 = atomic_reg_data[60] & atomic_mem_data[60];
  assign N427 = atomic_reg_data[59] & atomic_mem_data[59];
  assign N428 = atomic_reg_data[58] & atomic_mem_data[58];
  assign N429 = atomic_reg_data[57] & atomic_mem_data[57];
  assign N430 = atomic_reg_data[56] & atomic_mem_data[56];
  assign N431 = atomic_reg_data[55] & atomic_mem_data[55];
  assign N432 = atomic_reg_data[54] & atomic_mem_data[54];
  assign N433 = atomic_reg_data[53] & atomic_mem_data[53];
  assign N434 = atomic_reg_data[52] & atomic_mem_data[52];
  assign N435 = atomic_reg_data[51] & atomic_mem_data[51];
  assign N436 = atomic_reg_data[50] & atomic_mem_data[50];
  assign N437 = atomic_reg_data[49] & atomic_mem_data[49];
  assign N438 = atomic_reg_data[48] & atomic_mem_data[48];
  assign N439 = atomic_reg_data[47] & atomic_mem_data[47];
  assign N440 = atomic_reg_data[46] & atomic_mem_data[46];
  assign N441 = atomic_reg_data[45] & atomic_mem_data[45];
  assign N442 = atomic_reg_data[44] & atomic_mem_data[44];
  assign N443 = atomic_reg_data[43] & atomic_mem_data[43];
  assign N444 = atomic_reg_data[42] & atomic_mem_data[42];
  assign N445 = atomic_reg_data[41] & atomic_mem_data[41];
  assign N446 = atomic_reg_data[40] & atomic_mem_data[40];
  assign N447 = atomic_reg_data[39] & atomic_mem_data[39];
  assign N448 = atomic_reg_data[38] & atomic_mem_data[38];
  assign N449 = atomic_reg_data[37] & atomic_mem_data[37];
  assign N450 = atomic_reg_data[36] & atomic_mem_data[36];
  assign N451 = atomic_reg_data[35] & atomic_mem_data[35];
  assign N452 = atomic_reg_data[34] & atomic_mem_data[34];
  assign N453 = atomic_reg_data[33] & atomic_mem_data[33];
  assign N454 = atomic_reg_data[32] & atomic_mem_data[32];
  assign N455 = atomic_reg_data[31] & atomic_mem_data[31];
  assign N456 = atomic_reg_data[30] & atomic_mem_data[30];
  assign N457 = atomic_reg_data[29] & atomic_mem_data[29];
  assign N458 = atomic_reg_data[28] & atomic_mem_data[28];
  assign N459 = atomic_reg_data[27] & atomic_mem_data[27];
  assign N460 = atomic_reg_data[26] & atomic_mem_data[26];
  assign N461 = atomic_reg_data[25] & atomic_mem_data[25];
  assign N462 = atomic_reg_data[24] & atomic_mem_data[24];
  assign N463 = atomic_reg_data[23] & atomic_mem_data[23];
  assign N464 = atomic_reg_data[22] & atomic_mem_data[22];
  assign N465 = atomic_reg_data[21] & atomic_mem_data[21];
  assign N466 = atomic_reg_data[20] & atomic_mem_data[20];
  assign N467 = atomic_reg_data[19] & atomic_mem_data[19];
  assign N468 = atomic_reg_data[18] & atomic_mem_data[18];
  assign N469 = atomic_reg_data[17] & atomic_mem_data[17];
  assign N470 = atomic_reg_data[16] & atomic_mem_data[16];
  assign N471 = atomic_reg_data[15] & atomic_mem_data[15];
  assign N472 = atomic_reg_data[14] & atomic_mem_data[14];
  assign N473 = atomic_reg_data[13] & atomic_mem_data[13];
  assign N474 = atomic_reg_data[12] & atomic_mem_data[12];
  assign N475 = atomic_reg_data[11] & atomic_mem_data[11];
  assign N476 = atomic_reg_data[10] & atomic_mem_data[10];
  assign N477 = atomic_reg_data[9] & atomic_mem_data[9];
  assign N478 = atomic_reg_data[8] & atomic_mem_data[8];
  assign N479 = atomic_reg_data[7] & atomic_mem_data[7];
  assign N480 = atomic_reg_data[6] & atomic_mem_data[6];
  assign N481 = atomic_reg_data[5] & atomic_mem_data[5];
  assign N482 = atomic_reg_data[4] & atomic_mem_data[4];
  assign N483 = atomic_reg_data[3] & atomic_mem_data[3];
  assign N484 = atomic_reg_data[2] & atomic_mem_data[2];
  assign N485 = atomic_reg_data[1] & atomic_mem_data[1];
  assign N486 = atomic_reg_data[0] & atomic_mem_data[0];
  assign N487 = atomic_reg_data[63] | atomic_mem_data[63];
  assign N488 = atomic_reg_data[62] | atomic_mem_data[62];
  assign N489 = atomic_reg_data[61] | atomic_mem_data[61];
  assign N490 = atomic_reg_data[60] | atomic_mem_data[60];
  assign N491 = atomic_reg_data[59] | atomic_mem_data[59];
  assign N492 = atomic_reg_data[58] | atomic_mem_data[58];
  assign N493 = atomic_reg_data[57] | atomic_mem_data[57];
  assign N494 = atomic_reg_data[56] | atomic_mem_data[56];
  assign N495 = atomic_reg_data[55] | atomic_mem_data[55];
  assign N496 = atomic_reg_data[54] | atomic_mem_data[54];
  assign N497 = atomic_reg_data[53] | atomic_mem_data[53];
  assign N498 = atomic_reg_data[52] | atomic_mem_data[52];
  assign N499 = atomic_reg_data[51] | atomic_mem_data[51];
  assign N500 = atomic_reg_data[50] | atomic_mem_data[50];
  assign N501 = atomic_reg_data[49] | atomic_mem_data[49];
  assign N502 = atomic_reg_data[48] | atomic_mem_data[48];
  assign N503 = atomic_reg_data[47] | atomic_mem_data[47];
  assign N504 = atomic_reg_data[46] | atomic_mem_data[46];
  assign N505 = atomic_reg_data[45] | atomic_mem_data[45];
  assign N506 = atomic_reg_data[44] | atomic_mem_data[44];
  assign N507 = atomic_reg_data[43] | atomic_mem_data[43];
  assign N508 = atomic_reg_data[42] | atomic_mem_data[42];
  assign N509 = atomic_reg_data[41] | atomic_mem_data[41];
  assign N510 = atomic_reg_data[40] | atomic_mem_data[40];
  assign N511 = atomic_reg_data[39] | atomic_mem_data[39];
  assign N512 = atomic_reg_data[38] | atomic_mem_data[38];
  assign N513 = atomic_reg_data[37] | atomic_mem_data[37];
  assign N514 = atomic_reg_data[36] | atomic_mem_data[36];
  assign N515 = atomic_reg_data[35] | atomic_mem_data[35];
  assign N516 = atomic_reg_data[34] | atomic_mem_data[34];
  assign N517 = atomic_reg_data[33] | atomic_mem_data[33];
  assign N518 = atomic_reg_data[32] | atomic_mem_data[32];
  assign N519 = atomic_reg_data[31] | atomic_mem_data[31];
  assign N520 = atomic_reg_data[30] | atomic_mem_data[30];
  assign N521 = atomic_reg_data[29] | atomic_mem_data[29];
  assign N522 = atomic_reg_data[28] | atomic_mem_data[28];
  assign N523 = atomic_reg_data[27] | atomic_mem_data[27];
  assign N524 = atomic_reg_data[26] | atomic_mem_data[26];
  assign N525 = atomic_reg_data[25] | atomic_mem_data[25];
  assign N526 = atomic_reg_data[24] | atomic_mem_data[24];
  assign N527 = atomic_reg_data[23] | atomic_mem_data[23];
  assign N528 = atomic_reg_data[22] | atomic_mem_data[22];
  assign N529 = atomic_reg_data[21] | atomic_mem_data[21];
  assign N530 = atomic_reg_data[20] | atomic_mem_data[20];
  assign N531 = atomic_reg_data[19] | atomic_mem_data[19];
  assign N532 = atomic_reg_data[18] | atomic_mem_data[18];
  assign N533 = atomic_reg_data[17] | atomic_mem_data[17];
  assign N534 = atomic_reg_data[16] | atomic_mem_data[16];
  assign N535 = atomic_reg_data[15] | atomic_mem_data[15];
  assign N536 = atomic_reg_data[14] | atomic_mem_data[14];
  assign N537 = atomic_reg_data[13] | atomic_mem_data[13];
  assign N538 = atomic_reg_data[12] | atomic_mem_data[12];
  assign N539 = atomic_reg_data[11] | atomic_mem_data[11];
  assign N540 = atomic_reg_data[10] | atomic_mem_data[10];
  assign N541 = atomic_reg_data[9] | atomic_mem_data[9];
  assign N542 = atomic_reg_data[8] | atomic_mem_data[8];
  assign N543 = atomic_reg_data[7] | atomic_mem_data[7];
  assign N544 = atomic_reg_data[6] | atomic_mem_data[6];
  assign N545 = atomic_reg_data[5] | atomic_mem_data[5];
  assign N546 = atomic_reg_data[4] | atomic_mem_data[4];
  assign N547 = atomic_reg_data[3] | atomic_mem_data[3];
  assign N548 = atomic_reg_data[2] | atomic_mem_data[2];
  assign N549 = atomic_reg_data[1] | atomic_mem_data[1];
  assign N550 = atomic_reg_data[0] | atomic_mem_data[0];
  assign N551 = atomic_reg_data[63] ^ atomic_mem_data[63];
  assign N552 = atomic_reg_data[62] ^ atomic_mem_data[62];
  assign N553 = atomic_reg_data[61] ^ atomic_mem_data[61];
  assign N554 = atomic_reg_data[60] ^ atomic_mem_data[60];
  assign N555 = atomic_reg_data[59] ^ atomic_mem_data[59];
  assign N556 = atomic_reg_data[58] ^ atomic_mem_data[58];
  assign N557 = atomic_reg_data[57] ^ atomic_mem_data[57];
  assign N558 = atomic_reg_data[56] ^ atomic_mem_data[56];
  assign N559 = atomic_reg_data[55] ^ atomic_mem_data[55];
  assign N560 = atomic_reg_data[54] ^ atomic_mem_data[54];
  assign N561 = atomic_reg_data[53] ^ atomic_mem_data[53];
  assign N562 = atomic_reg_data[52] ^ atomic_mem_data[52];
  assign N563 = atomic_reg_data[51] ^ atomic_mem_data[51];
  assign N564 = atomic_reg_data[50] ^ atomic_mem_data[50];
  assign N565 = atomic_reg_data[49] ^ atomic_mem_data[49];
  assign N566 = atomic_reg_data[48] ^ atomic_mem_data[48];
  assign N567 = atomic_reg_data[47] ^ atomic_mem_data[47];
  assign N568 = atomic_reg_data[46] ^ atomic_mem_data[46];
  assign N569 = atomic_reg_data[45] ^ atomic_mem_data[45];
  assign N570 = atomic_reg_data[44] ^ atomic_mem_data[44];
  assign N571 = atomic_reg_data[43] ^ atomic_mem_data[43];
  assign N572 = atomic_reg_data[42] ^ atomic_mem_data[42];
  assign N573 = atomic_reg_data[41] ^ atomic_mem_data[41];
  assign N574 = atomic_reg_data[40] ^ atomic_mem_data[40];
  assign N575 = atomic_reg_data[39] ^ atomic_mem_data[39];
  assign N576 = atomic_reg_data[38] ^ atomic_mem_data[38];
  assign N577 = atomic_reg_data[37] ^ atomic_mem_data[37];
  assign N578 = atomic_reg_data[36] ^ atomic_mem_data[36];
  assign N579 = atomic_reg_data[35] ^ atomic_mem_data[35];
  assign N580 = atomic_reg_data[34] ^ atomic_mem_data[34];
  assign N581 = atomic_reg_data[33] ^ atomic_mem_data[33];
  assign N582 = atomic_reg_data[32] ^ atomic_mem_data[32];
  assign N583 = atomic_reg_data[31] ^ atomic_mem_data[31];
  assign N584 = atomic_reg_data[30] ^ atomic_mem_data[30];
  assign N585 = atomic_reg_data[29] ^ atomic_mem_data[29];
  assign N586 = atomic_reg_data[28] ^ atomic_mem_data[28];
  assign N587 = atomic_reg_data[27] ^ atomic_mem_data[27];
  assign N588 = atomic_reg_data[26] ^ atomic_mem_data[26];
  assign N589 = atomic_reg_data[25] ^ atomic_mem_data[25];
  assign N590 = atomic_reg_data[24] ^ atomic_mem_data[24];
  assign N591 = atomic_reg_data[23] ^ atomic_mem_data[23];
  assign N592 = atomic_reg_data[22] ^ atomic_mem_data[22];
  assign N593 = atomic_reg_data[21] ^ atomic_mem_data[21];
  assign N594 = atomic_reg_data[20] ^ atomic_mem_data[20];
  assign N595 = atomic_reg_data[19] ^ atomic_mem_data[19];
  assign N596 = atomic_reg_data[18] ^ atomic_mem_data[18];
  assign N597 = atomic_reg_data[17] ^ atomic_mem_data[17];
  assign N598 = atomic_reg_data[16] ^ atomic_mem_data[16];
  assign N599 = atomic_reg_data[15] ^ atomic_mem_data[15];
  assign N600 = atomic_reg_data[14] ^ atomic_mem_data[14];
  assign N601 = atomic_reg_data[13] ^ atomic_mem_data[13];
  assign N602 = atomic_reg_data[12] ^ atomic_mem_data[12];
  assign N603 = atomic_reg_data[11] ^ atomic_mem_data[11];
  assign N604 = atomic_reg_data[10] ^ atomic_mem_data[10];
  assign N605 = atomic_reg_data[9] ^ atomic_mem_data[9];
  assign N606 = atomic_reg_data[8] ^ atomic_mem_data[8];
  assign N607 = atomic_reg_data[7] ^ atomic_mem_data[7];
  assign N608 = atomic_reg_data[6] ^ atomic_mem_data[6];
  assign N609 = atomic_reg_data[5] ^ atomic_mem_data[5];
  assign N610 = atomic_reg_data[4] ^ atomic_mem_data[4];
  assign N611 = atomic_reg_data[3] ^ atomic_mem_data[3];
  assign N612 = atomic_reg_data[2] ^ atomic_mem_data[2];
  assign N613 = atomic_reg_data[1] ^ atomic_mem_data[1];
  assign N614 = atomic_reg_data[0] ^ atomic_mem_data[0];
  assign N680 = ~N679;
  assign N746 = ~N745;
  assign N812 = ~N811;
  assign N878 = ~N877;
  assign N943 = decode_v_r[19];
  assign N944 = ~N943;
  assign N945 = decode_v_r[4];
  assign N946 = ~N945;
  assign N947 = decode_v_r[4];
  assign N948 = ~N947;
  assign N949 = decode_v_r[17];
  assign N950 = ~N949;
  assign N951 = ~tbuf_way_decode[0];
  assign N952 = ~tbuf_way_decode[1];
  assign N953 = ~tbuf_way_decode[2];
  assign N954 = ~tbuf_way_decode[3];
  assign N955 = ~tbuf_way_decode[4];
  assign N956 = ~tbuf_way_decode[5];
  assign N957 = ~tbuf_way_decode[6];
  assign N958 = ~tbuf_way_decode[7];
  assign N959 = ~select_snoop_data_r_lo;
  assign ld_data_masked[127] = snoop_or_ld_data[127] & expanded_mask_v[127];
  assign ld_data_masked[126] = snoop_or_ld_data[126] & expanded_mask_v[126];
  assign ld_data_masked[125] = snoop_or_ld_data[125] & expanded_mask_v[125];
  assign ld_data_masked[124] = snoop_or_ld_data[124] & expanded_mask_v[124];
  assign ld_data_masked[123] = snoop_or_ld_data[123] & expanded_mask_v[123];
  assign ld_data_masked[122] = snoop_or_ld_data[122] & expanded_mask_v[122];
  assign ld_data_masked[121] = snoop_or_ld_data[121] & expanded_mask_v[121];
  assign ld_data_masked[120] = snoop_or_ld_data[120] & expanded_mask_v[120];
  assign ld_data_masked[119] = snoop_or_ld_data[119] & expanded_mask_v[119];
  assign ld_data_masked[118] = snoop_or_ld_data[118] & expanded_mask_v[118];
  assign ld_data_masked[117] = snoop_or_ld_data[117] & expanded_mask_v[117];
  assign ld_data_masked[116] = snoop_or_ld_data[116] & expanded_mask_v[116];
  assign ld_data_masked[115] = snoop_or_ld_data[115] & expanded_mask_v[115];
  assign ld_data_masked[114] = snoop_or_ld_data[114] & expanded_mask_v[114];
  assign ld_data_masked[113] = snoop_or_ld_data[113] & expanded_mask_v[113];
  assign ld_data_masked[112] = snoop_or_ld_data[112] & expanded_mask_v[112];
  assign ld_data_masked[111] = snoop_or_ld_data[111] & expanded_mask_v[111];
  assign ld_data_masked[110] = snoop_or_ld_data[110] & expanded_mask_v[110];
  assign ld_data_masked[109] = snoop_or_ld_data[109] & expanded_mask_v[109];
  assign ld_data_masked[108] = snoop_or_ld_data[108] & expanded_mask_v[108];
  assign ld_data_masked[107] = snoop_or_ld_data[107] & expanded_mask_v[107];
  assign ld_data_masked[106] = snoop_or_ld_data[106] & expanded_mask_v[106];
  assign ld_data_masked[105] = snoop_or_ld_data[105] & expanded_mask_v[105];
  assign ld_data_masked[104] = snoop_or_ld_data[104] & expanded_mask_v[104];
  assign ld_data_masked[103] = snoop_or_ld_data[103] & expanded_mask_v[103];
  assign ld_data_masked[102] = snoop_or_ld_data[102] & expanded_mask_v[102];
  assign ld_data_masked[101] = snoop_or_ld_data[101] & expanded_mask_v[101];
  assign ld_data_masked[100] = snoop_or_ld_data[100] & expanded_mask_v[100];
  assign ld_data_masked[99] = snoop_or_ld_data[99] & expanded_mask_v[99];
  assign ld_data_masked[98] = snoop_or_ld_data[98] & expanded_mask_v[98];
  assign ld_data_masked[97] = snoop_or_ld_data[97] & expanded_mask_v[97];
  assign ld_data_masked[96] = snoop_or_ld_data[96] & expanded_mask_v[96];
  assign ld_data_masked[95] = snoop_or_ld_data[95] & expanded_mask_v[95];
  assign ld_data_masked[94] = snoop_or_ld_data[94] & expanded_mask_v[94];
  assign ld_data_masked[93] = snoop_or_ld_data[93] & expanded_mask_v[93];
  assign ld_data_masked[92] = snoop_or_ld_data[92] & expanded_mask_v[92];
  assign ld_data_masked[91] = snoop_or_ld_data[91] & expanded_mask_v[91];
  assign ld_data_masked[90] = snoop_or_ld_data[90] & expanded_mask_v[90];
  assign ld_data_masked[89] = snoop_or_ld_data[89] & expanded_mask_v[89];
  assign ld_data_masked[88] = snoop_or_ld_data[88] & expanded_mask_v[88];
  assign ld_data_masked[87] = snoop_or_ld_data[87] & expanded_mask_v[87];
  assign ld_data_masked[86] = snoop_or_ld_data[86] & expanded_mask_v[86];
  assign ld_data_masked[85] = snoop_or_ld_data[85] & expanded_mask_v[85];
  assign ld_data_masked[84] = snoop_or_ld_data[84] & expanded_mask_v[84];
  assign ld_data_masked[83] = snoop_or_ld_data[83] & expanded_mask_v[83];
  assign ld_data_masked[82] = snoop_or_ld_data[82] & expanded_mask_v[82];
  assign ld_data_masked[81] = snoop_or_ld_data[81] & expanded_mask_v[81];
  assign ld_data_masked[80] = snoop_or_ld_data[80] & expanded_mask_v[80];
  assign ld_data_masked[79] = snoop_or_ld_data[79] & expanded_mask_v[79];
  assign ld_data_masked[78] = snoop_or_ld_data[78] & expanded_mask_v[78];
  assign ld_data_masked[77] = snoop_or_ld_data[77] & expanded_mask_v[77];
  assign ld_data_masked[76] = snoop_or_ld_data[76] & expanded_mask_v[76];
  assign ld_data_masked[75] = snoop_or_ld_data[75] & expanded_mask_v[75];
  assign ld_data_masked[74] = snoop_or_ld_data[74] & expanded_mask_v[74];
  assign ld_data_masked[73] = snoop_or_ld_data[73] & expanded_mask_v[73];
  assign ld_data_masked[72] = snoop_or_ld_data[72] & expanded_mask_v[72];
  assign ld_data_masked[71] = snoop_or_ld_data[71] & expanded_mask_v[71];
  assign ld_data_masked[70] = snoop_or_ld_data[70] & expanded_mask_v[70];
  assign ld_data_masked[69] = snoop_or_ld_data[69] & expanded_mask_v[69];
  assign ld_data_masked[68] = snoop_or_ld_data[68] & expanded_mask_v[68];
  assign ld_data_masked[67] = snoop_or_ld_data[67] & expanded_mask_v[67];
  assign ld_data_masked[66] = snoop_or_ld_data[66] & expanded_mask_v[66];
  assign ld_data_masked[65] = snoop_or_ld_data[65] & expanded_mask_v[65];
  assign ld_data_masked[64] = snoop_or_ld_data[64] & expanded_mask_v[64];
  assign ld_data_masked[63] = snoop_or_ld_data[63] & expanded_mask_v[63];
  assign ld_data_masked[62] = snoop_or_ld_data[62] & expanded_mask_v[62];
  assign ld_data_masked[61] = snoop_or_ld_data[61] & expanded_mask_v[61];
  assign ld_data_masked[60] = snoop_or_ld_data[60] & expanded_mask_v[60];
  assign ld_data_masked[59] = snoop_or_ld_data[59] & expanded_mask_v[59];
  assign ld_data_masked[58] = snoop_or_ld_data[58] & expanded_mask_v[58];
  assign ld_data_masked[57] = snoop_or_ld_data[57] & expanded_mask_v[57];
  assign ld_data_masked[56] = snoop_or_ld_data[56] & expanded_mask_v[56];
  assign ld_data_masked[55] = snoop_or_ld_data[55] & expanded_mask_v[55];
  assign ld_data_masked[54] = snoop_or_ld_data[54] & expanded_mask_v[54];
  assign ld_data_masked[53] = snoop_or_ld_data[53] & expanded_mask_v[53];
  assign ld_data_masked[52] = snoop_or_ld_data[52] & expanded_mask_v[52];
  assign ld_data_masked[51] = snoop_or_ld_data[51] & expanded_mask_v[51];
  assign ld_data_masked[50] = snoop_or_ld_data[50] & expanded_mask_v[50];
  assign ld_data_masked[49] = snoop_or_ld_data[49] & expanded_mask_v[49];
  assign ld_data_masked[48] = snoop_or_ld_data[48] & expanded_mask_v[48];
  assign ld_data_masked[47] = snoop_or_ld_data[47] & expanded_mask_v[47];
  assign ld_data_masked[46] = snoop_or_ld_data[46] & expanded_mask_v[46];
  assign ld_data_masked[45] = snoop_or_ld_data[45] & expanded_mask_v[45];
  assign ld_data_masked[44] = snoop_or_ld_data[44] & expanded_mask_v[44];
  assign ld_data_masked[43] = snoop_or_ld_data[43] & expanded_mask_v[43];
  assign ld_data_masked[42] = snoop_or_ld_data[42] & expanded_mask_v[42];
  assign ld_data_masked[41] = snoop_or_ld_data[41] & expanded_mask_v[41];
  assign ld_data_masked[40] = snoop_or_ld_data[40] & expanded_mask_v[40];
  assign ld_data_masked[39] = snoop_or_ld_data[39] & expanded_mask_v[39];
  assign ld_data_masked[38] = snoop_or_ld_data[38] & expanded_mask_v[38];
  assign ld_data_masked[37] = snoop_or_ld_data[37] & expanded_mask_v[37];
  assign ld_data_masked[36] = snoop_or_ld_data[36] & expanded_mask_v[36];
  assign ld_data_masked[35] = snoop_or_ld_data[35] & expanded_mask_v[35];
  assign ld_data_masked[34] = snoop_or_ld_data[34] & expanded_mask_v[34];
  assign ld_data_masked[33] = snoop_or_ld_data[33] & expanded_mask_v[33];
  assign ld_data_masked[32] = snoop_or_ld_data[32] & expanded_mask_v[32];
  assign ld_data_masked[31] = snoop_or_ld_data[31] & expanded_mask_v[31];
  assign ld_data_masked[30] = snoop_or_ld_data[30] & expanded_mask_v[30];
  assign ld_data_masked[29] = snoop_or_ld_data[29] & expanded_mask_v[29];
  assign ld_data_masked[28] = snoop_or_ld_data[28] & expanded_mask_v[28];
  assign ld_data_masked[27] = snoop_or_ld_data[27] & expanded_mask_v[27];
  assign ld_data_masked[26] = snoop_or_ld_data[26] & expanded_mask_v[26];
  assign ld_data_masked[25] = snoop_or_ld_data[25] & expanded_mask_v[25];
  assign ld_data_masked[24] = snoop_or_ld_data[24] & expanded_mask_v[24];
  assign ld_data_masked[23] = snoop_or_ld_data[23] & expanded_mask_v[23];
  assign ld_data_masked[22] = snoop_or_ld_data[22] & expanded_mask_v[22];
  assign ld_data_masked[21] = snoop_or_ld_data[21] & expanded_mask_v[21];
  assign ld_data_masked[20] = snoop_or_ld_data[20] & expanded_mask_v[20];
  assign ld_data_masked[19] = snoop_or_ld_data[19] & expanded_mask_v[19];
  assign ld_data_masked[18] = snoop_or_ld_data[18] & expanded_mask_v[18];
  assign ld_data_masked[17] = snoop_or_ld_data[17] & expanded_mask_v[17];
  assign ld_data_masked[16] = snoop_or_ld_data[16] & expanded_mask_v[16];
  assign ld_data_masked[15] = snoop_or_ld_data[15] & expanded_mask_v[15];
  assign ld_data_masked[14] = snoop_or_ld_data[14] & expanded_mask_v[14];
  assign ld_data_masked[13] = snoop_or_ld_data[13] & expanded_mask_v[13];
  assign ld_data_masked[12] = snoop_or_ld_data[12] & expanded_mask_v[12];
  assign ld_data_masked[11] = snoop_or_ld_data[11] & expanded_mask_v[11];
  assign ld_data_masked[10] = snoop_or_ld_data[10] & expanded_mask_v[10];
  assign ld_data_masked[9] = snoop_or_ld_data[9] & expanded_mask_v[9];
  assign ld_data_masked[8] = snoop_or_ld_data[8] & expanded_mask_v[8];
  assign ld_data_masked[7] = snoop_or_ld_data[7] & expanded_mask_v[7];
  assign ld_data_masked[6] = snoop_or_ld_data[6] & expanded_mask_v[6];
  assign ld_data_masked[5] = snoop_or_ld_data[5] & expanded_mask_v[5];
  assign ld_data_masked[4] = snoop_or_ld_data[4] & expanded_mask_v[4];
  assign ld_data_masked[3] = snoop_or_ld_data[3] & expanded_mask_v[3];
  assign ld_data_masked[2] = snoop_or_ld_data[2] & expanded_mask_v[2];
  assign ld_data_masked[1] = snoop_or_ld_data[1] & expanded_mask_v[1];
  assign ld_data_masked[0] = snoop_or_ld_data[0] & expanded_mask_v[0];
  assign ld_data_final_li_0__127_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__126_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__125_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__124_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__123_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__122_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__121_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__120_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__119_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__118_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__117_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__116_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__115_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__114_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__113_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__112_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__111_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__110_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__109_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__108_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__107_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__106_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__105_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__104_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__103_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__102_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__101_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__100_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__99_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__98_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__97_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__96_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__95_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__94_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__93_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__92_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__91_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__90_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__89_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__88_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__87_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__86_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__85_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__84_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__83_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__82_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__81_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__80_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__79_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__78_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__77_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__76_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__75_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__74_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__73_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__72_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__71_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__70_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__69_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__68_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__67_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__66_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__65_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__64_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__63_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__62_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__61_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__60_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__59_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__58_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__57_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__56_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__55_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__54_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__53_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__52_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__51_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__50_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__49_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__48_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__47_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__46_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__45_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__44_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__43_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__42_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__41_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__40_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__39_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__38_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__37_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__36_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__35_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__34_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__33_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__32_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__31_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__30_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__29_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__28_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__27_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__26_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__25_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__24_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__23_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__22_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__21_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__20_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__19_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__18_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__17_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__16_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__15_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__14_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__13_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__12_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__11_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__10_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__9_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__8_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_1__127_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__126_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__125_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__124_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__123_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__122_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__121_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__120_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__119_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__118_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__117_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__116_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__115_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__114_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__113_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__112_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__111_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__110_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__109_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__108_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__107_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__106_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__105_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__104_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__103_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__102_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__101_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__100_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__99_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__98_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__97_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__96_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__95_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__94_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__93_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__92_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__91_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__90_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__89_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__88_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__87_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__86_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__85_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__84_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__83_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__82_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__81_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__80_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__79_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__78_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__77_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__76_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__75_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__74_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__73_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__72_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__71_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__70_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__69_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__68_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__67_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__66_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__65_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__64_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__63_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__62_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__61_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__60_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__59_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__58_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__57_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__56_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__55_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__54_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__53_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__52_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__51_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__50_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__49_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__48_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__47_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__46_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__45_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__44_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__43_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__42_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__41_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__40_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__39_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__38_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__37_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__36_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__35_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__34_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__33_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__32_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__31_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__30_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__29_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__28_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__27_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__26_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__25_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__24_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__23_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__22_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__21_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__20_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__19_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__18_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__17_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__16_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_2__127_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__126_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__125_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__124_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__123_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__122_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__121_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__120_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__119_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__118_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__117_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__116_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__115_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__114_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__113_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__112_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__111_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__110_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__109_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__108_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__107_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__106_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__105_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__104_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__103_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__102_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__101_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__100_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__99_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__98_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__97_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__96_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__95_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__94_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__93_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__92_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__91_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__90_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__89_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__88_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__87_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__86_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__85_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__84_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__83_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__82_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__81_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__80_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__79_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__78_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__77_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__76_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__75_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__74_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__73_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__72_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__71_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__70_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__69_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__68_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__67_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__66_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__65_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__64_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__63_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__62_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__61_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__60_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__59_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__58_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__57_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__56_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__55_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__54_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__53_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__52_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__51_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__50_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__49_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__48_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__47_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__46_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__45_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__44_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__43_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__42_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__41_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__40_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__39_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__38_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__37_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__36_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__35_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__34_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__33_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_2__32_ = decode_v_r[18] & \atomic_64.amo32_mem_in [63];
  assign ld_data_final_li_3__127_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__126_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__125_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__124_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__123_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__122_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__121_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__120_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__119_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__118_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__117_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__116_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__115_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__114_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__113_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__112_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__111_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__110_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__109_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__108_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__107_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__106_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__105_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__104_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__103_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__102_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__101_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__100_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__99_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__98_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__97_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__96_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__95_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__94_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__93_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__92_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__91_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__90_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__89_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__88_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__87_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__86_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__85_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__84_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__83_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__82_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__81_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__80_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__79_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__78_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__77_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__76_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__75_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__74_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__73_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__72_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__71_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__70_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__69_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__68_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__67_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__66_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__65_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign ld_data_final_li_3__64_ = decode_v_r[18] & \atomic_64.amo64_mem_in [63];
  assign N960 = ~retval_op_v;
  assign N961 = decode_v_r[12];
  assign N962 = decode_v_r[11];
  assign N963 = decode_v_r[17];
  assign N964 = N962 | N961;
  assign N965 = N963 | N964;
  assign N966 = ~N965;
  assign N967 = ~addr_v_r[13];
  assign N968 = ~addr_v_r[14];
  assign N969 = N967 & N968;
  assign N970 = N967 & addr_v_r[14];
  assign N971 = addr_v_r[13] & N968;
  assign N972 = addr_v_r[13] & addr_v_r[14];
  assign N973 = ~addr_v_r[15];
  assign N974 = N969 & N973;
  assign N975 = N969 & addr_v_r[15];
  assign N976 = N971 & N973;
  assign N977 = N971 & addr_v_r[15];
  assign N978 = N970 & N973;
  assign N979 = N970 & addr_v_r[15];
  assign N980 = N972 & N973;
  assign N981 = N972 & addr_v_r[15];
  assign N983 = ~addr_v_r[13];
  assign N984 = ~addr_v_r[14];
  assign N985 = N983 & N984;
  assign N986 = N983 & addr_v_r[14];
  assign N987 = addr_v_r[13] & N984;
  assign N988 = addr_v_r[13] & addr_v_r[14];
  assign N989 = ~addr_v_r[15];
  assign N990 = N985 & N989;
  assign N991 = N985 & addr_v_r[15];
  assign N992 = N987 & N989;
  assign N993 = N987 & addr_v_r[15];
  assign N994 = N986 & N989;
  assign N995 = N986 & addr_v_r[15];
  assign N996 = N988 & N989;
  assign N997 = N988 & addr_v_r[15];
  assign N999 = ~addr_v_r[13];
  assign N1000 = ~addr_v_r[14];
  assign N1001 = N999 & N1000;
  assign N1002 = N999 & addr_v_r[14];
  assign N1003 = addr_v_r[13] & N1000;
  assign N1004 = addr_v_r[13] & addr_v_r[14];
  assign N1005 = ~addr_v_r[15];
  assign N1006 = N1001 & N1005;
  assign N1007 = N1001 & addr_v_r[15];
  assign N1008 = N1003 & N1005;
  assign N1009 = N1003 & addr_v_r[15];
  assign N1010 = N1002 & N1005;
  assign N1011 = N1002 & addr_v_r[15];
  assign N1012 = N1004 & N1005;
  assign N1013 = N1004 & addr_v_r[15];
  assign N1162 = ~N961;
  assign N1163 = N962 & N1162;
  assign N1164 = ~N962;
  assign N1165 = N1162 & N1164;
  assign N1166 = N963 & N1165;
  assign N1167 = ~miss_v;
  assign N1168 = miss_v;
  assign v_o = v_v_r & N1169;
  assign N1170 = ~v_v_r;
  assign N1171 = v_o & yumi_i;
  assign sbuf_hazard = N1368 & N1370;
  assign N1368 = sbuf_full_lo & N1367;
  assign N1367 = N1365 & N1366;
  assign N1365 = v_o & yumi_i;
  assign N1366 = decode_v_r[15] | decode_v_r[4];
  assign N1370 = v_i & N1369;
  assign N1369 = decode[16] | decode[4];
  assign N1172 = ~miss_v;
  assign N1173 = miss_v;
  assign N1174 = N1380 & N1381;
  assign N1380 = N1378 & N1379;
  assign N1378 = N1376 & N1377;
  assign N1376 = N1374 & N1375;
  assign N1374 = N1372 & N1373;
  assign N1372 = ~N1371;
  assign N1371 = decode[14] & v_i;
  assign N1373 = ~miss_tag_mem_v_lo;
  assign N1375 = ~miss_track_mem_v_lo;
  assign N1377 = ~dma_data_mem_v_lo;
  assign N1379 = ~recover_lo;
  assign N1381 = ~dma_evict_lo;
  assign tl_ready = N1175 & N1382;
  assign N1382 = ~sbuf_hazard;
  assign N1176 = ~v_tl_r;
  assign tl_we = tl_ready & N1177;
  assign yumi_o = v_i & tl_we;
  assign tagst_write_en = decode[14] & yumi_o;
  assign tag_mem_v_li = N1387 | N1388;
  assign N1387 = N1386 | miss_tag_mem_v_lo;
  assign N1386 = N1383 | N1385;
  assign N1383 = decode[5] & yumi_o;
  assign N1385 = N1384 & v_tl_r;
  assign N1384 = recover_lo & decode_tl_r[5];
  assign N1388 = decode[14] & yumi_o;
  assign N1178 = ~miss_v;
  assign N1179 = miss_v;
  assign N1180 = miss_tag_mem_v_lo & miss_tag_mem_w_lo;
  assign N1181 = ~miss_v;
  assign N1182 = miss_v;
  assign N1183 = miss_tag_mem_v_lo | recover_lo;
  assign N1184 = ~N1183;
  assign N1192 = ~recover_lo;
  assign N1193 = miss_tag_mem_v_lo & N1192;
  assign data_mem_v_li = N1395 | N1396;
  assign N1395 = N1394 | dma_data_mem_v_lo;
  assign N1394 = N1390 | N1393;
  assign N1390 = yumi_o & N1389;
  assign N1389 = decode[16] | decode[4];
  assign N1393 = N1391 & N1392;
  assign N1391 = v_tl_r & recover_lo;
  assign N1392 = decode_tl_r[16] | decode_tl_r[4];
  assign N1396 = sbuf_v_lo & sbuf_yumi_li;
  assign data_mem_w_li = dma_data_mem_w_lo | N1397;
  assign N1397 = sbuf_v_lo & sbuf_yumi_li;
  assign N1194 = ~dma_data_mem_w_lo;
  assign N1195 = N1398 & yumi_o;
  assign N1398 = decode[16] | decode[4];
  assign N1196 = dma_data_mem_v_lo | recover_lo;
  assign N1197 = N1195 | N1196;
  assign N1198 = ~N1197;
  assign N1199 = dma_data_mem_v_lo & N1192;
  assign N1200 = ~dma_data_mem_v_lo;
  assign N1201 = N1192 & N1200;
  assign N1202 = N1195 & N1201;
  assign track_mem_v_li = N1407 | N1408;
  assign N1407 = N1406 | miss_track_mem_v_lo;
  assign N1406 = N1401 | N1405;
  assign N1401 = yumi_o & N1400;
  assign N1400 = N1399 | partial_st;
  assign N1399 = decode[16] | decode[4];
  assign N1405 = N1402 & N1404;
  assign N1402 = v_tl_r & recover_lo;
  assign N1404 = N1403 | partial_st_tl;
  assign N1403 = decode_tl_r[16] | decode_tl_r[4];
  assign N1408 = tbuf_v_lo & tbuf_yumi_li;
  assign N1203 = tbuf_v_lo & tbuf_yumi_li;
  assign N1204 = N1410 & yumi_o;
  assign N1410 = N1409 | partial_st;
  assign N1409 = decode[16] | decode[4];
  assign N1205 = miss_track_mem_v_lo | recover_lo;
  assign N1206 = N1204 | N1205;
  assign N1207 = ~N1206;
  assign N1208 = miss_track_mem_v_lo & N1192;
  assign N1209 = ~miss_track_mem_v_lo;
  assign N1210 = N1192 & N1209;
  assign N1211 = N1204 & N1210;
  assign N1212 = ~miss_v;
  assign N1213 = miss_v;
  assign N1214 = N1414 & yumi_i;
  assign N1414 = N1413 & v_o;
  assign N1413 = N1412 | decode_v_r[4];
  assign N1412 = N1411 | decode_v_r[14];
  assign N1411 = decode_v_r[15] | decode_v_r[16];
  assign N1215 = N1418 & yumi_i;
  assign N1418 = N1417 & v_o;
  assign N1417 = N1416 | decode_v_r[4];
  assign N1416 = N1415 | decode_v_r[14];
  assign N1415 = decode_v_r[15] | decode_v_r[16];
  assign N1216 = decode_v_r[14];
  assign N1217 = ~N1216;
  assign N1218 = decode_v_r[15] | decode_v_r[4];
  assign N1219 = decode_v_r[15] | decode_v_r[4];
  assign N1220 = decode_v_r[15] | decode_v_r[4];
  assign N1221 = decode_v_r[15] | decode_v_r[4];
  assign N1222 = decode_v_r[15] | decode_v_r[4];
  assign N1223 = decode_v_r[15] | decode_v_r[4];
  assign N1224 = decode_v_r[15] | decode_v_r[4];
  assign N1225 = decode_v_r[15] | decode_v_r[4];
  assign N1226 = N1419 & tag_hit_v[7];
  assign N1419 = decode_v_r[15] | decode_v_r[4];
  assign N1227 = N1420 & tag_hit_v[6];
  assign N1420 = decode_v_r[15] | decode_v_r[4];
  assign N1228 = N1421 & tag_hit_v[5];
  assign N1421 = decode_v_r[15] | decode_v_r[4];
  assign N1229 = N1422 & tag_hit_v[4];
  assign N1422 = decode_v_r[15] | decode_v_r[4];
  assign N1230 = N1423 & tag_hit_v[3];
  assign N1423 = decode_v_r[15] | decode_v_r[4];
  assign N1231 = N1424 & tag_hit_v[2];
  assign N1424 = decode_v_r[15] | decode_v_r[4];
  assign N1232 = N1425 & tag_hit_v[1];
  assign N1425 = decode_v_r[15] | decode_v_r[4];
  assign N1233 = N1426 & tag_hit_v[0];
  assign N1426 = decode_v_r[15] | decode_v_r[4];
  assign sbuf_v_li = N1428 & yumi_i;
  assign N1428 = N1427 & v_o;
  assign N1427 = decode_v_r[15] | decode_v_r[4];
  assign N1264 = ~miss_v;
  assign N1265 = miss_v;
  assign sbuf_yumi_li = N1433 & N1440;
  assign N1433 = N1432 & N1377;
  assign N1432 = sbuf_v_lo & N1431;
  assign N1431 = ~N1430;
  assign N1430 = N1429 & yumi_o;
  assign N1429 = decode[16] | decode[4];
  assign N1440 = ~N1439;
  assign N1439 = N1437 & N1438;
  assign N1437 = N1435 & N1436;
  assign N1435 = v_tl_r & N1434;
  assign N1434 = decode_tl_r[16] | decode_tl_r[4];
  assign N1436 = ~v_we_o;
  assign N1438 = ~miss_v;
  assign sbuf_bypass_v_li = N1442 & v_we_o;
  assign N1442 = N1441 & v_tl_r;
  assign N1441 = decode_tl_r[16] | decode_tl_r[4];
  assign tbuf_v_li = N1445 & yumi_i;
  assign N1445 = N1444 & v_o;
  assign N1444 = decode_v_r[15] & N1443;
  assign N1443 = ~partial_st_v;
  assign N1266 = ~miss_v;
  assign N1267 = miss_v;
  assign tbuf_yumi_li = N1451 & N1458;
  assign N1451 = N1450 & N1375;
  assign N1450 = tbuf_v_lo & N1449;
  assign N1449 = ~N1448;
  assign N1448 = N1447 & yumi_o;
  assign N1447 = N1446 | partial_st;
  assign N1446 = decode[16] | decode[4];
  assign N1458 = ~N1457;
  assign N1457 = N1455 & N1456;
  assign N1455 = N1454 & N1436;
  assign N1454 = v_tl_r & N1453;
  assign N1453 = N1452 | partial_st_tl;
  assign N1452 = decode_tl_r[16] | decode_tl_r[4];
  assign N1456 = ~miss_v;
  assign tbuf_bypass_v_li = N1461 & v_we_o;
  assign N1461 = N1460 & v_tl_r;
  assign N1460 = N1459 | partial_st_tl;
  assign N1459 = decode_tl_r[16] | decode_tl_r[4];
  assign N2 = ~v_we_o;
  assign N1268 = ~decode_v_r[0];
  assign N1269 = ~decode_v_r[1];
  assign N1270 = N1268 & N1269;
  assign N1271 = N1268 & decode_v_r[1];
  assign N1272 = decode_v_r[0] & N1269;
  assign N1273 = decode_v_r[0] & decode_v_r[1];
  assign N1274 = ~decode_v_r[2];
  assign N1275 = N1270 & N1274;
  assign N1276 = N1270 & decode_v_r[2];
  assign N1277 = N1272 & N1274;
  assign N1278 = N1272 & decode_v_r[2];
  assign N1279 = N1271 & N1274;
  assign N1280 = N1271 & decode_v_r[2];
  assign N1281 = N1273 & N1274;
  assign N1282 = N1273 & decode_v_r[2];
  assign N1283 = ~decode_v_r[3];
  assign N1284 = N1275 & N1283;
  assign N1285 = N1275 & decode_v_r[3];
  assign N1286 = N1277 & N1283;
  assign N1287 = N1277 & decode_v_r[3];
  assign N1288 = N1279 & N1283;
  assign N1289 = N1279 & decode_v_r[3];
  assign N1290 = N1281 & N1283;
  assign N1291 = N1281 & decode_v_r[3];
  assign N1292 = N1276 & N1283;
  assign N1293 = N1276 & decode_v_r[3];
  assign N1294 = N1278 & N1283;
  assign N1295 = N1278 & decode_v_r[3];
  assign N1296 = N1280 & N1283;
  assign N1297 = N1280 & decode_v_r[3];
  assign N1298 = N1282 & N1283;
  assign N1299 = N1282 & decode_v_r[3];

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_tl_r_127_sv2v_reg <= 1'b0;
      data_tl_r_126_sv2v_reg <= 1'b0;
      data_tl_r_125_sv2v_reg <= 1'b0;
      data_tl_r_124_sv2v_reg <= 1'b0;
      data_tl_r_123_sv2v_reg <= 1'b0;
      data_tl_r_122_sv2v_reg <= 1'b0;
      data_tl_r_121_sv2v_reg <= 1'b0;
      data_tl_r_120_sv2v_reg <= 1'b0;
      data_tl_r_119_sv2v_reg <= 1'b0;
      data_tl_r_118_sv2v_reg <= 1'b0;
      data_tl_r_117_sv2v_reg <= 1'b0;
      data_tl_r_116_sv2v_reg <= 1'b0;
      data_tl_r_115_sv2v_reg <= 1'b0;
      data_tl_r_114_sv2v_reg <= 1'b0;
      data_tl_r_113_sv2v_reg <= 1'b0;
      data_tl_r_112_sv2v_reg <= 1'b0;
      data_tl_r_111_sv2v_reg <= 1'b0;
      data_tl_r_110_sv2v_reg <= 1'b0;
      data_tl_r_109_sv2v_reg <= 1'b0;
      data_tl_r_108_sv2v_reg <= 1'b0;
      data_tl_r_107_sv2v_reg <= 1'b0;
      data_tl_r_106_sv2v_reg <= 1'b0;
      data_tl_r_105_sv2v_reg <= 1'b0;
      data_tl_r_104_sv2v_reg <= 1'b0;
      data_tl_r_103_sv2v_reg <= 1'b0;
      data_tl_r_102_sv2v_reg <= 1'b0;
      data_tl_r_101_sv2v_reg <= 1'b0;
      data_tl_r_100_sv2v_reg <= 1'b0;
      data_tl_r_99_sv2v_reg <= 1'b0;
      data_tl_r_98_sv2v_reg <= 1'b0;
      data_tl_r_97_sv2v_reg <= 1'b0;
      data_tl_r_96_sv2v_reg <= 1'b0;
      data_tl_r_95_sv2v_reg <= 1'b0;
      data_tl_r_94_sv2v_reg <= 1'b0;
      data_tl_r_93_sv2v_reg <= 1'b0;
      data_tl_r_92_sv2v_reg <= 1'b0;
      data_tl_r_91_sv2v_reg <= 1'b0;
      data_tl_r_90_sv2v_reg <= 1'b0;
      data_tl_r_89_sv2v_reg <= 1'b0;
      data_tl_r_88_sv2v_reg <= 1'b0;
      data_tl_r_87_sv2v_reg <= 1'b0;
      data_tl_r_86_sv2v_reg <= 1'b0;
      data_tl_r_85_sv2v_reg <= 1'b0;
      data_tl_r_84_sv2v_reg <= 1'b0;
      data_tl_r_83_sv2v_reg <= 1'b0;
      data_tl_r_82_sv2v_reg <= 1'b0;
      data_tl_r_81_sv2v_reg <= 1'b0;
      data_tl_r_80_sv2v_reg <= 1'b0;
      data_tl_r_79_sv2v_reg <= 1'b0;
      data_tl_r_78_sv2v_reg <= 1'b0;
      data_tl_r_77_sv2v_reg <= 1'b0;
      data_tl_r_76_sv2v_reg <= 1'b0;
      data_tl_r_75_sv2v_reg <= 1'b0;
      data_tl_r_74_sv2v_reg <= 1'b0;
      data_tl_r_73_sv2v_reg <= 1'b0;
      data_tl_r_72_sv2v_reg <= 1'b0;
      data_tl_r_71_sv2v_reg <= 1'b0;
      data_tl_r_70_sv2v_reg <= 1'b0;
      data_tl_r_69_sv2v_reg <= 1'b0;
      data_tl_r_68_sv2v_reg <= 1'b0;
      data_tl_r_67_sv2v_reg <= 1'b0;
      data_tl_r_66_sv2v_reg <= 1'b0;
      data_tl_r_65_sv2v_reg <= 1'b0;
      data_tl_r_64_sv2v_reg <= 1'b0;
      data_tl_r_63_sv2v_reg <= 1'b0;
      data_tl_r_62_sv2v_reg <= 1'b0;
      data_tl_r_61_sv2v_reg <= 1'b0;
      data_tl_r_60_sv2v_reg <= 1'b0;
      data_tl_r_59_sv2v_reg <= 1'b0;
      data_tl_r_58_sv2v_reg <= 1'b0;
      data_tl_r_57_sv2v_reg <= 1'b0;
      data_tl_r_56_sv2v_reg <= 1'b0;
      data_tl_r_55_sv2v_reg <= 1'b0;
      data_tl_r_54_sv2v_reg <= 1'b0;
      data_tl_r_53_sv2v_reg <= 1'b0;
      data_tl_r_52_sv2v_reg <= 1'b0;
      data_tl_r_51_sv2v_reg <= 1'b0;
      data_tl_r_50_sv2v_reg <= 1'b0;
      decode_tl_r_20_sv2v_reg <= 1'b0;
      decode_tl_r_19_sv2v_reg <= 1'b0;
      decode_tl_r_18_sv2v_reg <= 1'b0;
      decode_tl_r_17_sv2v_reg <= 1'b0;
      decode_tl_r_16_sv2v_reg <= 1'b0;
      decode_tl_r_15_sv2v_reg <= 1'b0;
      decode_tl_r_14_sv2v_reg <= 1'b0;
      decode_tl_r_13_sv2v_reg <= 1'b0;
      decode_tl_r_12_sv2v_reg <= 1'b0;
      decode_tl_r_11_sv2v_reg <= 1'b0;
      decode_tl_r_10_sv2v_reg <= 1'b0;
      decode_tl_r_9_sv2v_reg <= 1'b0;
      decode_tl_r_8_sv2v_reg <= 1'b0;
      decode_tl_r_7_sv2v_reg <= 1'b0;
      decode_tl_r_6_sv2v_reg <= 1'b0;
      decode_tl_r_5_sv2v_reg <= 1'b0;
      decode_tl_r_4_sv2v_reg <= 1'b0;
      decode_tl_r_3_sv2v_reg <= 1'b0;
      decode_tl_r_2_sv2v_reg <= 1'b0;
      decode_tl_r_1_sv2v_reg <= 1'b0;
      decode_tl_r_0_sv2v_reg <= 1'b0;
      mask_tl_r_0_sv2v_reg <= 1'b0;
    end else if(N81) begin
      data_tl_r_127_sv2v_reg <= cache_pkt_i[143];
      data_tl_r_126_sv2v_reg <= cache_pkt_i[142];
      data_tl_r_125_sv2v_reg <= cache_pkt_i[141];
      data_tl_r_124_sv2v_reg <= cache_pkt_i[140];
      data_tl_r_123_sv2v_reg <= cache_pkt_i[139];
      data_tl_r_122_sv2v_reg <= cache_pkt_i[138];
      data_tl_r_121_sv2v_reg <= cache_pkt_i[137];
      data_tl_r_120_sv2v_reg <= cache_pkt_i[136];
      data_tl_r_119_sv2v_reg <= cache_pkt_i[135];
      data_tl_r_118_sv2v_reg <= cache_pkt_i[134];
      data_tl_r_117_sv2v_reg <= cache_pkt_i[133];
      data_tl_r_116_sv2v_reg <= cache_pkt_i[132];
      data_tl_r_115_sv2v_reg <= cache_pkt_i[131];
      data_tl_r_114_sv2v_reg <= cache_pkt_i[130];
      data_tl_r_113_sv2v_reg <= cache_pkt_i[129];
      data_tl_r_112_sv2v_reg <= cache_pkt_i[128];
      data_tl_r_111_sv2v_reg <= cache_pkt_i[127];
      data_tl_r_110_sv2v_reg <= cache_pkt_i[126];
      data_tl_r_109_sv2v_reg <= cache_pkt_i[125];
      data_tl_r_108_sv2v_reg <= cache_pkt_i[124];
      data_tl_r_107_sv2v_reg <= cache_pkt_i[123];
      data_tl_r_106_sv2v_reg <= cache_pkt_i[122];
      data_tl_r_105_sv2v_reg <= cache_pkt_i[121];
      data_tl_r_104_sv2v_reg <= cache_pkt_i[120];
      data_tl_r_103_sv2v_reg <= cache_pkt_i[119];
      data_tl_r_102_sv2v_reg <= cache_pkt_i[118];
      data_tl_r_101_sv2v_reg <= cache_pkt_i[117];
      data_tl_r_100_sv2v_reg <= cache_pkt_i[116];
      data_tl_r_99_sv2v_reg <= cache_pkt_i[115];
      data_tl_r_98_sv2v_reg <= cache_pkt_i[114];
      data_tl_r_97_sv2v_reg <= cache_pkt_i[113];
      data_tl_r_96_sv2v_reg <= cache_pkt_i[112];
      data_tl_r_95_sv2v_reg <= cache_pkt_i[111];
      data_tl_r_94_sv2v_reg <= cache_pkt_i[110];
      data_tl_r_93_sv2v_reg <= cache_pkt_i[109];
      data_tl_r_92_sv2v_reg <= cache_pkt_i[108];
      data_tl_r_91_sv2v_reg <= cache_pkt_i[107];
      data_tl_r_90_sv2v_reg <= cache_pkt_i[106];
      data_tl_r_89_sv2v_reg <= cache_pkt_i[105];
      data_tl_r_88_sv2v_reg <= cache_pkt_i[104];
      data_tl_r_87_sv2v_reg <= cache_pkt_i[103];
      data_tl_r_86_sv2v_reg <= cache_pkt_i[102];
      data_tl_r_85_sv2v_reg <= cache_pkt_i[101];
      data_tl_r_84_sv2v_reg <= cache_pkt_i[100];
      data_tl_r_83_sv2v_reg <= cache_pkt_i[99];
      data_tl_r_82_sv2v_reg <= cache_pkt_i[98];
      data_tl_r_81_sv2v_reg <= cache_pkt_i[97];
      data_tl_r_80_sv2v_reg <= cache_pkt_i[96];
      data_tl_r_79_sv2v_reg <= cache_pkt_i[95];
      data_tl_r_78_sv2v_reg <= cache_pkt_i[94];
      data_tl_r_77_sv2v_reg <= cache_pkt_i[93];
      data_tl_r_76_sv2v_reg <= cache_pkt_i[92];
      data_tl_r_75_sv2v_reg <= cache_pkt_i[91];
      data_tl_r_74_sv2v_reg <= cache_pkt_i[90];
      data_tl_r_73_sv2v_reg <= cache_pkt_i[89];
      data_tl_r_72_sv2v_reg <= cache_pkt_i[88];
      data_tl_r_71_sv2v_reg <= cache_pkt_i[87];
      data_tl_r_70_sv2v_reg <= cache_pkt_i[86];
      data_tl_r_69_sv2v_reg <= cache_pkt_i[85];
      data_tl_r_68_sv2v_reg <= cache_pkt_i[84];
      data_tl_r_67_sv2v_reg <= cache_pkt_i[83];
      data_tl_r_66_sv2v_reg <= cache_pkt_i[82];
      data_tl_r_65_sv2v_reg <= cache_pkt_i[81];
      data_tl_r_64_sv2v_reg <= cache_pkt_i[80];
      data_tl_r_63_sv2v_reg <= cache_pkt_i[79];
      data_tl_r_62_sv2v_reg <= cache_pkt_i[78];
      data_tl_r_61_sv2v_reg <= cache_pkt_i[77];
      data_tl_r_60_sv2v_reg <= cache_pkt_i[76];
      data_tl_r_59_sv2v_reg <= cache_pkt_i[75];
      data_tl_r_58_sv2v_reg <= cache_pkt_i[74];
      data_tl_r_57_sv2v_reg <= cache_pkt_i[73];
      data_tl_r_56_sv2v_reg <= cache_pkt_i[72];
      data_tl_r_55_sv2v_reg <= cache_pkt_i[71];
      data_tl_r_54_sv2v_reg <= cache_pkt_i[70];
      data_tl_r_53_sv2v_reg <= cache_pkt_i[69];
      data_tl_r_52_sv2v_reg <= cache_pkt_i[68];
      data_tl_r_51_sv2v_reg <= cache_pkt_i[67];
      data_tl_r_50_sv2v_reg <= cache_pkt_i[66];
      decode_tl_r_20_sv2v_reg <= decode[20];
      decode_tl_r_19_sv2v_reg <= decode[19];
      decode_tl_r_18_sv2v_reg <= decode[18];
      decode_tl_r_17_sv2v_reg <= decode[17];
      decode_tl_r_16_sv2v_reg <= decode[16];
      decode_tl_r_15_sv2v_reg <= decode[15];
      decode_tl_r_14_sv2v_reg <= decode[14];
      decode_tl_r_13_sv2v_reg <= decode[13];
      decode_tl_r_12_sv2v_reg <= decode[12];
      decode_tl_r_11_sv2v_reg <= decode[11];
      decode_tl_r_10_sv2v_reg <= decode[10];
      decode_tl_r_9_sv2v_reg <= decode[9];
      decode_tl_r_8_sv2v_reg <= decode[8];
      decode_tl_r_7_sv2v_reg <= decode[7];
      decode_tl_r_6_sv2v_reg <= decode[6];
      decode_tl_r_5_sv2v_reg <= decode[5];
      decode_tl_r_4_sv2v_reg <= decode[4];
      decode_tl_r_3_sv2v_reg <= decode[3];
      decode_tl_r_2_sv2v_reg <= decode[2];
      decode_tl_r_1_sv2v_reg <= decode[1];
      decode_tl_r_0_sv2v_reg <= decode[0];
      mask_tl_r_0_sv2v_reg <= cache_pkt_i[0];
    end 
    if(reset_i) begin
      data_tl_r_49_sv2v_reg <= 1'b0;
      data_tl_r_48_sv2v_reg <= 1'b0;
      data_tl_r_47_sv2v_reg <= 1'b0;
      data_tl_r_46_sv2v_reg <= 1'b0;
      data_tl_r_45_sv2v_reg <= 1'b0;
      data_tl_r_44_sv2v_reg <= 1'b0;
      data_tl_r_43_sv2v_reg <= 1'b0;
      data_tl_r_42_sv2v_reg <= 1'b0;
      data_tl_r_41_sv2v_reg <= 1'b0;
      data_tl_r_40_sv2v_reg <= 1'b0;
      data_tl_r_39_sv2v_reg <= 1'b0;
      data_tl_r_38_sv2v_reg <= 1'b0;
      data_tl_r_37_sv2v_reg <= 1'b0;
      data_tl_r_36_sv2v_reg <= 1'b0;
      data_tl_r_35_sv2v_reg <= 1'b0;
      data_tl_r_34_sv2v_reg <= 1'b0;
      data_tl_r_33_sv2v_reg <= 1'b0;
      data_tl_r_32_sv2v_reg <= 1'b0;
      data_tl_r_31_sv2v_reg <= 1'b0;
      data_tl_r_30_sv2v_reg <= 1'b0;
      data_tl_r_29_sv2v_reg <= 1'b0;
      data_tl_r_28_sv2v_reg <= 1'b0;
      data_tl_r_27_sv2v_reg <= 1'b0;
      data_tl_r_26_sv2v_reg <= 1'b0;
      data_tl_r_25_sv2v_reg <= 1'b0;
      data_tl_r_24_sv2v_reg <= 1'b0;
      data_tl_r_23_sv2v_reg <= 1'b0;
      data_tl_r_22_sv2v_reg <= 1'b0;
      data_tl_r_21_sv2v_reg <= 1'b0;
      data_tl_r_20_sv2v_reg <= 1'b0;
      data_tl_r_19_sv2v_reg <= 1'b0;
      data_tl_r_18_sv2v_reg <= 1'b0;
      data_tl_r_17_sv2v_reg <= 1'b0;
      data_tl_r_16_sv2v_reg <= 1'b0;
      data_tl_r_15_sv2v_reg <= 1'b0;
      data_tl_r_14_sv2v_reg <= 1'b0;
      data_tl_r_13_sv2v_reg <= 1'b0;
      data_tl_r_12_sv2v_reg <= 1'b0;
      data_tl_r_11_sv2v_reg <= 1'b0;
      data_tl_r_10_sv2v_reg <= 1'b0;
      data_tl_r_9_sv2v_reg <= 1'b0;
      data_tl_r_8_sv2v_reg <= 1'b0;
      data_tl_r_7_sv2v_reg <= 1'b0;
      data_tl_r_6_sv2v_reg <= 1'b0;
      data_tl_r_5_sv2v_reg <= 1'b0;
      data_tl_r_4_sv2v_reg <= 1'b0;
      data_tl_r_3_sv2v_reg <= 1'b0;
      data_tl_r_2_sv2v_reg <= 1'b0;
      data_tl_r_1_sv2v_reg <= 1'b0;
      data_tl_r_0_sv2v_reg <= 1'b0;
      mask_tl_r_15_sv2v_reg <= 1'b0;
      mask_tl_r_14_sv2v_reg <= 1'b0;
      mask_tl_r_13_sv2v_reg <= 1'b0;
      mask_tl_r_12_sv2v_reg <= 1'b0;
      mask_tl_r_11_sv2v_reg <= 1'b0;
      mask_tl_r_10_sv2v_reg <= 1'b0;
      mask_tl_r_9_sv2v_reg <= 1'b0;
      mask_tl_r_8_sv2v_reg <= 1'b0;
      mask_tl_r_7_sv2v_reg <= 1'b0;
      mask_tl_r_6_sv2v_reg <= 1'b0;
      mask_tl_r_5_sv2v_reg <= 1'b0;
      mask_tl_r_4_sv2v_reg <= 1'b0;
      mask_tl_r_3_sv2v_reg <= 1'b0;
      mask_tl_r_2_sv2v_reg <= 1'b0;
      mask_tl_r_1_sv2v_reg <= 1'b0;
      addr_tl_r_32_sv2v_reg <= 1'b0;
      addr_tl_r_31_sv2v_reg <= 1'b0;
      addr_tl_r_30_sv2v_reg <= 1'b0;
      addr_tl_r_29_sv2v_reg <= 1'b0;
      addr_tl_r_28_sv2v_reg <= 1'b0;
      addr_tl_r_27_sv2v_reg <= 1'b0;
      addr_tl_r_26_sv2v_reg <= 1'b0;
      addr_tl_r_25_sv2v_reg <= 1'b0;
      addr_tl_r_24_sv2v_reg <= 1'b0;
      addr_tl_r_23_sv2v_reg <= 1'b0;
      addr_tl_r_22_sv2v_reg <= 1'b0;
      addr_tl_r_21_sv2v_reg <= 1'b0;
      addr_tl_r_20_sv2v_reg <= 1'b0;
      addr_tl_r_19_sv2v_reg <= 1'b0;
      addr_tl_r_18_sv2v_reg <= 1'b0;
      addr_tl_r_17_sv2v_reg <= 1'b0;
      addr_tl_r_16_sv2v_reg <= 1'b0;
      addr_tl_r_15_sv2v_reg <= 1'b0;
      addr_tl_r_14_sv2v_reg <= 1'b0;
      addr_tl_r_13_sv2v_reg <= 1'b0;
      addr_tl_r_12_sv2v_reg <= 1'b0;
      addr_tl_r_11_sv2v_reg <= 1'b0;
      addr_tl_r_10_sv2v_reg <= 1'b0;
      addr_tl_r_9_sv2v_reg <= 1'b0;
      addr_tl_r_8_sv2v_reg <= 1'b0;
      addr_tl_r_7_sv2v_reg <= 1'b0;
      addr_tl_r_6_sv2v_reg <= 1'b0;
      addr_tl_r_5_sv2v_reg <= 1'b0;
      addr_tl_r_4_sv2v_reg <= 1'b0;
      addr_tl_r_3_sv2v_reg <= 1'b0;
      addr_tl_r_2_sv2v_reg <= 1'b0;
      addr_tl_r_1_sv2v_reg <= 1'b0;
      addr_tl_r_0_sv2v_reg <= 1'b0;
    end else if(N82) begin
      data_tl_r_49_sv2v_reg <= cache_pkt_i[65];
      data_tl_r_48_sv2v_reg <= cache_pkt_i[64];
      data_tl_r_47_sv2v_reg <= cache_pkt_i[63];
      data_tl_r_46_sv2v_reg <= cache_pkt_i[62];
      data_tl_r_45_sv2v_reg <= cache_pkt_i[61];
      data_tl_r_44_sv2v_reg <= cache_pkt_i[60];
      data_tl_r_43_sv2v_reg <= cache_pkt_i[59];
      data_tl_r_42_sv2v_reg <= cache_pkt_i[58];
      data_tl_r_41_sv2v_reg <= cache_pkt_i[57];
      data_tl_r_40_sv2v_reg <= cache_pkt_i[56];
      data_tl_r_39_sv2v_reg <= cache_pkt_i[55];
      data_tl_r_38_sv2v_reg <= cache_pkt_i[54];
      data_tl_r_37_sv2v_reg <= cache_pkt_i[53];
      data_tl_r_36_sv2v_reg <= cache_pkt_i[52];
      data_tl_r_35_sv2v_reg <= cache_pkt_i[51];
      data_tl_r_34_sv2v_reg <= cache_pkt_i[50];
      data_tl_r_33_sv2v_reg <= cache_pkt_i[49];
      data_tl_r_32_sv2v_reg <= cache_pkt_i[48];
      data_tl_r_31_sv2v_reg <= cache_pkt_i[47];
      data_tl_r_30_sv2v_reg <= cache_pkt_i[46];
      data_tl_r_29_sv2v_reg <= cache_pkt_i[45];
      data_tl_r_28_sv2v_reg <= cache_pkt_i[44];
      data_tl_r_27_sv2v_reg <= cache_pkt_i[43];
      data_tl_r_26_sv2v_reg <= cache_pkt_i[42];
      data_tl_r_25_sv2v_reg <= cache_pkt_i[41];
      data_tl_r_24_sv2v_reg <= cache_pkt_i[40];
      data_tl_r_23_sv2v_reg <= cache_pkt_i[39];
      data_tl_r_22_sv2v_reg <= cache_pkt_i[38];
      data_tl_r_21_sv2v_reg <= cache_pkt_i[37];
      data_tl_r_20_sv2v_reg <= cache_pkt_i[36];
      data_tl_r_19_sv2v_reg <= cache_pkt_i[35];
      data_tl_r_18_sv2v_reg <= cache_pkt_i[34];
      data_tl_r_17_sv2v_reg <= cache_pkt_i[33];
      data_tl_r_16_sv2v_reg <= cache_pkt_i[32];
      data_tl_r_15_sv2v_reg <= cache_pkt_i[31];
      data_tl_r_14_sv2v_reg <= cache_pkt_i[30];
      data_tl_r_13_sv2v_reg <= cache_pkt_i[29];
      data_tl_r_12_sv2v_reg <= cache_pkt_i[28];
      data_tl_r_11_sv2v_reg <= cache_pkt_i[27];
      data_tl_r_10_sv2v_reg <= cache_pkt_i[26];
      data_tl_r_9_sv2v_reg <= cache_pkt_i[25];
      data_tl_r_8_sv2v_reg <= cache_pkt_i[24];
      data_tl_r_7_sv2v_reg <= cache_pkt_i[23];
      data_tl_r_6_sv2v_reg <= cache_pkt_i[22];
      data_tl_r_5_sv2v_reg <= cache_pkt_i[21];
      data_tl_r_4_sv2v_reg <= cache_pkt_i[20];
      data_tl_r_3_sv2v_reg <= cache_pkt_i[19];
      data_tl_r_2_sv2v_reg <= cache_pkt_i[18];
      data_tl_r_1_sv2v_reg <= cache_pkt_i[17];
      data_tl_r_0_sv2v_reg <= cache_pkt_i[16];
      mask_tl_r_15_sv2v_reg <= cache_pkt_i[15];
      mask_tl_r_14_sv2v_reg <= cache_pkt_i[14];
      mask_tl_r_13_sv2v_reg <= cache_pkt_i[13];
      mask_tl_r_12_sv2v_reg <= cache_pkt_i[12];
      mask_tl_r_11_sv2v_reg <= cache_pkt_i[11];
      mask_tl_r_10_sv2v_reg <= cache_pkt_i[10];
      mask_tl_r_9_sv2v_reg <= cache_pkt_i[9];
      mask_tl_r_8_sv2v_reg <= cache_pkt_i[8];
      mask_tl_r_7_sv2v_reg <= cache_pkt_i[7];
      mask_tl_r_6_sv2v_reg <= cache_pkt_i[6];
      mask_tl_r_5_sv2v_reg <= cache_pkt_i[5];
      mask_tl_r_4_sv2v_reg <= cache_pkt_i[4];
      mask_tl_r_3_sv2v_reg <= cache_pkt_i[3];
      mask_tl_r_2_sv2v_reg <= cache_pkt_i[2];
      mask_tl_r_1_sv2v_reg <= cache_pkt_i[1];
      addr_tl_r_32_sv2v_reg <= cache_pkt_i[176];
      addr_tl_r_31_sv2v_reg <= cache_pkt_i[175];
      addr_tl_r_30_sv2v_reg <= cache_pkt_i[174];
      addr_tl_r_29_sv2v_reg <= cache_pkt_i[173];
      addr_tl_r_28_sv2v_reg <= cache_pkt_i[172];
      addr_tl_r_27_sv2v_reg <= cache_pkt_i[171];
      addr_tl_r_26_sv2v_reg <= cache_pkt_i[170];
      addr_tl_r_25_sv2v_reg <= cache_pkt_i[169];
      addr_tl_r_24_sv2v_reg <= cache_pkt_i[168];
      addr_tl_r_23_sv2v_reg <= cache_pkt_i[167];
      addr_tl_r_22_sv2v_reg <= cache_pkt_i[166];
      addr_tl_r_21_sv2v_reg <= cache_pkt_i[165];
      addr_tl_r_20_sv2v_reg <= cache_pkt_i[164];
      addr_tl_r_19_sv2v_reg <= cache_pkt_i[163];
      addr_tl_r_18_sv2v_reg <= cache_pkt_i[162];
      addr_tl_r_17_sv2v_reg <= cache_pkt_i[161];
      addr_tl_r_16_sv2v_reg <= cache_pkt_i[160];
      addr_tl_r_15_sv2v_reg <= cache_pkt_i[159];
      addr_tl_r_14_sv2v_reg <= cache_pkt_i[158];
      addr_tl_r_13_sv2v_reg <= cache_pkt_i[157];
      addr_tl_r_12_sv2v_reg <= cache_pkt_i[156];
      addr_tl_r_11_sv2v_reg <= cache_pkt_i[155];
      addr_tl_r_10_sv2v_reg <= cache_pkt_i[154];
      addr_tl_r_9_sv2v_reg <= cache_pkt_i[153];
      addr_tl_r_8_sv2v_reg <= cache_pkt_i[152];
      addr_tl_r_7_sv2v_reg <= cache_pkt_i[151];
      addr_tl_r_6_sv2v_reg <= cache_pkt_i[150];
      addr_tl_r_5_sv2v_reg <= cache_pkt_i[149];
      addr_tl_r_4_sv2v_reg <= cache_pkt_i[148];
      addr_tl_r_3_sv2v_reg <= cache_pkt_i[147];
      addr_tl_r_2_sv2v_reg <= cache_pkt_i[146];
      addr_tl_r_1_sv2v_reg <= cache_pkt_i[145];
      addr_tl_r_0_sv2v_reg <= cache_pkt_i[144];
    end 
    if(reset_i) begin
      v_tl_r_sv2v_reg <= 1'b0;
    end else if(N79) begin
      v_tl_r_sv2v_reg <= N80;
    end 
    if(N114) begin
      ld_data_v_r_1023_sv2v_reg <= data_mem_data_lo[1023];
      ld_data_v_r_1022_sv2v_reg <= data_mem_data_lo[1022];
      ld_data_v_r_1021_sv2v_reg <= data_mem_data_lo[1021];
      ld_data_v_r_1020_sv2v_reg <= data_mem_data_lo[1020];
      ld_data_v_r_1019_sv2v_reg <= data_mem_data_lo[1019];
      ld_data_v_r_1018_sv2v_reg <= data_mem_data_lo[1018];
      ld_data_v_r_1017_sv2v_reg <= data_mem_data_lo[1017];
      ld_data_v_r_1016_sv2v_reg <= data_mem_data_lo[1016];
      ld_data_v_r_1015_sv2v_reg <= data_mem_data_lo[1015];
      ld_data_v_r_1014_sv2v_reg <= data_mem_data_lo[1014];
      ld_data_v_r_1013_sv2v_reg <= data_mem_data_lo[1013];
      ld_data_v_r_1012_sv2v_reg <= data_mem_data_lo[1012];
      ld_data_v_r_1011_sv2v_reg <= data_mem_data_lo[1011];
      ld_data_v_r_1010_sv2v_reg <= data_mem_data_lo[1010];
      ld_data_v_r_1009_sv2v_reg <= data_mem_data_lo[1009];
      ld_data_v_r_1008_sv2v_reg <= data_mem_data_lo[1008];
      ld_data_v_r_1007_sv2v_reg <= data_mem_data_lo[1007];
      ld_data_v_r_1006_sv2v_reg <= data_mem_data_lo[1006];
      ld_data_v_r_1005_sv2v_reg <= data_mem_data_lo[1005];
      ld_data_v_r_1004_sv2v_reg <= data_mem_data_lo[1004];
      ld_data_v_r_1003_sv2v_reg <= data_mem_data_lo[1003];
      ld_data_v_r_1002_sv2v_reg <= data_mem_data_lo[1002];
      ld_data_v_r_1001_sv2v_reg <= data_mem_data_lo[1001];
      ld_data_v_r_1000_sv2v_reg <= data_mem_data_lo[1000];
      ld_data_v_r_999_sv2v_reg <= data_mem_data_lo[999];
      ld_data_v_r_998_sv2v_reg <= data_mem_data_lo[998];
      ld_data_v_r_997_sv2v_reg <= data_mem_data_lo[997];
      ld_data_v_r_996_sv2v_reg <= data_mem_data_lo[996];
      ld_data_v_r_995_sv2v_reg <= data_mem_data_lo[995];
      ld_data_v_r_994_sv2v_reg <= data_mem_data_lo[994];
      ld_data_v_r_993_sv2v_reg <= data_mem_data_lo[993];
      ld_data_v_r_992_sv2v_reg <= data_mem_data_lo[992];
      ld_data_v_r_991_sv2v_reg <= data_mem_data_lo[991];
      ld_data_v_r_990_sv2v_reg <= data_mem_data_lo[990];
      ld_data_v_r_989_sv2v_reg <= data_mem_data_lo[989];
      ld_data_v_r_988_sv2v_reg <= data_mem_data_lo[988];
      ld_data_v_r_987_sv2v_reg <= data_mem_data_lo[987];
      ld_data_v_r_986_sv2v_reg <= data_mem_data_lo[986];
      ld_data_v_r_985_sv2v_reg <= data_mem_data_lo[985];
      ld_data_v_r_984_sv2v_reg <= data_mem_data_lo[984];
      ld_data_v_r_983_sv2v_reg <= data_mem_data_lo[983];
      ld_data_v_r_982_sv2v_reg <= data_mem_data_lo[982];
      ld_data_v_r_981_sv2v_reg <= data_mem_data_lo[981];
      ld_data_v_r_980_sv2v_reg <= data_mem_data_lo[980];
      ld_data_v_r_979_sv2v_reg <= data_mem_data_lo[979];
      ld_data_v_r_978_sv2v_reg <= data_mem_data_lo[978];
      ld_data_v_r_977_sv2v_reg <= data_mem_data_lo[977];
      ld_data_v_r_976_sv2v_reg <= data_mem_data_lo[976];
      ld_data_v_r_975_sv2v_reg <= data_mem_data_lo[975];
      ld_data_v_r_974_sv2v_reg <= data_mem_data_lo[974];
      ld_data_v_r_973_sv2v_reg <= data_mem_data_lo[973];
      ld_data_v_r_972_sv2v_reg <= data_mem_data_lo[972];
      ld_data_v_r_971_sv2v_reg <= data_mem_data_lo[971];
      ld_data_v_r_970_sv2v_reg <= data_mem_data_lo[970];
      ld_data_v_r_969_sv2v_reg <= data_mem_data_lo[969];
      ld_data_v_r_968_sv2v_reg <= data_mem_data_lo[968];
      ld_data_v_r_967_sv2v_reg <= data_mem_data_lo[967];
      ld_data_v_r_966_sv2v_reg <= data_mem_data_lo[966];
      ld_data_v_r_965_sv2v_reg <= data_mem_data_lo[965];
      ld_data_v_r_964_sv2v_reg <= data_mem_data_lo[964];
      ld_data_v_r_963_sv2v_reg <= data_mem_data_lo[963];
      ld_data_v_r_962_sv2v_reg <= data_mem_data_lo[962];
      ld_data_v_r_961_sv2v_reg <= data_mem_data_lo[961];
      ld_data_v_r_960_sv2v_reg <= data_mem_data_lo[960];
      ld_data_v_r_959_sv2v_reg <= data_mem_data_lo[959];
      ld_data_v_r_958_sv2v_reg <= data_mem_data_lo[958];
      ld_data_v_r_957_sv2v_reg <= data_mem_data_lo[957];
    end 
    if(N113) begin
      ld_data_v_r_956_sv2v_reg <= data_mem_data_lo[956];
      ld_data_v_r_955_sv2v_reg <= data_mem_data_lo[955];
      ld_data_v_r_954_sv2v_reg <= data_mem_data_lo[954];
      ld_data_v_r_953_sv2v_reg <= data_mem_data_lo[953];
      ld_data_v_r_952_sv2v_reg <= data_mem_data_lo[952];
      ld_data_v_r_951_sv2v_reg <= data_mem_data_lo[951];
      ld_data_v_r_950_sv2v_reg <= data_mem_data_lo[950];
      ld_data_v_r_949_sv2v_reg <= data_mem_data_lo[949];
      ld_data_v_r_948_sv2v_reg <= data_mem_data_lo[948];
      ld_data_v_r_947_sv2v_reg <= data_mem_data_lo[947];
      ld_data_v_r_946_sv2v_reg <= data_mem_data_lo[946];
      ld_data_v_r_945_sv2v_reg <= data_mem_data_lo[945];
      ld_data_v_r_944_sv2v_reg <= data_mem_data_lo[944];
      ld_data_v_r_943_sv2v_reg <= data_mem_data_lo[943];
      ld_data_v_r_942_sv2v_reg <= data_mem_data_lo[942];
      ld_data_v_r_941_sv2v_reg <= data_mem_data_lo[941];
      ld_data_v_r_940_sv2v_reg <= data_mem_data_lo[940];
      ld_data_v_r_939_sv2v_reg <= data_mem_data_lo[939];
      ld_data_v_r_938_sv2v_reg <= data_mem_data_lo[938];
      ld_data_v_r_937_sv2v_reg <= data_mem_data_lo[937];
      ld_data_v_r_936_sv2v_reg <= data_mem_data_lo[936];
      ld_data_v_r_935_sv2v_reg <= data_mem_data_lo[935];
      ld_data_v_r_934_sv2v_reg <= data_mem_data_lo[934];
      ld_data_v_r_933_sv2v_reg <= data_mem_data_lo[933];
      ld_data_v_r_932_sv2v_reg <= data_mem_data_lo[932];
      ld_data_v_r_931_sv2v_reg <= data_mem_data_lo[931];
      ld_data_v_r_930_sv2v_reg <= data_mem_data_lo[930];
      ld_data_v_r_929_sv2v_reg <= data_mem_data_lo[929];
      ld_data_v_r_928_sv2v_reg <= data_mem_data_lo[928];
      ld_data_v_r_927_sv2v_reg <= data_mem_data_lo[927];
      ld_data_v_r_926_sv2v_reg <= data_mem_data_lo[926];
      ld_data_v_r_925_sv2v_reg <= data_mem_data_lo[925];
      ld_data_v_r_924_sv2v_reg <= data_mem_data_lo[924];
      ld_data_v_r_923_sv2v_reg <= data_mem_data_lo[923];
      ld_data_v_r_922_sv2v_reg <= data_mem_data_lo[922];
      ld_data_v_r_921_sv2v_reg <= data_mem_data_lo[921];
      ld_data_v_r_920_sv2v_reg <= data_mem_data_lo[920];
      ld_data_v_r_919_sv2v_reg <= data_mem_data_lo[919];
      ld_data_v_r_918_sv2v_reg <= data_mem_data_lo[918];
      ld_data_v_r_917_sv2v_reg <= data_mem_data_lo[917];
      ld_data_v_r_916_sv2v_reg <= data_mem_data_lo[916];
      ld_data_v_r_915_sv2v_reg <= data_mem_data_lo[915];
      ld_data_v_r_914_sv2v_reg <= data_mem_data_lo[914];
      ld_data_v_r_913_sv2v_reg <= data_mem_data_lo[913];
      ld_data_v_r_912_sv2v_reg <= data_mem_data_lo[912];
      ld_data_v_r_911_sv2v_reg <= data_mem_data_lo[911];
      ld_data_v_r_910_sv2v_reg <= data_mem_data_lo[910];
      ld_data_v_r_909_sv2v_reg <= data_mem_data_lo[909];
      ld_data_v_r_908_sv2v_reg <= data_mem_data_lo[908];
      ld_data_v_r_907_sv2v_reg <= data_mem_data_lo[907];
      ld_data_v_r_906_sv2v_reg <= data_mem_data_lo[906];
      ld_data_v_r_905_sv2v_reg <= data_mem_data_lo[905];
      ld_data_v_r_904_sv2v_reg <= data_mem_data_lo[904];
      ld_data_v_r_903_sv2v_reg <= data_mem_data_lo[903];
      ld_data_v_r_902_sv2v_reg <= data_mem_data_lo[902];
      ld_data_v_r_901_sv2v_reg <= data_mem_data_lo[901];
      ld_data_v_r_900_sv2v_reg <= data_mem_data_lo[900];
      ld_data_v_r_899_sv2v_reg <= data_mem_data_lo[899];
      ld_data_v_r_898_sv2v_reg <= data_mem_data_lo[898];
      ld_data_v_r_897_sv2v_reg <= data_mem_data_lo[897];
      ld_data_v_r_896_sv2v_reg <= data_mem_data_lo[896];
      ld_data_v_r_895_sv2v_reg <= data_mem_data_lo[895];
      ld_data_v_r_894_sv2v_reg <= data_mem_data_lo[894];
      ld_data_v_r_893_sv2v_reg <= data_mem_data_lo[893];
      ld_data_v_r_892_sv2v_reg <= data_mem_data_lo[892];
      ld_data_v_r_891_sv2v_reg <= data_mem_data_lo[891];
      ld_data_v_r_890_sv2v_reg <= data_mem_data_lo[890];
      ld_data_v_r_889_sv2v_reg <= data_mem_data_lo[889];
      ld_data_v_r_888_sv2v_reg <= data_mem_data_lo[888];
      ld_data_v_r_887_sv2v_reg <= data_mem_data_lo[887];
      ld_data_v_r_886_sv2v_reg <= data_mem_data_lo[886];
      ld_data_v_r_885_sv2v_reg <= data_mem_data_lo[885];
      ld_data_v_r_884_sv2v_reg <= data_mem_data_lo[884];
      ld_data_v_r_883_sv2v_reg <= data_mem_data_lo[883];
      ld_data_v_r_882_sv2v_reg <= data_mem_data_lo[882];
      ld_data_v_r_881_sv2v_reg <= data_mem_data_lo[881];
      ld_data_v_r_880_sv2v_reg <= data_mem_data_lo[880];
      ld_data_v_r_879_sv2v_reg <= data_mem_data_lo[879];
      ld_data_v_r_878_sv2v_reg <= data_mem_data_lo[878];
      ld_data_v_r_877_sv2v_reg <= data_mem_data_lo[877];
      ld_data_v_r_876_sv2v_reg <= data_mem_data_lo[876];
      ld_data_v_r_875_sv2v_reg <= data_mem_data_lo[875];
      ld_data_v_r_874_sv2v_reg <= data_mem_data_lo[874];
      ld_data_v_r_873_sv2v_reg <= data_mem_data_lo[873];
      ld_data_v_r_872_sv2v_reg <= data_mem_data_lo[872];
      ld_data_v_r_871_sv2v_reg <= data_mem_data_lo[871];
      ld_data_v_r_870_sv2v_reg <= data_mem_data_lo[870];
      ld_data_v_r_869_sv2v_reg <= data_mem_data_lo[869];
      ld_data_v_r_868_sv2v_reg <= data_mem_data_lo[868];
      ld_data_v_r_867_sv2v_reg <= data_mem_data_lo[867];
      ld_data_v_r_866_sv2v_reg <= data_mem_data_lo[866];
      ld_data_v_r_865_sv2v_reg <= data_mem_data_lo[865];
      ld_data_v_r_864_sv2v_reg <= data_mem_data_lo[864];
      ld_data_v_r_863_sv2v_reg <= data_mem_data_lo[863];
      ld_data_v_r_862_sv2v_reg <= data_mem_data_lo[862];
      ld_data_v_r_861_sv2v_reg <= data_mem_data_lo[861];
      ld_data_v_r_860_sv2v_reg <= data_mem_data_lo[860];
      ld_data_v_r_859_sv2v_reg <= data_mem_data_lo[859];
      ld_data_v_r_858_sv2v_reg <= data_mem_data_lo[858];
    end 
    if(N112) begin
      ld_data_v_r_857_sv2v_reg <= data_mem_data_lo[857];
      ld_data_v_r_856_sv2v_reg <= data_mem_data_lo[856];
      ld_data_v_r_855_sv2v_reg <= data_mem_data_lo[855];
      ld_data_v_r_854_sv2v_reg <= data_mem_data_lo[854];
      ld_data_v_r_853_sv2v_reg <= data_mem_data_lo[853];
      ld_data_v_r_852_sv2v_reg <= data_mem_data_lo[852];
      ld_data_v_r_851_sv2v_reg <= data_mem_data_lo[851];
      ld_data_v_r_850_sv2v_reg <= data_mem_data_lo[850];
      ld_data_v_r_849_sv2v_reg <= data_mem_data_lo[849];
      ld_data_v_r_848_sv2v_reg <= data_mem_data_lo[848];
      ld_data_v_r_847_sv2v_reg <= data_mem_data_lo[847];
      ld_data_v_r_846_sv2v_reg <= data_mem_data_lo[846];
      ld_data_v_r_845_sv2v_reg <= data_mem_data_lo[845];
      ld_data_v_r_844_sv2v_reg <= data_mem_data_lo[844];
      ld_data_v_r_843_sv2v_reg <= data_mem_data_lo[843];
      ld_data_v_r_842_sv2v_reg <= data_mem_data_lo[842];
      ld_data_v_r_841_sv2v_reg <= data_mem_data_lo[841];
      ld_data_v_r_840_sv2v_reg <= data_mem_data_lo[840];
      ld_data_v_r_839_sv2v_reg <= data_mem_data_lo[839];
      ld_data_v_r_838_sv2v_reg <= data_mem_data_lo[838];
      ld_data_v_r_837_sv2v_reg <= data_mem_data_lo[837];
      ld_data_v_r_836_sv2v_reg <= data_mem_data_lo[836];
      ld_data_v_r_835_sv2v_reg <= data_mem_data_lo[835];
      ld_data_v_r_834_sv2v_reg <= data_mem_data_lo[834];
      ld_data_v_r_833_sv2v_reg <= data_mem_data_lo[833];
      ld_data_v_r_832_sv2v_reg <= data_mem_data_lo[832];
      ld_data_v_r_831_sv2v_reg <= data_mem_data_lo[831];
      ld_data_v_r_830_sv2v_reg <= data_mem_data_lo[830];
      ld_data_v_r_829_sv2v_reg <= data_mem_data_lo[829];
      ld_data_v_r_828_sv2v_reg <= data_mem_data_lo[828];
      ld_data_v_r_827_sv2v_reg <= data_mem_data_lo[827];
      ld_data_v_r_826_sv2v_reg <= data_mem_data_lo[826];
      ld_data_v_r_825_sv2v_reg <= data_mem_data_lo[825];
      ld_data_v_r_824_sv2v_reg <= data_mem_data_lo[824];
      ld_data_v_r_823_sv2v_reg <= data_mem_data_lo[823];
      ld_data_v_r_822_sv2v_reg <= data_mem_data_lo[822];
      ld_data_v_r_821_sv2v_reg <= data_mem_data_lo[821];
      ld_data_v_r_820_sv2v_reg <= data_mem_data_lo[820];
      ld_data_v_r_819_sv2v_reg <= data_mem_data_lo[819];
      ld_data_v_r_818_sv2v_reg <= data_mem_data_lo[818];
      ld_data_v_r_817_sv2v_reg <= data_mem_data_lo[817];
      ld_data_v_r_816_sv2v_reg <= data_mem_data_lo[816];
      ld_data_v_r_815_sv2v_reg <= data_mem_data_lo[815];
      ld_data_v_r_814_sv2v_reg <= data_mem_data_lo[814];
      ld_data_v_r_813_sv2v_reg <= data_mem_data_lo[813];
      ld_data_v_r_812_sv2v_reg <= data_mem_data_lo[812];
      ld_data_v_r_811_sv2v_reg <= data_mem_data_lo[811];
      ld_data_v_r_810_sv2v_reg <= data_mem_data_lo[810];
      ld_data_v_r_809_sv2v_reg <= data_mem_data_lo[809];
      ld_data_v_r_808_sv2v_reg <= data_mem_data_lo[808];
      ld_data_v_r_807_sv2v_reg <= data_mem_data_lo[807];
      ld_data_v_r_806_sv2v_reg <= data_mem_data_lo[806];
      ld_data_v_r_805_sv2v_reg <= data_mem_data_lo[805];
      ld_data_v_r_804_sv2v_reg <= data_mem_data_lo[804];
      ld_data_v_r_803_sv2v_reg <= data_mem_data_lo[803];
      ld_data_v_r_802_sv2v_reg <= data_mem_data_lo[802];
      ld_data_v_r_801_sv2v_reg <= data_mem_data_lo[801];
      ld_data_v_r_800_sv2v_reg <= data_mem_data_lo[800];
      ld_data_v_r_799_sv2v_reg <= data_mem_data_lo[799];
      ld_data_v_r_798_sv2v_reg <= data_mem_data_lo[798];
      ld_data_v_r_797_sv2v_reg <= data_mem_data_lo[797];
      ld_data_v_r_796_sv2v_reg <= data_mem_data_lo[796];
      ld_data_v_r_795_sv2v_reg <= data_mem_data_lo[795];
      ld_data_v_r_794_sv2v_reg <= data_mem_data_lo[794];
      ld_data_v_r_793_sv2v_reg <= data_mem_data_lo[793];
      ld_data_v_r_792_sv2v_reg <= data_mem_data_lo[792];
      ld_data_v_r_791_sv2v_reg <= data_mem_data_lo[791];
      ld_data_v_r_790_sv2v_reg <= data_mem_data_lo[790];
      ld_data_v_r_789_sv2v_reg <= data_mem_data_lo[789];
      ld_data_v_r_788_sv2v_reg <= data_mem_data_lo[788];
      ld_data_v_r_787_sv2v_reg <= data_mem_data_lo[787];
      ld_data_v_r_786_sv2v_reg <= data_mem_data_lo[786];
      ld_data_v_r_785_sv2v_reg <= data_mem_data_lo[785];
      ld_data_v_r_784_sv2v_reg <= data_mem_data_lo[784];
      ld_data_v_r_783_sv2v_reg <= data_mem_data_lo[783];
      ld_data_v_r_782_sv2v_reg <= data_mem_data_lo[782];
      ld_data_v_r_781_sv2v_reg <= data_mem_data_lo[781];
      ld_data_v_r_780_sv2v_reg <= data_mem_data_lo[780];
      ld_data_v_r_779_sv2v_reg <= data_mem_data_lo[779];
      ld_data_v_r_778_sv2v_reg <= data_mem_data_lo[778];
      ld_data_v_r_777_sv2v_reg <= data_mem_data_lo[777];
      ld_data_v_r_776_sv2v_reg <= data_mem_data_lo[776];
      ld_data_v_r_775_sv2v_reg <= data_mem_data_lo[775];
      ld_data_v_r_774_sv2v_reg <= data_mem_data_lo[774];
      ld_data_v_r_773_sv2v_reg <= data_mem_data_lo[773];
      ld_data_v_r_772_sv2v_reg <= data_mem_data_lo[772];
      ld_data_v_r_771_sv2v_reg <= data_mem_data_lo[771];
      ld_data_v_r_770_sv2v_reg <= data_mem_data_lo[770];
      ld_data_v_r_769_sv2v_reg <= data_mem_data_lo[769];
      ld_data_v_r_768_sv2v_reg <= data_mem_data_lo[768];
      ld_data_v_r_767_sv2v_reg <= data_mem_data_lo[767];
      ld_data_v_r_766_sv2v_reg <= data_mem_data_lo[766];
      ld_data_v_r_765_sv2v_reg <= data_mem_data_lo[765];
      ld_data_v_r_764_sv2v_reg <= data_mem_data_lo[764];
      ld_data_v_r_763_sv2v_reg <= data_mem_data_lo[763];
      ld_data_v_r_762_sv2v_reg <= data_mem_data_lo[762];
      ld_data_v_r_761_sv2v_reg <= data_mem_data_lo[761];
      ld_data_v_r_760_sv2v_reg <= data_mem_data_lo[760];
      ld_data_v_r_759_sv2v_reg <= data_mem_data_lo[759];
    end 
    if(N111) begin
      ld_data_v_r_758_sv2v_reg <= data_mem_data_lo[758];
      ld_data_v_r_757_sv2v_reg <= data_mem_data_lo[757];
      ld_data_v_r_756_sv2v_reg <= data_mem_data_lo[756];
      ld_data_v_r_755_sv2v_reg <= data_mem_data_lo[755];
      ld_data_v_r_754_sv2v_reg <= data_mem_data_lo[754];
      ld_data_v_r_753_sv2v_reg <= data_mem_data_lo[753];
      ld_data_v_r_752_sv2v_reg <= data_mem_data_lo[752];
      ld_data_v_r_751_sv2v_reg <= data_mem_data_lo[751];
      ld_data_v_r_750_sv2v_reg <= data_mem_data_lo[750];
      ld_data_v_r_749_sv2v_reg <= data_mem_data_lo[749];
      ld_data_v_r_748_sv2v_reg <= data_mem_data_lo[748];
      ld_data_v_r_747_sv2v_reg <= data_mem_data_lo[747];
      ld_data_v_r_746_sv2v_reg <= data_mem_data_lo[746];
      ld_data_v_r_745_sv2v_reg <= data_mem_data_lo[745];
      ld_data_v_r_744_sv2v_reg <= data_mem_data_lo[744];
      ld_data_v_r_743_sv2v_reg <= data_mem_data_lo[743];
      ld_data_v_r_742_sv2v_reg <= data_mem_data_lo[742];
      ld_data_v_r_741_sv2v_reg <= data_mem_data_lo[741];
      ld_data_v_r_740_sv2v_reg <= data_mem_data_lo[740];
      ld_data_v_r_739_sv2v_reg <= data_mem_data_lo[739];
      ld_data_v_r_738_sv2v_reg <= data_mem_data_lo[738];
      ld_data_v_r_737_sv2v_reg <= data_mem_data_lo[737];
      ld_data_v_r_736_sv2v_reg <= data_mem_data_lo[736];
      ld_data_v_r_735_sv2v_reg <= data_mem_data_lo[735];
      ld_data_v_r_734_sv2v_reg <= data_mem_data_lo[734];
      ld_data_v_r_733_sv2v_reg <= data_mem_data_lo[733];
      ld_data_v_r_732_sv2v_reg <= data_mem_data_lo[732];
      ld_data_v_r_731_sv2v_reg <= data_mem_data_lo[731];
      ld_data_v_r_730_sv2v_reg <= data_mem_data_lo[730];
      ld_data_v_r_729_sv2v_reg <= data_mem_data_lo[729];
      ld_data_v_r_728_sv2v_reg <= data_mem_data_lo[728];
      ld_data_v_r_727_sv2v_reg <= data_mem_data_lo[727];
      ld_data_v_r_726_sv2v_reg <= data_mem_data_lo[726];
      ld_data_v_r_725_sv2v_reg <= data_mem_data_lo[725];
      ld_data_v_r_724_sv2v_reg <= data_mem_data_lo[724];
      ld_data_v_r_723_sv2v_reg <= data_mem_data_lo[723];
      ld_data_v_r_722_sv2v_reg <= data_mem_data_lo[722];
      ld_data_v_r_721_sv2v_reg <= data_mem_data_lo[721];
      ld_data_v_r_720_sv2v_reg <= data_mem_data_lo[720];
      ld_data_v_r_719_sv2v_reg <= data_mem_data_lo[719];
      ld_data_v_r_718_sv2v_reg <= data_mem_data_lo[718];
      ld_data_v_r_717_sv2v_reg <= data_mem_data_lo[717];
      ld_data_v_r_716_sv2v_reg <= data_mem_data_lo[716];
      ld_data_v_r_715_sv2v_reg <= data_mem_data_lo[715];
      ld_data_v_r_714_sv2v_reg <= data_mem_data_lo[714];
      ld_data_v_r_713_sv2v_reg <= data_mem_data_lo[713];
      ld_data_v_r_712_sv2v_reg <= data_mem_data_lo[712];
      ld_data_v_r_711_sv2v_reg <= data_mem_data_lo[711];
      ld_data_v_r_710_sv2v_reg <= data_mem_data_lo[710];
      ld_data_v_r_709_sv2v_reg <= data_mem_data_lo[709];
      ld_data_v_r_708_sv2v_reg <= data_mem_data_lo[708];
      ld_data_v_r_707_sv2v_reg <= data_mem_data_lo[707];
      ld_data_v_r_706_sv2v_reg <= data_mem_data_lo[706];
      ld_data_v_r_705_sv2v_reg <= data_mem_data_lo[705];
      ld_data_v_r_704_sv2v_reg <= data_mem_data_lo[704];
      ld_data_v_r_703_sv2v_reg <= data_mem_data_lo[703];
      ld_data_v_r_702_sv2v_reg <= data_mem_data_lo[702];
      ld_data_v_r_701_sv2v_reg <= data_mem_data_lo[701];
      ld_data_v_r_700_sv2v_reg <= data_mem_data_lo[700];
      ld_data_v_r_699_sv2v_reg <= data_mem_data_lo[699];
      ld_data_v_r_698_sv2v_reg <= data_mem_data_lo[698];
      ld_data_v_r_697_sv2v_reg <= data_mem_data_lo[697];
      ld_data_v_r_696_sv2v_reg <= data_mem_data_lo[696];
      ld_data_v_r_695_sv2v_reg <= data_mem_data_lo[695];
      ld_data_v_r_694_sv2v_reg <= data_mem_data_lo[694];
      ld_data_v_r_693_sv2v_reg <= data_mem_data_lo[693];
      ld_data_v_r_692_sv2v_reg <= data_mem_data_lo[692];
      ld_data_v_r_691_sv2v_reg <= data_mem_data_lo[691];
      ld_data_v_r_690_sv2v_reg <= data_mem_data_lo[690];
      ld_data_v_r_689_sv2v_reg <= data_mem_data_lo[689];
      ld_data_v_r_688_sv2v_reg <= data_mem_data_lo[688];
      ld_data_v_r_687_sv2v_reg <= data_mem_data_lo[687];
      ld_data_v_r_686_sv2v_reg <= data_mem_data_lo[686];
      ld_data_v_r_685_sv2v_reg <= data_mem_data_lo[685];
      ld_data_v_r_684_sv2v_reg <= data_mem_data_lo[684];
      ld_data_v_r_683_sv2v_reg <= data_mem_data_lo[683];
      ld_data_v_r_682_sv2v_reg <= data_mem_data_lo[682];
      ld_data_v_r_681_sv2v_reg <= data_mem_data_lo[681];
      ld_data_v_r_680_sv2v_reg <= data_mem_data_lo[680];
      ld_data_v_r_679_sv2v_reg <= data_mem_data_lo[679];
      ld_data_v_r_678_sv2v_reg <= data_mem_data_lo[678];
      ld_data_v_r_677_sv2v_reg <= data_mem_data_lo[677];
      ld_data_v_r_676_sv2v_reg <= data_mem_data_lo[676];
      ld_data_v_r_675_sv2v_reg <= data_mem_data_lo[675];
      ld_data_v_r_674_sv2v_reg <= data_mem_data_lo[674];
      ld_data_v_r_673_sv2v_reg <= data_mem_data_lo[673];
      ld_data_v_r_672_sv2v_reg <= data_mem_data_lo[672];
      ld_data_v_r_671_sv2v_reg <= data_mem_data_lo[671];
      ld_data_v_r_670_sv2v_reg <= data_mem_data_lo[670];
      ld_data_v_r_669_sv2v_reg <= data_mem_data_lo[669];
      ld_data_v_r_668_sv2v_reg <= data_mem_data_lo[668];
      ld_data_v_r_667_sv2v_reg <= data_mem_data_lo[667];
      ld_data_v_r_666_sv2v_reg <= data_mem_data_lo[666];
      ld_data_v_r_665_sv2v_reg <= data_mem_data_lo[665];
      ld_data_v_r_664_sv2v_reg <= data_mem_data_lo[664];
      ld_data_v_r_663_sv2v_reg <= data_mem_data_lo[663];
      ld_data_v_r_662_sv2v_reg <= data_mem_data_lo[662];
      ld_data_v_r_661_sv2v_reg <= data_mem_data_lo[661];
      ld_data_v_r_660_sv2v_reg <= data_mem_data_lo[660];
    end 
    if(N110) begin
      ld_data_v_r_659_sv2v_reg <= data_mem_data_lo[659];
      ld_data_v_r_658_sv2v_reg <= data_mem_data_lo[658];
      ld_data_v_r_657_sv2v_reg <= data_mem_data_lo[657];
      ld_data_v_r_656_sv2v_reg <= data_mem_data_lo[656];
      ld_data_v_r_655_sv2v_reg <= data_mem_data_lo[655];
      ld_data_v_r_654_sv2v_reg <= data_mem_data_lo[654];
      ld_data_v_r_653_sv2v_reg <= data_mem_data_lo[653];
      ld_data_v_r_652_sv2v_reg <= data_mem_data_lo[652];
      ld_data_v_r_651_sv2v_reg <= data_mem_data_lo[651];
      ld_data_v_r_650_sv2v_reg <= data_mem_data_lo[650];
      ld_data_v_r_649_sv2v_reg <= data_mem_data_lo[649];
      ld_data_v_r_648_sv2v_reg <= data_mem_data_lo[648];
      ld_data_v_r_647_sv2v_reg <= data_mem_data_lo[647];
      ld_data_v_r_646_sv2v_reg <= data_mem_data_lo[646];
      ld_data_v_r_645_sv2v_reg <= data_mem_data_lo[645];
      ld_data_v_r_644_sv2v_reg <= data_mem_data_lo[644];
      ld_data_v_r_643_sv2v_reg <= data_mem_data_lo[643];
      ld_data_v_r_642_sv2v_reg <= data_mem_data_lo[642];
      ld_data_v_r_641_sv2v_reg <= data_mem_data_lo[641];
      ld_data_v_r_640_sv2v_reg <= data_mem_data_lo[640];
      ld_data_v_r_639_sv2v_reg <= data_mem_data_lo[639];
      ld_data_v_r_638_sv2v_reg <= data_mem_data_lo[638];
      ld_data_v_r_637_sv2v_reg <= data_mem_data_lo[637];
      ld_data_v_r_636_sv2v_reg <= data_mem_data_lo[636];
      ld_data_v_r_635_sv2v_reg <= data_mem_data_lo[635];
      ld_data_v_r_634_sv2v_reg <= data_mem_data_lo[634];
      ld_data_v_r_633_sv2v_reg <= data_mem_data_lo[633];
      ld_data_v_r_632_sv2v_reg <= data_mem_data_lo[632];
      ld_data_v_r_631_sv2v_reg <= data_mem_data_lo[631];
      ld_data_v_r_630_sv2v_reg <= data_mem_data_lo[630];
      ld_data_v_r_629_sv2v_reg <= data_mem_data_lo[629];
      ld_data_v_r_628_sv2v_reg <= data_mem_data_lo[628];
      ld_data_v_r_627_sv2v_reg <= data_mem_data_lo[627];
      ld_data_v_r_626_sv2v_reg <= data_mem_data_lo[626];
      ld_data_v_r_625_sv2v_reg <= data_mem_data_lo[625];
      ld_data_v_r_624_sv2v_reg <= data_mem_data_lo[624];
      ld_data_v_r_623_sv2v_reg <= data_mem_data_lo[623];
      ld_data_v_r_622_sv2v_reg <= data_mem_data_lo[622];
      ld_data_v_r_621_sv2v_reg <= data_mem_data_lo[621];
      ld_data_v_r_620_sv2v_reg <= data_mem_data_lo[620];
      ld_data_v_r_619_sv2v_reg <= data_mem_data_lo[619];
      ld_data_v_r_618_sv2v_reg <= data_mem_data_lo[618];
      ld_data_v_r_617_sv2v_reg <= data_mem_data_lo[617];
      ld_data_v_r_616_sv2v_reg <= data_mem_data_lo[616];
      ld_data_v_r_615_sv2v_reg <= data_mem_data_lo[615];
      ld_data_v_r_614_sv2v_reg <= data_mem_data_lo[614];
      ld_data_v_r_613_sv2v_reg <= data_mem_data_lo[613];
      ld_data_v_r_612_sv2v_reg <= data_mem_data_lo[612];
      ld_data_v_r_611_sv2v_reg <= data_mem_data_lo[611];
      ld_data_v_r_610_sv2v_reg <= data_mem_data_lo[610];
      ld_data_v_r_609_sv2v_reg <= data_mem_data_lo[609];
      ld_data_v_r_608_sv2v_reg <= data_mem_data_lo[608];
      ld_data_v_r_607_sv2v_reg <= data_mem_data_lo[607];
      ld_data_v_r_606_sv2v_reg <= data_mem_data_lo[606];
      ld_data_v_r_605_sv2v_reg <= data_mem_data_lo[605];
      ld_data_v_r_604_sv2v_reg <= data_mem_data_lo[604];
      ld_data_v_r_603_sv2v_reg <= data_mem_data_lo[603];
      ld_data_v_r_602_sv2v_reg <= data_mem_data_lo[602];
      ld_data_v_r_601_sv2v_reg <= data_mem_data_lo[601];
      ld_data_v_r_600_sv2v_reg <= data_mem_data_lo[600];
      ld_data_v_r_599_sv2v_reg <= data_mem_data_lo[599];
      ld_data_v_r_598_sv2v_reg <= data_mem_data_lo[598];
      ld_data_v_r_597_sv2v_reg <= data_mem_data_lo[597];
      ld_data_v_r_596_sv2v_reg <= data_mem_data_lo[596];
      ld_data_v_r_595_sv2v_reg <= data_mem_data_lo[595];
      ld_data_v_r_594_sv2v_reg <= data_mem_data_lo[594];
      ld_data_v_r_593_sv2v_reg <= data_mem_data_lo[593];
      ld_data_v_r_592_sv2v_reg <= data_mem_data_lo[592];
      ld_data_v_r_591_sv2v_reg <= data_mem_data_lo[591];
      ld_data_v_r_590_sv2v_reg <= data_mem_data_lo[590];
      ld_data_v_r_589_sv2v_reg <= data_mem_data_lo[589];
      ld_data_v_r_588_sv2v_reg <= data_mem_data_lo[588];
      ld_data_v_r_587_sv2v_reg <= data_mem_data_lo[587];
      ld_data_v_r_586_sv2v_reg <= data_mem_data_lo[586];
      ld_data_v_r_585_sv2v_reg <= data_mem_data_lo[585];
      ld_data_v_r_584_sv2v_reg <= data_mem_data_lo[584];
      ld_data_v_r_583_sv2v_reg <= data_mem_data_lo[583];
      ld_data_v_r_582_sv2v_reg <= data_mem_data_lo[582];
      ld_data_v_r_581_sv2v_reg <= data_mem_data_lo[581];
      ld_data_v_r_580_sv2v_reg <= data_mem_data_lo[580];
      ld_data_v_r_579_sv2v_reg <= data_mem_data_lo[579];
      ld_data_v_r_578_sv2v_reg <= data_mem_data_lo[578];
      ld_data_v_r_577_sv2v_reg <= data_mem_data_lo[577];
      ld_data_v_r_576_sv2v_reg <= data_mem_data_lo[576];
      ld_data_v_r_575_sv2v_reg <= data_mem_data_lo[575];
      ld_data_v_r_574_sv2v_reg <= data_mem_data_lo[574];
      ld_data_v_r_573_sv2v_reg <= data_mem_data_lo[573];
      ld_data_v_r_572_sv2v_reg <= data_mem_data_lo[572];
      ld_data_v_r_571_sv2v_reg <= data_mem_data_lo[571];
      ld_data_v_r_570_sv2v_reg <= data_mem_data_lo[570];
      ld_data_v_r_569_sv2v_reg <= data_mem_data_lo[569];
      ld_data_v_r_568_sv2v_reg <= data_mem_data_lo[568];
      ld_data_v_r_567_sv2v_reg <= data_mem_data_lo[567];
      ld_data_v_r_566_sv2v_reg <= data_mem_data_lo[566];
      ld_data_v_r_565_sv2v_reg <= data_mem_data_lo[565];
      ld_data_v_r_564_sv2v_reg <= data_mem_data_lo[564];
      ld_data_v_r_563_sv2v_reg <= data_mem_data_lo[563];
      ld_data_v_r_562_sv2v_reg <= data_mem_data_lo[562];
      ld_data_v_r_561_sv2v_reg <= data_mem_data_lo[561];
    end 
    if(N109) begin
      ld_data_v_r_560_sv2v_reg <= data_mem_data_lo[560];
      ld_data_v_r_559_sv2v_reg <= data_mem_data_lo[559];
      ld_data_v_r_558_sv2v_reg <= data_mem_data_lo[558];
      ld_data_v_r_557_sv2v_reg <= data_mem_data_lo[557];
      ld_data_v_r_556_sv2v_reg <= data_mem_data_lo[556];
      ld_data_v_r_555_sv2v_reg <= data_mem_data_lo[555];
      ld_data_v_r_554_sv2v_reg <= data_mem_data_lo[554];
      ld_data_v_r_553_sv2v_reg <= data_mem_data_lo[553];
      ld_data_v_r_552_sv2v_reg <= data_mem_data_lo[552];
      ld_data_v_r_551_sv2v_reg <= data_mem_data_lo[551];
      ld_data_v_r_550_sv2v_reg <= data_mem_data_lo[550];
      ld_data_v_r_549_sv2v_reg <= data_mem_data_lo[549];
      ld_data_v_r_548_sv2v_reg <= data_mem_data_lo[548];
      ld_data_v_r_547_sv2v_reg <= data_mem_data_lo[547];
      ld_data_v_r_546_sv2v_reg <= data_mem_data_lo[546];
      ld_data_v_r_545_sv2v_reg <= data_mem_data_lo[545];
      ld_data_v_r_544_sv2v_reg <= data_mem_data_lo[544];
      ld_data_v_r_543_sv2v_reg <= data_mem_data_lo[543];
      ld_data_v_r_542_sv2v_reg <= data_mem_data_lo[542];
      ld_data_v_r_541_sv2v_reg <= data_mem_data_lo[541];
      ld_data_v_r_540_sv2v_reg <= data_mem_data_lo[540];
      ld_data_v_r_539_sv2v_reg <= data_mem_data_lo[539];
      ld_data_v_r_538_sv2v_reg <= data_mem_data_lo[538];
      ld_data_v_r_537_sv2v_reg <= data_mem_data_lo[537];
      ld_data_v_r_536_sv2v_reg <= data_mem_data_lo[536];
      ld_data_v_r_535_sv2v_reg <= data_mem_data_lo[535];
      ld_data_v_r_534_sv2v_reg <= data_mem_data_lo[534];
      ld_data_v_r_533_sv2v_reg <= data_mem_data_lo[533];
      ld_data_v_r_532_sv2v_reg <= data_mem_data_lo[532];
      ld_data_v_r_531_sv2v_reg <= data_mem_data_lo[531];
      ld_data_v_r_530_sv2v_reg <= data_mem_data_lo[530];
      ld_data_v_r_529_sv2v_reg <= data_mem_data_lo[529];
      ld_data_v_r_528_sv2v_reg <= data_mem_data_lo[528];
      ld_data_v_r_527_sv2v_reg <= data_mem_data_lo[527];
      ld_data_v_r_526_sv2v_reg <= data_mem_data_lo[526];
      ld_data_v_r_525_sv2v_reg <= data_mem_data_lo[525];
      ld_data_v_r_524_sv2v_reg <= data_mem_data_lo[524];
      ld_data_v_r_523_sv2v_reg <= data_mem_data_lo[523];
      ld_data_v_r_522_sv2v_reg <= data_mem_data_lo[522];
      ld_data_v_r_521_sv2v_reg <= data_mem_data_lo[521];
      ld_data_v_r_520_sv2v_reg <= data_mem_data_lo[520];
      ld_data_v_r_519_sv2v_reg <= data_mem_data_lo[519];
      ld_data_v_r_518_sv2v_reg <= data_mem_data_lo[518];
      ld_data_v_r_517_sv2v_reg <= data_mem_data_lo[517];
      ld_data_v_r_516_sv2v_reg <= data_mem_data_lo[516];
      ld_data_v_r_515_sv2v_reg <= data_mem_data_lo[515];
      ld_data_v_r_514_sv2v_reg <= data_mem_data_lo[514];
      ld_data_v_r_513_sv2v_reg <= data_mem_data_lo[513];
      ld_data_v_r_512_sv2v_reg <= data_mem_data_lo[512];
      ld_data_v_r_511_sv2v_reg <= data_mem_data_lo[511];
      ld_data_v_r_510_sv2v_reg <= data_mem_data_lo[510];
      ld_data_v_r_509_sv2v_reg <= data_mem_data_lo[509];
      ld_data_v_r_508_sv2v_reg <= data_mem_data_lo[508];
      ld_data_v_r_507_sv2v_reg <= data_mem_data_lo[507];
      ld_data_v_r_506_sv2v_reg <= data_mem_data_lo[506];
      ld_data_v_r_505_sv2v_reg <= data_mem_data_lo[505];
      ld_data_v_r_504_sv2v_reg <= data_mem_data_lo[504];
      ld_data_v_r_503_sv2v_reg <= data_mem_data_lo[503];
      ld_data_v_r_502_sv2v_reg <= data_mem_data_lo[502];
      ld_data_v_r_501_sv2v_reg <= data_mem_data_lo[501];
      ld_data_v_r_500_sv2v_reg <= data_mem_data_lo[500];
      ld_data_v_r_499_sv2v_reg <= data_mem_data_lo[499];
      ld_data_v_r_498_sv2v_reg <= data_mem_data_lo[498];
      ld_data_v_r_497_sv2v_reg <= data_mem_data_lo[497];
      ld_data_v_r_496_sv2v_reg <= data_mem_data_lo[496];
      ld_data_v_r_495_sv2v_reg <= data_mem_data_lo[495];
      ld_data_v_r_494_sv2v_reg <= data_mem_data_lo[494];
      ld_data_v_r_493_sv2v_reg <= data_mem_data_lo[493];
      ld_data_v_r_492_sv2v_reg <= data_mem_data_lo[492];
      ld_data_v_r_491_sv2v_reg <= data_mem_data_lo[491];
      ld_data_v_r_490_sv2v_reg <= data_mem_data_lo[490];
      ld_data_v_r_489_sv2v_reg <= data_mem_data_lo[489];
      ld_data_v_r_488_sv2v_reg <= data_mem_data_lo[488];
      ld_data_v_r_487_sv2v_reg <= data_mem_data_lo[487];
      ld_data_v_r_486_sv2v_reg <= data_mem_data_lo[486];
      ld_data_v_r_485_sv2v_reg <= data_mem_data_lo[485];
      ld_data_v_r_484_sv2v_reg <= data_mem_data_lo[484];
      ld_data_v_r_483_sv2v_reg <= data_mem_data_lo[483];
      ld_data_v_r_482_sv2v_reg <= data_mem_data_lo[482];
      ld_data_v_r_481_sv2v_reg <= data_mem_data_lo[481];
      ld_data_v_r_480_sv2v_reg <= data_mem_data_lo[480];
      ld_data_v_r_479_sv2v_reg <= data_mem_data_lo[479];
      ld_data_v_r_478_sv2v_reg <= data_mem_data_lo[478];
      ld_data_v_r_477_sv2v_reg <= data_mem_data_lo[477];
      ld_data_v_r_476_sv2v_reg <= data_mem_data_lo[476];
      ld_data_v_r_475_sv2v_reg <= data_mem_data_lo[475];
      ld_data_v_r_474_sv2v_reg <= data_mem_data_lo[474];
      ld_data_v_r_473_sv2v_reg <= data_mem_data_lo[473];
      ld_data_v_r_472_sv2v_reg <= data_mem_data_lo[472];
      ld_data_v_r_471_sv2v_reg <= data_mem_data_lo[471];
      ld_data_v_r_470_sv2v_reg <= data_mem_data_lo[470];
      ld_data_v_r_469_sv2v_reg <= data_mem_data_lo[469];
      ld_data_v_r_468_sv2v_reg <= data_mem_data_lo[468];
      ld_data_v_r_467_sv2v_reg <= data_mem_data_lo[467];
      ld_data_v_r_466_sv2v_reg <= data_mem_data_lo[466];
      ld_data_v_r_465_sv2v_reg <= data_mem_data_lo[465];
      ld_data_v_r_464_sv2v_reg <= data_mem_data_lo[464];
      ld_data_v_r_463_sv2v_reg <= data_mem_data_lo[463];
      ld_data_v_r_462_sv2v_reg <= data_mem_data_lo[462];
    end 
    if(N108) begin
      ld_data_v_r_461_sv2v_reg <= data_mem_data_lo[461];
      ld_data_v_r_460_sv2v_reg <= data_mem_data_lo[460];
      ld_data_v_r_459_sv2v_reg <= data_mem_data_lo[459];
      ld_data_v_r_458_sv2v_reg <= data_mem_data_lo[458];
      ld_data_v_r_457_sv2v_reg <= data_mem_data_lo[457];
      ld_data_v_r_456_sv2v_reg <= data_mem_data_lo[456];
      ld_data_v_r_455_sv2v_reg <= data_mem_data_lo[455];
      ld_data_v_r_454_sv2v_reg <= data_mem_data_lo[454];
      ld_data_v_r_453_sv2v_reg <= data_mem_data_lo[453];
      ld_data_v_r_452_sv2v_reg <= data_mem_data_lo[452];
      ld_data_v_r_451_sv2v_reg <= data_mem_data_lo[451];
      ld_data_v_r_450_sv2v_reg <= data_mem_data_lo[450];
      ld_data_v_r_449_sv2v_reg <= data_mem_data_lo[449];
      ld_data_v_r_448_sv2v_reg <= data_mem_data_lo[448];
      ld_data_v_r_447_sv2v_reg <= data_mem_data_lo[447];
      ld_data_v_r_446_sv2v_reg <= data_mem_data_lo[446];
      ld_data_v_r_445_sv2v_reg <= data_mem_data_lo[445];
      ld_data_v_r_444_sv2v_reg <= data_mem_data_lo[444];
      ld_data_v_r_443_sv2v_reg <= data_mem_data_lo[443];
      ld_data_v_r_442_sv2v_reg <= data_mem_data_lo[442];
      ld_data_v_r_441_sv2v_reg <= data_mem_data_lo[441];
      ld_data_v_r_440_sv2v_reg <= data_mem_data_lo[440];
      ld_data_v_r_439_sv2v_reg <= data_mem_data_lo[439];
      ld_data_v_r_438_sv2v_reg <= data_mem_data_lo[438];
      ld_data_v_r_437_sv2v_reg <= data_mem_data_lo[437];
      ld_data_v_r_436_sv2v_reg <= data_mem_data_lo[436];
      ld_data_v_r_435_sv2v_reg <= data_mem_data_lo[435];
      ld_data_v_r_434_sv2v_reg <= data_mem_data_lo[434];
      ld_data_v_r_433_sv2v_reg <= data_mem_data_lo[433];
      ld_data_v_r_432_sv2v_reg <= data_mem_data_lo[432];
      ld_data_v_r_431_sv2v_reg <= data_mem_data_lo[431];
      ld_data_v_r_430_sv2v_reg <= data_mem_data_lo[430];
      ld_data_v_r_429_sv2v_reg <= data_mem_data_lo[429];
      ld_data_v_r_428_sv2v_reg <= data_mem_data_lo[428];
      ld_data_v_r_427_sv2v_reg <= data_mem_data_lo[427];
      ld_data_v_r_426_sv2v_reg <= data_mem_data_lo[426];
      ld_data_v_r_425_sv2v_reg <= data_mem_data_lo[425];
      ld_data_v_r_424_sv2v_reg <= data_mem_data_lo[424];
      ld_data_v_r_423_sv2v_reg <= data_mem_data_lo[423];
      ld_data_v_r_422_sv2v_reg <= data_mem_data_lo[422];
      ld_data_v_r_421_sv2v_reg <= data_mem_data_lo[421];
      ld_data_v_r_420_sv2v_reg <= data_mem_data_lo[420];
      ld_data_v_r_419_sv2v_reg <= data_mem_data_lo[419];
      ld_data_v_r_418_sv2v_reg <= data_mem_data_lo[418];
      ld_data_v_r_417_sv2v_reg <= data_mem_data_lo[417];
      ld_data_v_r_416_sv2v_reg <= data_mem_data_lo[416];
      ld_data_v_r_415_sv2v_reg <= data_mem_data_lo[415];
      ld_data_v_r_414_sv2v_reg <= data_mem_data_lo[414];
      ld_data_v_r_413_sv2v_reg <= data_mem_data_lo[413];
      ld_data_v_r_412_sv2v_reg <= data_mem_data_lo[412];
      ld_data_v_r_411_sv2v_reg <= data_mem_data_lo[411];
      ld_data_v_r_410_sv2v_reg <= data_mem_data_lo[410];
      ld_data_v_r_409_sv2v_reg <= data_mem_data_lo[409];
      ld_data_v_r_408_sv2v_reg <= data_mem_data_lo[408];
      ld_data_v_r_407_sv2v_reg <= data_mem_data_lo[407];
      ld_data_v_r_406_sv2v_reg <= data_mem_data_lo[406];
      ld_data_v_r_405_sv2v_reg <= data_mem_data_lo[405];
      ld_data_v_r_404_sv2v_reg <= data_mem_data_lo[404];
      ld_data_v_r_403_sv2v_reg <= data_mem_data_lo[403];
      ld_data_v_r_402_sv2v_reg <= data_mem_data_lo[402];
      ld_data_v_r_401_sv2v_reg <= data_mem_data_lo[401];
      ld_data_v_r_400_sv2v_reg <= data_mem_data_lo[400];
      ld_data_v_r_399_sv2v_reg <= data_mem_data_lo[399];
      ld_data_v_r_398_sv2v_reg <= data_mem_data_lo[398];
      ld_data_v_r_397_sv2v_reg <= data_mem_data_lo[397];
      ld_data_v_r_396_sv2v_reg <= data_mem_data_lo[396];
      ld_data_v_r_395_sv2v_reg <= data_mem_data_lo[395];
      ld_data_v_r_394_sv2v_reg <= data_mem_data_lo[394];
      ld_data_v_r_393_sv2v_reg <= data_mem_data_lo[393];
      ld_data_v_r_392_sv2v_reg <= data_mem_data_lo[392];
      ld_data_v_r_391_sv2v_reg <= data_mem_data_lo[391];
      ld_data_v_r_390_sv2v_reg <= data_mem_data_lo[390];
      ld_data_v_r_389_sv2v_reg <= data_mem_data_lo[389];
      ld_data_v_r_388_sv2v_reg <= data_mem_data_lo[388];
      ld_data_v_r_387_sv2v_reg <= data_mem_data_lo[387];
      ld_data_v_r_386_sv2v_reg <= data_mem_data_lo[386];
      ld_data_v_r_385_sv2v_reg <= data_mem_data_lo[385];
      ld_data_v_r_384_sv2v_reg <= data_mem_data_lo[384];
      ld_data_v_r_383_sv2v_reg <= data_mem_data_lo[383];
      ld_data_v_r_382_sv2v_reg <= data_mem_data_lo[382];
      ld_data_v_r_381_sv2v_reg <= data_mem_data_lo[381];
      ld_data_v_r_380_sv2v_reg <= data_mem_data_lo[380];
      ld_data_v_r_379_sv2v_reg <= data_mem_data_lo[379];
      ld_data_v_r_378_sv2v_reg <= data_mem_data_lo[378];
      ld_data_v_r_377_sv2v_reg <= data_mem_data_lo[377];
      ld_data_v_r_376_sv2v_reg <= data_mem_data_lo[376];
      ld_data_v_r_375_sv2v_reg <= data_mem_data_lo[375];
      ld_data_v_r_374_sv2v_reg <= data_mem_data_lo[374];
      ld_data_v_r_373_sv2v_reg <= data_mem_data_lo[373];
      ld_data_v_r_372_sv2v_reg <= data_mem_data_lo[372];
      ld_data_v_r_371_sv2v_reg <= data_mem_data_lo[371];
      ld_data_v_r_370_sv2v_reg <= data_mem_data_lo[370];
      ld_data_v_r_369_sv2v_reg <= data_mem_data_lo[369];
      ld_data_v_r_368_sv2v_reg <= data_mem_data_lo[368];
      ld_data_v_r_367_sv2v_reg <= data_mem_data_lo[367];
      ld_data_v_r_366_sv2v_reg <= data_mem_data_lo[366];
      ld_data_v_r_365_sv2v_reg <= data_mem_data_lo[365];
      ld_data_v_r_364_sv2v_reg <= data_mem_data_lo[364];
      ld_data_v_r_363_sv2v_reg <= data_mem_data_lo[363];
    end 
    if(N107) begin
      ld_data_v_r_362_sv2v_reg <= data_mem_data_lo[362];
      ld_data_v_r_361_sv2v_reg <= data_mem_data_lo[361];
      ld_data_v_r_360_sv2v_reg <= data_mem_data_lo[360];
      ld_data_v_r_359_sv2v_reg <= data_mem_data_lo[359];
      ld_data_v_r_358_sv2v_reg <= data_mem_data_lo[358];
      ld_data_v_r_357_sv2v_reg <= data_mem_data_lo[357];
      ld_data_v_r_356_sv2v_reg <= data_mem_data_lo[356];
      ld_data_v_r_355_sv2v_reg <= data_mem_data_lo[355];
      ld_data_v_r_354_sv2v_reg <= data_mem_data_lo[354];
      ld_data_v_r_353_sv2v_reg <= data_mem_data_lo[353];
      ld_data_v_r_352_sv2v_reg <= data_mem_data_lo[352];
      ld_data_v_r_351_sv2v_reg <= data_mem_data_lo[351];
      ld_data_v_r_350_sv2v_reg <= data_mem_data_lo[350];
      ld_data_v_r_349_sv2v_reg <= data_mem_data_lo[349];
      ld_data_v_r_348_sv2v_reg <= data_mem_data_lo[348];
      ld_data_v_r_347_sv2v_reg <= data_mem_data_lo[347];
      ld_data_v_r_346_sv2v_reg <= data_mem_data_lo[346];
      ld_data_v_r_345_sv2v_reg <= data_mem_data_lo[345];
      ld_data_v_r_344_sv2v_reg <= data_mem_data_lo[344];
      ld_data_v_r_343_sv2v_reg <= data_mem_data_lo[343];
      ld_data_v_r_342_sv2v_reg <= data_mem_data_lo[342];
      ld_data_v_r_341_sv2v_reg <= data_mem_data_lo[341];
      ld_data_v_r_340_sv2v_reg <= data_mem_data_lo[340];
      ld_data_v_r_339_sv2v_reg <= data_mem_data_lo[339];
      ld_data_v_r_338_sv2v_reg <= data_mem_data_lo[338];
      ld_data_v_r_337_sv2v_reg <= data_mem_data_lo[337];
      ld_data_v_r_336_sv2v_reg <= data_mem_data_lo[336];
      ld_data_v_r_335_sv2v_reg <= data_mem_data_lo[335];
      ld_data_v_r_334_sv2v_reg <= data_mem_data_lo[334];
      ld_data_v_r_333_sv2v_reg <= data_mem_data_lo[333];
      ld_data_v_r_332_sv2v_reg <= data_mem_data_lo[332];
      ld_data_v_r_331_sv2v_reg <= data_mem_data_lo[331];
      ld_data_v_r_330_sv2v_reg <= data_mem_data_lo[330];
      ld_data_v_r_329_sv2v_reg <= data_mem_data_lo[329];
      ld_data_v_r_328_sv2v_reg <= data_mem_data_lo[328];
      ld_data_v_r_327_sv2v_reg <= data_mem_data_lo[327];
      ld_data_v_r_326_sv2v_reg <= data_mem_data_lo[326];
      ld_data_v_r_325_sv2v_reg <= data_mem_data_lo[325];
      ld_data_v_r_324_sv2v_reg <= data_mem_data_lo[324];
      ld_data_v_r_323_sv2v_reg <= data_mem_data_lo[323];
      ld_data_v_r_322_sv2v_reg <= data_mem_data_lo[322];
      ld_data_v_r_321_sv2v_reg <= data_mem_data_lo[321];
      ld_data_v_r_320_sv2v_reg <= data_mem_data_lo[320];
      ld_data_v_r_319_sv2v_reg <= data_mem_data_lo[319];
      ld_data_v_r_318_sv2v_reg <= data_mem_data_lo[318];
      ld_data_v_r_317_sv2v_reg <= data_mem_data_lo[317];
      ld_data_v_r_316_sv2v_reg <= data_mem_data_lo[316];
      ld_data_v_r_315_sv2v_reg <= data_mem_data_lo[315];
      ld_data_v_r_314_sv2v_reg <= data_mem_data_lo[314];
      ld_data_v_r_313_sv2v_reg <= data_mem_data_lo[313];
      ld_data_v_r_312_sv2v_reg <= data_mem_data_lo[312];
      ld_data_v_r_311_sv2v_reg <= data_mem_data_lo[311];
      ld_data_v_r_310_sv2v_reg <= data_mem_data_lo[310];
      ld_data_v_r_309_sv2v_reg <= data_mem_data_lo[309];
      ld_data_v_r_308_sv2v_reg <= data_mem_data_lo[308];
      ld_data_v_r_307_sv2v_reg <= data_mem_data_lo[307];
      ld_data_v_r_306_sv2v_reg <= data_mem_data_lo[306];
      ld_data_v_r_305_sv2v_reg <= data_mem_data_lo[305];
      ld_data_v_r_304_sv2v_reg <= data_mem_data_lo[304];
      ld_data_v_r_303_sv2v_reg <= data_mem_data_lo[303];
      ld_data_v_r_302_sv2v_reg <= data_mem_data_lo[302];
      ld_data_v_r_301_sv2v_reg <= data_mem_data_lo[301];
      ld_data_v_r_300_sv2v_reg <= data_mem_data_lo[300];
      ld_data_v_r_299_sv2v_reg <= data_mem_data_lo[299];
      ld_data_v_r_298_sv2v_reg <= data_mem_data_lo[298];
      ld_data_v_r_297_sv2v_reg <= data_mem_data_lo[297];
      ld_data_v_r_296_sv2v_reg <= data_mem_data_lo[296];
      ld_data_v_r_295_sv2v_reg <= data_mem_data_lo[295];
      ld_data_v_r_294_sv2v_reg <= data_mem_data_lo[294];
      ld_data_v_r_293_sv2v_reg <= data_mem_data_lo[293];
      ld_data_v_r_292_sv2v_reg <= data_mem_data_lo[292];
      ld_data_v_r_291_sv2v_reg <= data_mem_data_lo[291];
      ld_data_v_r_290_sv2v_reg <= data_mem_data_lo[290];
      ld_data_v_r_289_sv2v_reg <= data_mem_data_lo[289];
      ld_data_v_r_288_sv2v_reg <= data_mem_data_lo[288];
      ld_data_v_r_287_sv2v_reg <= data_mem_data_lo[287];
      ld_data_v_r_286_sv2v_reg <= data_mem_data_lo[286];
      ld_data_v_r_285_sv2v_reg <= data_mem_data_lo[285];
      ld_data_v_r_284_sv2v_reg <= data_mem_data_lo[284];
      ld_data_v_r_283_sv2v_reg <= data_mem_data_lo[283];
      ld_data_v_r_282_sv2v_reg <= data_mem_data_lo[282];
      ld_data_v_r_281_sv2v_reg <= data_mem_data_lo[281];
      ld_data_v_r_280_sv2v_reg <= data_mem_data_lo[280];
      ld_data_v_r_279_sv2v_reg <= data_mem_data_lo[279];
      ld_data_v_r_278_sv2v_reg <= data_mem_data_lo[278];
      ld_data_v_r_277_sv2v_reg <= data_mem_data_lo[277];
      ld_data_v_r_276_sv2v_reg <= data_mem_data_lo[276];
      ld_data_v_r_275_sv2v_reg <= data_mem_data_lo[275];
      ld_data_v_r_274_sv2v_reg <= data_mem_data_lo[274];
      ld_data_v_r_273_sv2v_reg <= data_mem_data_lo[273];
      ld_data_v_r_272_sv2v_reg <= data_mem_data_lo[272];
      ld_data_v_r_271_sv2v_reg <= data_mem_data_lo[271];
      ld_data_v_r_270_sv2v_reg <= data_mem_data_lo[270];
      ld_data_v_r_269_sv2v_reg <= data_mem_data_lo[269];
      ld_data_v_r_268_sv2v_reg <= data_mem_data_lo[268];
      ld_data_v_r_267_sv2v_reg <= data_mem_data_lo[267];
      ld_data_v_r_266_sv2v_reg <= data_mem_data_lo[266];
      ld_data_v_r_265_sv2v_reg <= data_mem_data_lo[265];
      ld_data_v_r_264_sv2v_reg <= data_mem_data_lo[264];
    end 
    if(N106) begin
      ld_data_v_r_263_sv2v_reg <= data_mem_data_lo[263];
      ld_data_v_r_262_sv2v_reg <= data_mem_data_lo[262];
      ld_data_v_r_261_sv2v_reg <= data_mem_data_lo[261];
      ld_data_v_r_260_sv2v_reg <= data_mem_data_lo[260];
      ld_data_v_r_259_sv2v_reg <= data_mem_data_lo[259];
      ld_data_v_r_258_sv2v_reg <= data_mem_data_lo[258];
      ld_data_v_r_257_sv2v_reg <= data_mem_data_lo[257];
      ld_data_v_r_256_sv2v_reg <= data_mem_data_lo[256];
      ld_data_v_r_255_sv2v_reg <= data_mem_data_lo[255];
      ld_data_v_r_254_sv2v_reg <= data_mem_data_lo[254];
      ld_data_v_r_253_sv2v_reg <= data_mem_data_lo[253];
      ld_data_v_r_252_sv2v_reg <= data_mem_data_lo[252];
      ld_data_v_r_251_sv2v_reg <= data_mem_data_lo[251];
      ld_data_v_r_250_sv2v_reg <= data_mem_data_lo[250];
      ld_data_v_r_249_sv2v_reg <= data_mem_data_lo[249];
      ld_data_v_r_248_sv2v_reg <= data_mem_data_lo[248];
      ld_data_v_r_247_sv2v_reg <= data_mem_data_lo[247];
      ld_data_v_r_246_sv2v_reg <= data_mem_data_lo[246];
      ld_data_v_r_245_sv2v_reg <= data_mem_data_lo[245];
      ld_data_v_r_244_sv2v_reg <= data_mem_data_lo[244];
      ld_data_v_r_243_sv2v_reg <= data_mem_data_lo[243];
      ld_data_v_r_242_sv2v_reg <= data_mem_data_lo[242];
      ld_data_v_r_241_sv2v_reg <= data_mem_data_lo[241];
      ld_data_v_r_240_sv2v_reg <= data_mem_data_lo[240];
      ld_data_v_r_239_sv2v_reg <= data_mem_data_lo[239];
      ld_data_v_r_238_sv2v_reg <= data_mem_data_lo[238];
      ld_data_v_r_237_sv2v_reg <= data_mem_data_lo[237];
      ld_data_v_r_236_sv2v_reg <= data_mem_data_lo[236];
      ld_data_v_r_235_sv2v_reg <= data_mem_data_lo[235];
      ld_data_v_r_234_sv2v_reg <= data_mem_data_lo[234];
      ld_data_v_r_233_sv2v_reg <= data_mem_data_lo[233];
      ld_data_v_r_232_sv2v_reg <= data_mem_data_lo[232];
      ld_data_v_r_231_sv2v_reg <= data_mem_data_lo[231];
      ld_data_v_r_230_sv2v_reg <= data_mem_data_lo[230];
      ld_data_v_r_229_sv2v_reg <= data_mem_data_lo[229];
      ld_data_v_r_228_sv2v_reg <= data_mem_data_lo[228];
      ld_data_v_r_227_sv2v_reg <= data_mem_data_lo[227];
      ld_data_v_r_226_sv2v_reg <= data_mem_data_lo[226];
      ld_data_v_r_225_sv2v_reg <= data_mem_data_lo[225];
      ld_data_v_r_224_sv2v_reg <= data_mem_data_lo[224];
      ld_data_v_r_223_sv2v_reg <= data_mem_data_lo[223];
      ld_data_v_r_222_sv2v_reg <= data_mem_data_lo[222];
      ld_data_v_r_221_sv2v_reg <= data_mem_data_lo[221];
      ld_data_v_r_220_sv2v_reg <= data_mem_data_lo[220];
      ld_data_v_r_219_sv2v_reg <= data_mem_data_lo[219];
      ld_data_v_r_218_sv2v_reg <= data_mem_data_lo[218];
      ld_data_v_r_217_sv2v_reg <= data_mem_data_lo[217];
      ld_data_v_r_216_sv2v_reg <= data_mem_data_lo[216];
      ld_data_v_r_215_sv2v_reg <= data_mem_data_lo[215];
      ld_data_v_r_214_sv2v_reg <= data_mem_data_lo[214];
      ld_data_v_r_213_sv2v_reg <= data_mem_data_lo[213];
      ld_data_v_r_212_sv2v_reg <= data_mem_data_lo[212];
      ld_data_v_r_211_sv2v_reg <= data_mem_data_lo[211];
      ld_data_v_r_210_sv2v_reg <= data_mem_data_lo[210];
      ld_data_v_r_209_sv2v_reg <= data_mem_data_lo[209];
      ld_data_v_r_208_sv2v_reg <= data_mem_data_lo[208];
      ld_data_v_r_207_sv2v_reg <= data_mem_data_lo[207];
      ld_data_v_r_206_sv2v_reg <= data_mem_data_lo[206];
      ld_data_v_r_205_sv2v_reg <= data_mem_data_lo[205];
      ld_data_v_r_204_sv2v_reg <= data_mem_data_lo[204];
      ld_data_v_r_203_sv2v_reg <= data_mem_data_lo[203];
      ld_data_v_r_202_sv2v_reg <= data_mem_data_lo[202];
      ld_data_v_r_201_sv2v_reg <= data_mem_data_lo[201];
      ld_data_v_r_200_sv2v_reg <= data_mem_data_lo[200];
      ld_data_v_r_199_sv2v_reg <= data_mem_data_lo[199];
      ld_data_v_r_198_sv2v_reg <= data_mem_data_lo[198];
      ld_data_v_r_197_sv2v_reg <= data_mem_data_lo[197];
      ld_data_v_r_196_sv2v_reg <= data_mem_data_lo[196];
      ld_data_v_r_195_sv2v_reg <= data_mem_data_lo[195];
      ld_data_v_r_194_sv2v_reg <= data_mem_data_lo[194];
      ld_data_v_r_193_sv2v_reg <= data_mem_data_lo[193];
      ld_data_v_r_192_sv2v_reg <= data_mem_data_lo[192];
      ld_data_v_r_191_sv2v_reg <= data_mem_data_lo[191];
      ld_data_v_r_190_sv2v_reg <= data_mem_data_lo[190];
      ld_data_v_r_189_sv2v_reg <= data_mem_data_lo[189];
      ld_data_v_r_188_sv2v_reg <= data_mem_data_lo[188];
      ld_data_v_r_187_sv2v_reg <= data_mem_data_lo[187];
      ld_data_v_r_186_sv2v_reg <= data_mem_data_lo[186];
      ld_data_v_r_185_sv2v_reg <= data_mem_data_lo[185];
      ld_data_v_r_184_sv2v_reg <= data_mem_data_lo[184];
      ld_data_v_r_183_sv2v_reg <= data_mem_data_lo[183];
      ld_data_v_r_182_sv2v_reg <= data_mem_data_lo[182];
      ld_data_v_r_181_sv2v_reg <= data_mem_data_lo[181];
      ld_data_v_r_180_sv2v_reg <= data_mem_data_lo[180];
      ld_data_v_r_179_sv2v_reg <= data_mem_data_lo[179];
      ld_data_v_r_178_sv2v_reg <= data_mem_data_lo[178];
      ld_data_v_r_177_sv2v_reg <= data_mem_data_lo[177];
      ld_data_v_r_176_sv2v_reg <= data_mem_data_lo[176];
      ld_data_v_r_175_sv2v_reg <= data_mem_data_lo[175];
      ld_data_v_r_174_sv2v_reg <= data_mem_data_lo[174];
      ld_data_v_r_173_sv2v_reg <= data_mem_data_lo[173];
      ld_data_v_r_172_sv2v_reg <= data_mem_data_lo[172];
      ld_data_v_r_171_sv2v_reg <= data_mem_data_lo[171];
      ld_data_v_r_170_sv2v_reg <= data_mem_data_lo[170];
      ld_data_v_r_169_sv2v_reg <= data_mem_data_lo[169];
      ld_data_v_r_168_sv2v_reg <= data_mem_data_lo[168];
      ld_data_v_r_167_sv2v_reg <= data_mem_data_lo[167];
      ld_data_v_r_166_sv2v_reg <= data_mem_data_lo[166];
      ld_data_v_r_165_sv2v_reg <= data_mem_data_lo[165];
    end 
    if(N105) begin
      ld_data_v_r_164_sv2v_reg <= data_mem_data_lo[164];
      ld_data_v_r_163_sv2v_reg <= data_mem_data_lo[163];
      ld_data_v_r_162_sv2v_reg <= data_mem_data_lo[162];
      ld_data_v_r_161_sv2v_reg <= data_mem_data_lo[161];
      ld_data_v_r_160_sv2v_reg <= data_mem_data_lo[160];
      ld_data_v_r_159_sv2v_reg <= data_mem_data_lo[159];
      ld_data_v_r_158_sv2v_reg <= data_mem_data_lo[158];
      ld_data_v_r_157_sv2v_reg <= data_mem_data_lo[157];
      ld_data_v_r_156_sv2v_reg <= data_mem_data_lo[156];
      ld_data_v_r_155_sv2v_reg <= data_mem_data_lo[155];
      ld_data_v_r_154_sv2v_reg <= data_mem_data_lo[154];
      ld_data_v_r_153_sv2v_reg <= data_mem_data_lo[153];
      ld_data_v_r_152_sv2v_reg <= data_mem_data_lo[152];
      ld_data_v_r_151_sv2v_reg <= data_mem_data_lo[151];
      ld_data_v_r_150_sv2v_reg <= data_mem_data_lo[150];
      ld_data_v_r_149_sv2v_reg <= data_mem_data_lo[149];
      ld_data_v_r_148_sv2v_reg <= data_mem_data_lo[148];
      ld_data_v_r_147_sv2v_reg <= data_mem_data_lo[147];
      ld_data_v_r_146_sv2v_reg <= data_mem_data_lo[146];
      ld_data_v_r_145_sv2v_reg <= data_mem_data_lo[145];
      ld_data_v_r_144_sv2v_reg <= data_mem_data_lo[144];
      ld_data_v_r_143_sv2v_reg <= data_mem_data_lo[143];
      ld_data_v_r_142_sv2v_reg <= data_mem_data_lo[142];
      ld_data_v_r_141_sv2v_reg <= data_mem_data_lo[141];
      ld_data_v_r_140_sv2v_reg <= data_mem_data_lo[140];
      ld_data_v_r_139_sv2v_reg <= data_mem_data_lo[139];
      ld_data_v_r_138_sv2v_reg <= data_mem_data_lo[138];
      ld_data_v_r_137_sv2v_reg <= data_mem_data_lo[137];
      ld_data_v_r_136_sv2v_reg <= data_mem_data_lo[136];
      ld_data_v_r_135_sv2v_reg <= data_mem_data_lo[135];
      ld_data_v_r_134_sv2v_reg <= data_mem_data_lo[134];
      ld_data_v_r_133_sv2v_reg <= data_mem_data_lo[133];
      ld_data_v_r_132_sv2v_reg <= data_mem_data_lo[132];
      ld_data_v_r_131_sv2v_reg <= data_mem_data_lo[131];
      ld_data_v_r_130_sv2v_reg <= data_mem_data_lo[130];
      ld_data_v_r_129_sv2v_reg <= data_mem_data_lo[129];
      ld_data_v_r_128_sv2v_reg <= data_mem_data_lo[128];
      ld_data_v_r_127_sv2v_reg <= data_mem_data_lo[127];
      ld_data_v_r_126_sv2v_reg <= data_mem_data_lo[126];
      ld_data_v_r_125_sv2v_reg <= data_mem_data_lo[125];
      ld_data_v_r_124_sv2v_reg <= data_mem_data_lo[124];
      ld_data_v_r_123_sv2v_reg <= data_mem_data_lo[123];
      ld_data_v_r_122_sv2v_reg <= data_mem_data_lo[122];
      ld_data_v_r_121_sv2v_reg <= data_mem_data_lo[121];
      ld_data_v_r_120_sv2v_reg <= data_mem_data_lo[120];
      ld_data_v_r_119_sv2v_reg <= data_mem_data_lo[119];
      ld_data_v_r_118_sv2v_reg <= data_mem_data_lo[118];
      ld_data_v_r_117_sv2v_reg <= data_mem_data_lo[117];
      ld_data_v_r_116_sv2v_reg <= data_mem_data_lo[116];
      ld_data_v_r_115_sv2v_reg <= data_mem_data_lo[115];
      ld_data_v_r_114_sv2v_reg <= data_mem_data_lo[114];
      ld_data_v_r_113_sv2v_reg <= data_mem_data_lo[113];
      ld_data_v_r_112_sv2v_reg <= data_mem_data_lo[112];
      ld_data_v_r_111_sv2v_reg <= data_mem_data_lo[111];
      ld_data_v_r_110_sv2v_reg <= data_mem_data_lo[110];
      ld_data_v_r_109_sv2v_reg <= data_mem_data_lo[109];
      ld_data_v_r_108_sv2v_reg <= data_mem_data_lo[108];
      ld_data_v_r_107_sv2v_reg <= data_mem_data_lo[107];
      ld_data_v_r_106_sv2v_reg <= data_mem_data_lo[106];
      ld_data_v_r_105_sv2v_reg <= data_mem_data_lo[105];
      ld_data_v_r_104_sv2v_reg <= data_mem_data_lo[104];
      ld_data_v_r_103_sv2v_reg <= data_mem_data_lo[103];
      ld_data_v_r_102_sv2v_reg <= data_mem_data_lo[102];
      ld_data_v_r_101_sv2v_reg <= data_mem_data_lo[101];
      ld_data_v_r_100_sv2v_reg <= data_mem_data_lo[100];
      ld_data_v_r_99_sv2v_reg <= data_mem_data_lo[99];
      ld_data_v_r_98_sv2v_reg <= data_mem_data_lo[98];
      ld_data_v_r_97_sv2v_reg <= data_mem_data_lo[97];
      ld_data_v_r_96_sv2v_reg <= data_mem_data_lo[96];
      ld_data_v_r_95_sv2v_reg <= data_mem_data_lo[95];
      ld_data_v_r_94_sv2v_reg <= data_mem_data_lo[94];
      ld_data_v_r_93_sv2v_reg <= data_mem_data_lo[93];
      ld_data_v_r_92_sv2v_reg <= data_mem_data_lo[92];
      ld_data_v_r_91_sv2v_reg <= data_mem_data_lo[91];
      ld_data_v_r_90_sv2v_reg <= data_mem_data_lo[90];
      ld_data_v_r_89_sv2v_reg <= data_mem_data_lo[89];
      ld_data_v_r_88_sv2v_reg <= data_mem_data_lo[88];
      ld_data_v_r_87_sv2v_reg <= data_mem_data_lo[87];
      ld_data_v_r_86_sv2v_reg <= data_mem_data_lo[86];
      ld_data_v_r_85_sv2v_reg <= data_mem_data_lo[85];
      ld_data_v_r_84_sv2v_reg <= data_mem_data_lo[84];
      ld_data_v_r_83_sv2v_reg <= data_mem_data_lo[83];
      ld_data_v_r_82_sv2v_reg <= data_mem_data_lo[82];
      ld_data_v_r_81_sv2v_reg <= data_mem_data_lo[81];
      ld_data_v_r_80_sv2v_reg <= data_mem_data_lo[80];
      ld_data_v_r_79_sv2v_reg <= data_mem_data_lo[79];
      ld_data_v_r_78_sv2v_reg <= data_mem_data_lo[78];
      ld_data_v_r_77_sv2v_reg <= data_mem_data_lo[77];
      ld_data_v_r_76_sv2v_reg <= data_mem_data_lo[76];
      ld_data_v_r_75_sv2v_reg <= data_mem_data_lo[75];
      ld_data_v_r_74_sv2v_reg <= data_mem_data_lo[74];
      ld_data_v_r_73_sv2v_reg <= data_mem_data_lo[73];
      ld_data_v_r_72_sv2v_reg <= data_mem_data_lo[72];
      ld_data_v_r_71_sv2v_reg <= data_mem_data_lo[71];
      ld_data_v_r_70_sv2v_reg <= data_mem_data_lo[70];
      ld_data_v_r_69_sv2v_reg <= data_mem_data_lo[69];
      ld_data_v_r_68_sv2v_reg <= data_mem_data_lo[68];
      ld_data_v_r_67_sv2v_reg <= data_mem_data_lo[67];
      ld_data_v_r_66_sv2v_reg <= data_mem_data_lo[66];
    end 
    if(N104) begin
      ld_data_v_r_65_sv2v_reg <= data_mem_data_lo[65];
      ld_data_v_r_64_sv2v_reg <= data_mem_data_lo[64];
      ld_data_v_r_63_sv2v_reg <= data_mem_data_lo[63];
      ld_data_v_r_62_sv2v_reg <= data_mem_data_lo[62];
      ld_data_v_r_61_sv2v_reg <= data_mem_data_lo[61];
      ld_data_v_r_60_sv2v_reg <= data_mem_data_lo[60];
      ld_data_v_r_59_sv2v_reg <= data_mem_data_lo[59];
      ld_data_v_r_58_sv2v_reg <= data_mem_data_lo[58];
      ld_data_v_r_57_sv2v_reg <= data_mem_data_lo[57];
      ld_data_v_r_56_sv2v_reg <= data_mem_data_lo[56];
      ld_data_v_r_55_sv2v_reg <= data_mem_data_lo[55];
      ld_data_v_r_54_sv2v_reg <= data_mem_data_lo[54];
      ld_data_v_r_53_sv2v_reg <= data_mem_data_lo[53];
      ld_data_v_r_52_sv2v_reg <= data_mem_data_lo[52];
      ld_data_v_r_51_sv2v_reg <= data_mem_data_lo[51];
      ld_data_v_r_50_sv2v_reg <= data_mem_data_lo[50];
      ld_data_v_r_49_sv2v_reg <= data_mem_data_lo[49];
      ld_data_v_r_48_sv2v_reg <= data_mem_data_lo[48];
      ld_data_v_r_47_sv2v_reg <= data_mem_data_lo[47];
      ld_data_v_r_46_sv2v_reg <= data_mem_data_lo[46];
      ld_data_v_r_45_sv2v_reg <= data_mem_data_lo[45];
      ld_data_v_r_44_sv2v_reg <= data_mem_data_lo[44];
      ld_data_v_r_43_sv2v_reg <= data_mem_data_lo[43];
      ld_data_v_r_42_sv2v_reg <= data_mem_data_lo[42];
      ld_data_v_r_41_sv2v_reg <= data_mem_data_lo[41];
      ld_data_v_r_40_sv2v_reg <= data_mem_data_lo[40];
      ld_data_v_r_39_sv2v_reg <= data_mem_data_lo[39];
      ld_data_v_r_38_sv2v_reg <= data_mem_data_lo[38];
      ld_data_v_r_37_sv2v_reg <= data_mem_data_lo[37];
      ld_data_v_r_36_sv2v_reg <= data_mem_data_lo[36];
      ld_data_v_r_35_sv2v_reg <= data_mem_data_lo[35];
      ld_data_v_r_34_sv2v_reg <= data_mem_data_lo[34];
      ld_data_v_r_33_sv2v_reg <= data_mem_data_lo[33];
      ld_data_v_r_32_sv2v_reg <= data_mem_data_lo[32];
      ld_data_v_r_31_sv2v_reg <= data_mem_data_lo[31];
      ld_data_v_r_30_sv2v_reg <= data_mem_data_lo[30];
      ld_data_v_r_29_sv2v_reg <= data_mem_data_lo[29];
      ld_data_v_r_28_sv2v_reg <= data_mem_data_lo[28];
      ld_data_v_r_27_sv2v_reg <= data_mem_data_lo[27];
      ld_data_v_r_26_sv2v_reg <= data_mem_data_lo[26];
      ld_data_v_r_25_sv2v_reg <= data_mem_data_lo[25];
      ld_data_v_r_24_sv2v_reg <= data_mem_data_lo[24];
      ld_data_v_r_23_sv2v_reg <= data_mem_data_lo[23];
      ld_data_v_r_22_sv2v_reg <= data_mem_data_lo[22];
      ld_data_v_r_21_sv2v_reg <= data_mem_data_lo[21];
      ld_data_v_r_20_sv2v_reg <= data_mem_data_lo[20];
      ld_data_v_r_19_sv2v_reg <= data_mem_data_lo[19];
      ld_data_v_r_18_sv2v_reg <= data_mem_data_lo[18];
      ld_data_v_r_17_sv2v_reg <= data_mem_data_lo[17];
      ld_data_v_r_16_sv2v_reg <= data_mem_data_lo[16];
      ld_data_v_r_15_sv2v_reg <= data_mem_data_lo[15];
      ld_data_v_r_14_sv2v_reg <= data_mem_data_lo[14];
      ld_data_v_r_13_sv2v_reg <= data_mem_data_lo[13];
      ld_data_v_r_12_sv2v_reg <= data_mem_data_lo[12];
      ld_data_v_r_11_sv2v_reg <= data_mem_data_lo[11];
      ld_data_v_r_10_sv2v_reg <= data_mem_data_lo[10];
      ld_data_v_r_9_sv2v_reg <= data_mem_data_lo[9];
      ld_data_v_r_8_sv2v_reg <= data_mem_data_lo[8];
      ld_data_v_r_7_sv2v_reg <= data_mem_data_lo[7];
      ld_data_v_r_6_sv2v_reg <= data_mem_data_lo[6];
      ld_data_v_r_5_sv2v_reg <= data_mem_data_lo[5];
      ld_data_v_r_4_sv2v_reg <= data_mem_data_lo[4];
      ld_data_v_r_3_sv2v_reg <= data_mem_data_lo[3];
      ld_data_v_r_2_sv2v_reg <= data_mem_data_lo[2];
      ld_data_v_r_1_sv2v_reg <= data_mem_data_lo[1];
      ld_data_v_r_0_sv2v_reg <= data_mem_data_lo[0];
    end 
    if(reset_i) begin
      v_v_r_sv2v_reg <= 1'b0;
    end else if(N88) begin
      v_v_r_sv2v_reg <= v_tl_r;
    end 
    if(reset_i) begin
      track_data_v_r_31_sv2v_reg <= 1'b0;
      track_data_v_r_30_sv2v_reg <= 1'b0;
      track_data_v_r_29_sv2v_reg <= 1'b0;
      track_data_v_r_28_sv2v_reg <= 1'b0;
      track_data_v_r_27_sv2v_reg <= 1'b0;
      track_data_v_r_26_sv2v_reg <= 1'b0;
      track_data_v_r_25_sv2v_reg <= 1'b0;
      track_data_v_r_24_sv2v_reg <= 1'b0;
      track_data_v_r_23_sv2v_reg <= 1'b0;
      track_data_v_r_22_sv2v_reg <= 1'b0;
      track_data_v_r_21_sv2v_reg <= 1'b0;
      track_data_v_r_20_sv2v_reg <= 1'b0;
      track_data_v_r_19_sv2v_reg <= 1'b0;
      track_data_v_r_18_sv2v_reg <= 1'b0;
      track_data_v_r_17_sv2v_reg <= 1'b0;
      track_data_v_r_16_sv2v_reg <= 1'b0;
      track_data_v_r_15_sv2v_reg <= 1'b0;
      track_data_v_r_14_sv2v_reg <= 1'b0;
      track_data_v_r_13_sv2v_reg <= 1'b0;
      track_data_v_r_12_sv2v_reg <= 1'b0;
      track_data_v_r_11_sv2v_reg <= 1'b0;
      track_data_v_r_10_sv2v_reg <= 1'b0;
      track_data_v_r_9_sv2v_reg <= 1'b0;
      track_data_v_r_8_sv2v_reg <= 1'b0;
      track_data_v_r_7_sv2v_reg <= 1'b0;
      track_data_v_r_6_sv2v_reg <= 1'b0;
      track_data_v_r_5_sv2v_reg <= 1'b0;
      track_data_v_r_4_sv2v_reg <= 1'b0;
      track_data_v_r_3_sv2v_reg <= 1'b0;
      track_data_v_r_2_sv2v_reg <= 1'b0;
      track_data_v_r_1_sv2v_reg <= 1'b0;
      track_data_v_r_0_sv2v_reg <= 1'b0;
      mask_v_r_0_sv2v_reg <= 1'b0;
    end else if(N89) begin
      track_data_v_r_31_sv2v_reg <= track_mem_data_lo[31];
      track_data_v_r_30_sv2v_reg <= track_mem_data_lo[30];
      track_data_v_r_29_sv2v_reg <= track_mem_data_lo[29];
      track_data_v_r_28_sv2v_reg <= track_mem_data_lo[28];
      track_data_v_r_27_sv2v_reg <= track_mem_data_lo[27];
      track_data_v_r_26_sv2v_reg <= track_mem_data_lo[26];
      track_data_v_r_25_sv2v_reg <= track_mem_data_lo[25];
      track_data_v_r_24_sv2v_reg <= track_mem_data_lo[24];
      track_data_v_r_23_sv2v_reg <= track_mem_data_lo[23];
      track_data_v_r_22_sv2v_reg <= track_mem_data_lo[22];
      track_data_v_r_21_sv2v_reg <= track_mem_data_lo[21];
      track_data_v_r_20_sv2v_reg <= track_mem_data_lo[20];
      track_data_v_r_19_sv2v_reg <= track_mem_data_lo[19];
      track_data_v_r_18_sv2v_reg <= track_mem_data_lo[18];
      track_data_v_r_17_sv2v_reg <= track_mem_data_lo[17];
      track_data_v_r_16_sv2v_reg <= track_mem_data_lo[16];
      track_data_v_r_15_sv2v_reg <= track_mem_data_lo[15];
      track_data_v_r_14_sv2v_reg <= track_mem_data_lo[14];
      track_data_v_r_13_sv2v_reg <= track_mem_data_lo[13];
      track_data_v_r_12_sv2v_reg <= track_mem_data_lo[12];
      track_data_v_r_11_sv2v_reg <= track_mem_data_lo[11];
      track_data_v_r_10_sv2v_reg <= track_mem_data_lo[10];
      track_data_v_r_9_sv2v_reg <= track_mem_data_lo[9];
      track_data_v_r_8_sv2v_reg <= track_mem_data_lo[8];
      track_data_v_r_7_sv2v_reg <= track_mem_data_lo[7];
      track_data_v_r_6_sv2v_reg <= track_mem_data_lo[6];
      track_data_v_r_5_sv2v_reg <= track_mem_data_lo[5];
      track_data_v_r_4_sv2v_reg <= track_mem_data_lo[4];
      track_data_v_r_3_sv2v_reg <= track_mem_data_lo[3];
      track_data_v_r_2_sv2v_reg <= track_mem_data_lo[2];
      track_data_v_r_1_sv2v_reg <= track_mem_data_lo[1];
      track_data_v_r_0_sv2v_reg <= track_mem_data_lo[0];
      mask_v_r_0_sv2v_reg <= mask_tl_r[0];
    end 
    if(reset_i) begin
      mask_v_r_15_sv2v_reg <= 1'b0;
      mask_v_r_14_sv2v_reg <= 1'b0;
      decode_v_r_20_sv2v_reg <= 1'b0;
      decode_v_r_19_sv2v_reg <= 1'b0;
      decode_v_r_18_sv2v_reg <= 1'b0;
      decode_v_r_17_sv2v_reg <= 1'b0;
      decode_v_r_16_sv2v_reg <= 1'b0;
      decode_v_r_15_sv2v_reg <= 1'b0;
      decode_v_r_14_sv2v_reg <= 1'b0;
      decode_v_r_13_sv2v_reg <= 1'b0;
      decode_v_r_12_sv2v_reg <= 1'b0;
      decode_v_r_11_sv2v_reg <= 1'b0;
      decode_v_r_10_sv2v_reg <= 1'b0;
      decode_v_r_9_sv2v_reg <= 1'b0;
      decode_v_r_8_sv2v_reg <= 1'b0;
      decode_v_r_7_sv2v_reg <= 1'b0;
      decode_v_r_6_sv2v_reg <= 1'b0;
      decode_v_r_5_sv2v_reg <= 1'b0;
      decode_v_r_4_sv2v_reg <= 1'b0;
      decode_v_r_3_sv2v_reg <= 1'b0;
      decode_v_r_2_sv2v_reg <= 1'b0;
      decode_v_r_1_sv2v_reg <= 1'b0;
      decode_v_r_0_sv2v_reg <= 1'b0;
      addr_v_r_6_sv2v_reg <= 1'b0;
      addr_v_r_5_sv2v_reg <= 1'b0;
      addr_v_r_4_sv2v_reg <= 1'b0;
      addr_v_r_3_sv2v_reg <= 1'b0;
      addr_v_r_2_sv2v_reg <= 1'b0;
      addr_v_r_1_sv2v_reg <= 1'b0;
      addr_v_r_0_sv2v_reg <= 1'b0;
    end else if(N103) begin
      mask_v_r_15_sv2v_reg <= mask_tl_r[15];
      mask_v_r_14_sv2v_reg <= mask_tl_r[14];
      decode_v_r_20_sv2v_reg <= decode_tl_r[20];
      decode_v_r_19_sv2v_reg <= decode_tl_r[19];
      decode_v_r_18_sv2v_reg <= decode_tl_r[18];
      decode_v_r_17_sv2v_reg <= decode_tl_r[17];
      decode_v_r_16_sv2v_reg <= decode_tl_r[16];
      decode_v_r_15_sv2v_reg <= decode_tl_r[15];
      decode_v_r_14_sv2v_reg <= decode_tl_r[14];
      decode_v_r_13_sv2v_reg <= decode_tl_r[13];
      decode_v_r_12_sv2v_reg <= decode_tl_r[12];
      decode_v_r_11_sv2v_reg <= decode_tl_r[11];
      decode_v_r_10_sv2v_reg <= decode_tl_r[10];
      decode_v_r_9_sv2v_reg <= decode_tl_r[9];
      decode_v_r_8_sv2v_reg <= decode_tl_r[8];
      decode_v_r_7_sv2v_reg <= decode_tl_r[7];
      decode_v_r_6_sv2v_reg <= decode_tl_r[6];
      decode_v_r_5_sv2v_reg <= decode_tl_r[5];
      decode_v_r_4_sv2v_reg <= decode_tl_r[4];
      decode_v_r_3_sv2v_reg <= decode_tl_r[3];
      decode_v_r_2_sv2v_reg <= decode_tl_r[2];
      decode_v_r_1_sv2v_reg <= decode_tl_r[1];
      decode_v_r_0_sv2v_reg <= decode_tl_r[0];
      addr_v_r_6_sv2v_reg <= addr_tl_r[6];
      addr_v_r_5_sv2v_reg <= addr_tl_r[5];
      addr_v_r_4_sv2v_reg <= addr_tl_r[4];
      addr_v_r_3_sv2v_reg <= addr_tl_r[3];
      addr_v_r_2_sv2v_reg <= addr_tl_r[2];
      addr_v_r_1_sv2v_reg <= addr_tl_r[1];
      addr_v_r_0_sv2v_reg <= addr_tl_r[0];
    end 
    if(reset_i) begin
      mask_v_r_13_sv2v_reg <= 1'b0;
      addr_v_r_32_sv2v_reg <= 1'b0;
      addr_v_r_31_sv2v_reg <= 1'b0;
      addr_v_r_30_sv2v_reg <= 1'b0;
      addr_v_r_29_sv2v_reg <= 1'b0;
      addr_v_r_28_sv2v_reg <= 1'b0;
      addr_v_r_27_sv2v_reg <= 1'b0;
      addr_v_r_26_sv2v_reg <= 1'b0;
      addr_v_r_25_sv2v_reg <= 1'b0;
      addr_v_r_24_sv2v_reg <= 1'b0;
      addr_v_r_23_sv2v_reg <= 1'b0;
      addr_v_r_22_sv2v_reg <= 1'b0;
      addr_v_r_21_sv2v_reg <= 1'b0;
      addr_v_r_20_sv2v_reg <= 1'b0;
      addr_v_r_19_sv2v_reg <= 1'b0;
      addr_v_r_18_sv2v_reg <= 1'b0;
      addr_v_r_17_sv2v_reg <= 1'b0;
      addr_v_r_16_sv2v_reg <= 1'b0;
      addr_v_r_15_sv2v_reg <= 1'b0;
      addr_v_r_14_sv2v_reg <= 1'b0;
      addr_v_r_13_sv2v_reg <= 1'b0;
      addr_v_r_12_sv2v_reg <= 1'b0;
      addr_v_r_11_sv2v_reg <= 1'b0;
      addr_v_r_10_sv2v_reg <= 1'b0;
      addr_v_r_9_sv2v_reg <= 1'b0;
      addr_v_r_8_sv2v_reg <= 1'b0;
      addr_v_r_7_sv2v_reg <= 1'b0;
      data_v_r_72_sv2v_reg <= 1'b0;
      data_v_r_71_sv2v_reg <= 1'b0;
      data_v_r_70_sv2v_reg <= 1'b0;
      data_v_r_69_sv2v_reg <= 1'b0;
      data_v_r_68_sv2v_reg <= 1'b0;
      data_v_r_67_sv2v_reg <= 1'b0;
      data_v_r_66_sv2v_reg <= 1'b0;
      data_v_r_65_sv2v_reg <= 1'b0;
      data_v_r_64_sv2v_reg <= 1'b0;
      data_v_r_63_sv2v_reg <= 1'b0;
      data_v_r_62_sv2v_reg <= 1'b0;
      data_v_r_61_sv2v_reg <= 1'b0;
      data_v_r_60_sv2v_reg <= 1'b0;
      data_v_r_59_sv2v_reg <= 1'b0;
      data_v_r_58_sv2v_reg <= 1'b0;
      data_v_r_57_sv2v_reg <= 1'b0;
      data_v_r_56_sv2v_reg <= 1'b0;
      data_v_r_55_sv2v_reg <= 1'b0;
      data_v_r_54_sv2v_reg <= 1'b0;
      data_v_r_53_sv2v_reg <= 1'b0;
      data_v_r_52_sv2v_reg <= 1'b0;
      data_v_r_51_sv2v_reg <= 1'b0;
      data_v_r_50_sv2v_reg <= 1'b0;
      data_v_r_49_sv2v_reg <= 1'b0;
      data_v_r_48_sv2v_reg <= 1'b0;
      data_v_r_47_sv2v_reg <= 1'b0;
      data_v_r_46_sv2v_reg <= 1'b0;
      data_v_r_45_sv2v_reg <= 1'b0;
      data_v_r_44_sv2v_reg <= 1'b0;
      data_v_r_43_sv2v_reg <= 1'b0;
      data_v_r_42_sv2v_reg <= 1'b0;
      data_v_r_41_sv2v_reg <= 1'b0;
      data_v_r_40_sv2v_reg <= 1'b0;
      data_v_r_39_sv2v_reg <= 1'b0;
      data_v_r_38_sv2v_reg <= 1'b0;
      data_v_r_37_sv2v_reg <= 1'b0;
      data_v_r_36_sv2v_reg <= 1'b0;
      data_v_r_35_sv2v_reg <= 1'b0;
      data_v_r_34_sv2v_reg <= 1'b0;
      data_v_r_33_sv2v_reg <= 1'b0;
      data_v_r_32_sv2v_reg <= 1'b0;
      data_v_r_31_sv2v_reg <= 1'b0;
      data_v_r_30_sv2v_reg <= 1'b0;
      data_v_r_29_sv2v_reg <= 1'b0;
      data_v_r_28_sv2v_reg <= 1'b0;
      data_v_r_27_sv2v_reg <= 1'b0;
      data_v_r_26_sv2v_reg <= 1'b0;
      data_v_r_25_sv2v_reg <= 1'b0;
      data_v_r_24_sv2v_reg <= 1'b0;
      data_v_r_23_sv2v_reg <= 1'b0;
      data_v_r_22_sv2v_reg <= 1'b0;
      data_v_r_21_sv2v_reg <= 1'b0;
      data_v_r_20_sv2v_reg <= 1'b0;
      data_v_r_19_sv2v_reg <= 1'b0;
      data_v_r_18_sv2v_reg <= 1'b0;
      data_v_r_17_sv2v_reg <= 1'b0;
      data_v_r_16_sv2v_reg <= 1'b0;
      data_v_r_15_sv2v_reg <= 1'b0;
      data_v_r_14_sv2v_reg <= 1'b0;
      data_v_r_13_sv2v_reg <= 1'b0;
      data_v_r_12_sv2v_reg <= 1'b0;
      data_v_r_11_sv2v_reg <= 1'b0;
      data_v_r_10_sv2v_reg <= 1'b0;
      data_v_r_9_sv2v_reg <= 1'b0;
      data_v_r_8_sv2v_reg <= 1'b0;
      data_v_r_7_sv2v_reg <= 1'b0;
      data_v_r_6_sv2v_reg <= 1'b0;
      data_v_r_5_sv2v_reg <= 1'b0;
      data_v_r_4_sv2v_reg <= 1'b0;
      data_v_r_3_sv2v_reg <= 1'b0;
      data_v_r_2_sv2v_reg <= 1'b0;
      data_v_r_1_sv2v_reg <= 1'b0;
      data_v_r_0_sv2v_reg <= 1'b0;
    end else if(N102) begin
      mask_v_r_13_sv2v_reg <= mask_tl_r[13];
      addr_v_r_32_sv2v_reg <= addr_tl_r[32];
      addr_v_r_31_sv2v_reg <= addr_tl_r[31];
      addr_v_r_30_sv2v_reg <= addr_tl_r[30];
      addr_v_r_29_sv2v_reg <= addr_tl_r[29];
      addr_v_r_28_sv2v_reg <= addr_tl_r[28];
      addr_v_r_27_sv2v_reg <= addr_tl_r[27];
      addr_v_r_26_sv2v_reg <= addr_tl_r[26];
      addr_v_r_25_sv2v_reg <= addr_tl_r[25];
      addr_v_r_24_sv2v_reg <= addr_tl_r[24];
      addr_v_r_23_sv2v_reg <= addr_tl_r[23];
      addr_v_r_22_sv2v_reg <= addr_tl_r[22];
      addr_v_r_21_sv2v_reg <= addr_tl_r[21];
      addr_v_r_20_sv2v_reg <= addr_tl_r[20];
      addr_v_r_19_sv2v_reg <= addr_tl_r[19];
      addr_v_r_18_sv2v_reg <= addr_tl_r[18];
      addr_v_r_17_sv2v_reg <= addr_tl_r[17];
      addr_v_r_16_sv2v_reg <= addr_tl_r[16];
      addr_v_r_15_sv2v_reg <= addr_tl_r[15];
      addr_v_r_14_sv2v_reg <= addr_tl_r[14];
      addr_v_r_13_sv2v_reg <= addr_tl_r[13];
      addr_v_r_12_sv2v_reg <= addr_tl_r[12];
      addr_v_r_11_sv2v_reg <= addr_tl_r[11];
      addr_v_r_10_sv2v_reg <= addr_tl_r[10];
      addr_v_r_9_sv2v_reg <= addr_tl_r[9];
      addr_v_r_8_sv2v_reg <= addr_tl_r[8];
      addr_v_r_7_sv2v_reg <= addr_tl_r[7];
      data_v_r_72_sv2v_reg <= data_tl_r[72];
      data_v_r_71_sv2v_reg <= data_tl_r[71];
      data_v_r_70_sv2v_reg <= data_tl_r[70];
      data_v_r_69_sv2v_reg <= data_tl_r[69];
      data_v_r_68_sv2v_reg <= data_tl_r[68];
      data_v_r_67_sv2v_reg <= data_tl_r[67];
      data_v_r_66_sv2v_reg <= data_tl_r[66];
      data_v_r_65_sv2v_reg <= data_tl_r[65];
      data_v_r_64_sv2v_reg <= data_tl_r[64];
      data_v_r_63_sv2v_reg <= data_tl_r[63];
      data_v_r_62_sv2v_reg <= data_tl_r[62];
      data_v_r_61_sv2v_reg <= data_tl_r[61];
      data_v_r_60_sv2v_reg <= data_tl_r[60];
      data_v_r_59_sv2v_reg <= data_tl_r[59];
      data_v_r_58_sv2v_reg <= data_tl_r[58];
      data_v_r_57_sv2v_reg <= data_tl_r[57];
      data_v_r_56_sv2v_reg <= data_tl_r[56];
      data_v_r_55_sv2v_reg <= data_tl_r[55];
      data_v_r_54_sv2v_reg <= data_tl_r[54];
      data_v_r_53_sv2v_reg <= data_tl_r[53];
      data_v_r_52_sv2v_reg <= data_tl_r[52];
      data_v_r_51_sv2v_reg <= data_tl_r[51];
      data_v_r_50_sv2v_reg <= data_tl_r[50];
      data_v_r_49_sv2v_reg <= data_tl_r[49];
      data_v_r_48_sv2v_reg <= data_tl_r[48];
      data_v_r_47_sv2v_reg <= data_tl_r[47];
      data_v_r_46_sv2v_reg <= data_tl_r[46];
      data_v_r_45_sv2v_reg <= data_tl_r[45];
      data_v_r_44_sv2v_reg <= data_tl_r[44];
      data_v_r_43_sv2v_reg <= data_tl_r[43];
      data_v_r_42_sv2v_reg <= data_tl_r[42];
      data_v_r_41_sv2v_reg <= data_tl_r[41];
      data_v_r_40_sv2v_reg <= data_tl_r[40];
      data_v_r_39_sv2v_reg <= data_tl_r[39];
      data_v_r_38_sv2v_reg <= data_tl_r[38];
      data_v_r_37_sv2v_reg <= data_tl_r[37];
      data_v_r_36_sv2v_reg <= data_tl_r[36];
      data_v_r_35_sv2v_reg <= data_tl_r[35];
      data_v_r_34_sv2v_reg <= data_tl_r[34];
      data_v_r_33_sv2v_reg <= data_tl_r[33];
      data_v_r_32_sv2v_reg <= data_tl_r[32];
      data_v_r_31_sv2v_reg <= data_tl_r[31];
      data_v_r_30_sv2v_reg <= data_tl_r[30];
      data_v_r_29_sv2v_reg <= data_tl_r[29];
      data_v_r_28_sv2v_reg <= data_tl_r[28];
      data_v_r_27_sv2v_reg <= data_tl_r[27];
      data_v_r_26_sv2v_reg <= data_tl_r[26];
      data_v_r_25_sv2v_reg <= data_tl_r[25];
      data_v_r_24_sv2v_reg <= data_tl_r[24];
      data_v_r_23_sv2v_reg <= data_tl_r[23];
      data_v_r_22_sv2v_reg <= data_tl_r[22];
      data_v_r_21_sv2v_reg <= data_tl_r[21];
      data_v_r_20_sv2v_reg <= data_tl_r[20];
      data_v_r_19_sv2v_reg <= data_tl_r[19];
      data_v_r_18_sv2v_reg <= data_tl_r[18];
      data_v_r_17_sv2v_reg <= data_tl_r[17];
      data_v_r_16_sv2v_reg <= data_tl_r[16];
      data_v_r_15_sv2v_reg <= data_tl_r[15];
      data_v_r_14_sv2v_reg <= data_tl_r[14];
      data_v_r_13_sv2v_reg <= data_tl_r[13];
      data_v_r_12_sv2v_reg <= data_tl_r[12];
      data_v_r_11_sv2v_reg <= data_tl_r[11];
      data_v_r_10_sv2v_reg <= data_tl_r[10];
      data_v_r_9_sv2v_reg <= data_tl_r[9];
      data_v_r_8_sv2v_reg <= data_tl_r[8];
      data_v_r_7_sv2v_reg <= data_tl_r[7];
      data_v_r_6_sv2v_reg <= data_tl_r[6];
      data_v_r_5_sv2v_reg <= data_tl_r[5];
      data_v_r_4_sv2v_reg <= data_tl_r[4];
      data_v_r_3_sv2v_reg <= data_tl_r[3];
      data_v_r_2_sv2v_reg <= data_tl_r[2];
      data_v_r_1_sv2v_reg <= data_tl_r[1];
      data_v_r_0_sv2v_reg <= data_tl_r[0];
    end 
    if(reset_i) begin
      mask_v_r_12_sv2v_reg <= 1'b0;
      data_v_r_127_sv2v_reg <= 1'b0;
      data_v_r_126_sv2v_reg <= 1'b0;
      data_v_r_125_sv2v_reg <= 1'b0;
      data_v_r_124_sv2v_reg <= 1'b0;
      data_v_r_123_sv2v_reg <= 1'b0;
      data_v_r_122_sv2v_reg <= 1'b0;
      data_v_r_121_sv2v_reg <= 1'b0;
      data_v_r_120_sv2v_reg <= 1'b0;
      data_v_r_119_sv2v_reg <= 1'b0;
      data_v_r_118_sv2v_reg <= 1'b0;
      data_v_r_117_sv2v_reg <= 1'b0;
      data_v_r_116_sv2v_reg <= 1'b0;
      data_v_r_115_sv2v_reg <= 1'b0;
      data_v_r_114_sv2v_reg <= 1'b0;
      data_v_r_113_sv2v_reg <= 1'b0;
      data_v_r_112_sv2v_reg <= 1'b0;
      data_v_r_111_sv2v_reg <= 1'b0;
      data_v_r_110_sv2v_reg <= 1'b0;
      data_v_r_109_sv2v_reg <= 1'b0;
      data_v_r_108_sv2v_reg <= 1'b0;
      data_v_r_107_sv2v_reg <= 1'b0;
      data_v_r_106_sv2v_reg <= 1'b0;
      data_v_r_105_sv2v_reg <= 1'b0;
      data_v_r_104_sv2v_reg <= 1'b0;
      data_v_r_103_sv2v_reg <= 1'b0;
      data_v_r_102_sv2v_reg <= 1'b0;
      data_v_r_101_sv2v_reg <= 1'b0;
      data_v_r_100_sv2v_reg <= 1'b0;
      data_v_r_99_sv2v_reg <= 1'b0;
      data_v_r_98_sv2v_reg <= 1'b0;
      data_v_r_97_sv2v_reg <= 1'b0;
      data_v_r_96_sv2v_reg <= 1'b0;
      data_v_r_95_sv2v_reg <= 1'b0;
      data_v_r_94_sv2v_reg <= 1'b0;
      data_v_r_93_sv2v_reg <= 1'b0;
      data_v_r_92_sv2v_reg <= 1'b0;
      data_v_r_91_sv2v_reg <= 1'b0;
      data_v_r_90_sv2v_reg <= 1'b0;
      data_v_r_89_sv2v_reg <= 1'b0;
      data_v_r_88_sv2v_reg <= 1'b0;
      data_v_r_87_sv2v_reg <= 1'b0;
      data_v_r_86_sv2v_reg <= 1'b0;
      data_v_r_85_sv2v_reg <= 1'b0;
      data_v_r_84_sv2v_reg <= 1'b0;
      data_v_r_83_sv2v_reg <= 1'b0;
      data_v_r_82_sv2v_reg <= 1'b0;
      data_v_r_81_sv2v_reg <= 1'b0;
      data_v_r_80_sv2v_reg <= 1'b0;
      data_v_r_79_sv2v_reg <= 1'b0;
      data_v_r_78_sv2v_reg <= 1'b0;
      data_v_r_77_sv2v_reg <= 1'b0;
      data_v_r_76_sv2v_reg <= 1'b0;
      data_v_r_75_sv2v_reg <= 1'b0;
      data_v_r_74_sv2v_reg <= 1'b0;
      data_v_r_73_sv2v_reg <= 1'b0;
      valid_v_r_7_sv2v_reg <= 1'b0;
      valid_v_r_6_sv2v_reg <= 1'b0;
      valid_v_r_5_sv2v_reg <= 1'b0;
      valid_v_r_4_sv2v_reg <= 1'b0;
      valid_v_r_3_sv2v_reg <= 1'b0;
      valid_v_r_2_sv2v_reg <= 1'b0;
      valid_v_r_1_sv2v_reg <= 1'b0;
      valid_v_r_0_sv2v_reg <= 1'b0;
      tag_v_r_35_sv2v_reg <= 1'b0;
      tag_v_r_34_sv2v_reg <= 1'b0;
      tag_v_r_33_sv2v_reg <= 1'b0;
      tag_v_r_32_sv2v_reg <= 1'b0;
      tag_v_r_31_sv2v_reg <= 1'b0;
      tag_v_r_30_sv2v_reg <= 1'b0;
      tag_v_r_29_sv2v_reg <= 1'b0;
      tag_v_r_28_sv2v_reg <= 1'b0;
      tag_v_r_27_sv2v_reg <= 1'b0;
      tag_v_r_26_sv2v_reg <= 1'b0;
      tag_v_r_25_sv2v_reg <= 1'b0;
      tag_v_r_24_sv2v_reg <= 1'b0;
      tag_v_r_23_sv2v_reg <= 1'b0;
      tag_v_r_22_sv2v_reg <= 1'b0;
      tag_v_r_21_sv2v_reg <= 1'b0;
      tag_v_r_20_sv2v_reg <= 1'b0;
      tag_v_r_19_sv2v_reg <= 1'b0;
      tag_v_r_18_sv2v_reg <= 1'b0;
      tag_v_r_17_sv2v_reg <= 1'b0;
      tag_v_r_16_sv2v_reg <= 1'b0;
      tag_v_r_15_sv2v_reg <= 1'b0;
      tag_v_r_14_sv2v_reg <= 1'b0;
      tag_v_r_13_sv2v_reg <= 1'b0;
      tag_v_r_12_sv2v_reg <= 1'b0;
      tag_v_r_11_sv2v_reg <= 1'b0;
      tag_v_r_10_sv2v_reg <= 1'b0;
      tag_v_r_9_sv2v_reg <= 1'b0;
      tag_v_r_8_sv2v_reg <= 1'b0;
      tag_v_r_7_sv2v_reg <= 1'b0;
      tag_v_r_6_sv2v_reg <= 1'b0;
      tag_v_r_5_sv2v_reg <= 1'b0;
      tag_v_r_4_sv2v_reg <= 1'b0;
      tag_v_r_3_sv2v_reg <= 1'b0;
      tag_v_r_2_sv2v_reg <= 1'b0;
      tag_v_r_1_sv2v_reg <= 1'b0;
      tag_v_r_0_sv2v_reg <= 1'b0;
    end else if(N101) begin
      mask_v_r_12_sv2v_reg <= mask_tl_r[12];
      data_v_r_127_sv2v_reg <= data_tl_r[127];
      data_v_r_126_sv2v_reg <= data_tl_r[126];
      data_v_r_125_sv2v_reg <= data_tl_r[125];
      data_v_r_124_sv2v_reg <= data_tl_r[124];
      data_v_r_123_sv2v_reg <= data_tl_r[123];
      data_v_r_122_sv2v_reg <= data_tl_r[122];
      data_v_r_121_sv2v_reg <= data_tl_r[121];
      data_v_r_120_sv2v_reg <= data_tl_r[120];
      data_v_r_119_sv2v_reg <= data_tl_r[119];
      data_v_r_118_sv2v_reg <= data_tl_r[118];
      data_v_r_117_sv2v_reg <= data_tl_r[117];
      data_v_r_116_sv2v_reg <= data_tl_r[116];
      data_v_r_115_sv2v_reg <= data_tl_r[115];
      data_v_r_114_sv2v_reg <= data_tl_r[114];
      data_v_r_113_sv2v_reg <= data_tl_r[113];
      data_v_r_112_sv2v_reg <= data_tl_r[112];
      data_v_r_111_sv2v_reg <= data_tl_r[111];
      data_v_r_110_sv2v_reg <= data_tl_r[110];
      data_v_r_109_sv2v_reg <= data_tl_r[109];
      data_v_r_108_sv2v_reg <= data_tl_r[108];
      data_v_r_107_sv2v_reg <= data_tl_r[107];
      data_v_r_106_sv2v_reg <= data_tl_r[106];
      data_v_r_105_sv2v_reg <= data_tl_r[105];
      data_v_r_104_sv2v_reg <= data_tl_r[104];
      data_v_r_103_sv2v_reg <= data_tl_r[103];
      data_v_r_102_sv2v_reg <= data_tl_r[102];
      data_v_r_101_sv2v_reg <= data_tl_r[101];
      data_v_r_100_sv2v_reg <= data_tl_r[100];
      data_v_r_99_sv2v_reg <= data_tl_r[99];
      data_v_r_98_sv2v_reg <= data_tl_r[98];
      data_v_r_97_sv2v_reg <= data_tl_r[97];
      data_v_r_96_sv2v_reg <= data_tl_r[96];
      data_v_r_95_sv2v_reg <= data_tl_r[95];
      data_v_r_94_sv2v_reg <= data_tl_r[94];
      data_v_r_93_sv2v_reg <= data_tl_r[93];
      data_v_r_92_sv2v_reg <= data_tl_r[92];
      data_v_r_91_sv2v_reg <= data_tl_r[91];
      data_v_r_90_sv2v_reg <= data_tl_r[90];
      data_v_r_89_sv2v_reg <= data_tl_r[89];
      data_v_r_88_sv2v_reg <= data_tl_r[88];
      data_v_r_87_sv2v_reg <= data_tl_r[87];
      data_v_r_86_sv2v_reg <= data_tl_r[86];
      data_v_r_85_sv2v_reg <= data_tl_r[85];
      data_v_r_84_sv2v_reg <= data_tl_r[84];
      data_v_r_83_sv2v_reg <= data_tl_r[83];
      data_v_r_82_sv2v_reg <= data_tl_r[82];
      data_v_r_81_sv2v_reg <= data_tl_r[81];
      data_v_r_80_sv2v_reg <= data_tl_r[80];
      data_v_r_79_sv2v_reg <= data_tl_r[79];
      data_v_r_78_sv2v_reg <= data_tl_r[78];
      data_v_r_77_sv2v_reg <= data_tl_r[77];
      data_v_r_76_sv2v_reg <= data_tl_r[76];
      data_v_r_75_sv2v_reg <= data_tl_r[75];
      data_v_r_74_sv2v_reg <= data_tl_r[74];
      data_v_r_73_sv2v_reg <= data_tl_r[73];
      valid_v_r_7_sv2v_reg <= tag_mem_data_lo[175];
      valid_v_r_6_sv2v_reg <= tag_mem_data_lo[153];
      valid_v_r_5_sv2v_reg <= tag_mem_data_lo[131];
      valid_v_r_4_sv2v_reg <= tag_mem_data_lo[109];
      valid_v_r_3_sv2v_reg <= tag_mem_data_lo[87];
      valid_v_r_2_sv2v_reg <= tag_mem_data_lo[65];
      valid_v_r_1_sv2v_reg <= tag_mem_data_lo[43];
      valid_v_r_0_sv2v_reg <= tag_mem_data_lo[21];
      tag_v_r_35_sv2v_reg <= tag_mem_data_lo[37];
      tag_v_r_34_sv2v_reg <= tag_mem_data_lo[36];
      tag_v_r_33_sv2v_reg <= tag_mem_data_lo[35];
      tag_v_r_32_sv2v_reg <= tag_mem_data_lo[34];
      tag_v_r_31_sv2v_reg <= tag_mem_data_lo[33];
      tag_v_r_30_sv2v_reg <= tag_mem_data_lo[32];
      tag_v_r_29_sv2v_reg <= tag_mem_data_lo[31];
      tag_v_r_28_sv2v_reg <= tag_mem_data_lo[30];
      tag_v_r_27_sv2v_reg <= tag_mem_data_lo[29];
      tag_v_r_26_sv2v_reg <= tag_mem_data_lo[28];
      tag_v_r_25_sv2v_reg <= tag_mem_data_lo[27];
      tag_v_r_24_sv2v_reg <= tag_mem_data_lo[26];
      tag_v_r_23_sv2v_reg <= tag_mem_data_lo[25];
      tag_v_r_22_sv2v_reg <= tag_mem_data_lo[24];
      tag_v_r_21_sv2v_reg <= tag_mem_data_lo[23];
      tag_v_r_20_sv2v_reg <= tag_mem_data_lo[22];
      tag_v_r_19_sv2v_reg <= tag_mem_data_lo[19];
      tag_v_r_18_sv2v_reg <= tag_mem_data_lo[18];
      tag_v_r_17_sv2v_reg <= tag_mem_data_lo[17];
      tag_v_r_16_sv2v_reg <= tag_mem_data_lo[16];
      tag_v_r_15_sv2v_reg <= tag_mem_data_lo[15];
      tag_v_r_14_sv2v_reg <= tag_mem_data_lo[14];
      tag_v_r_13_sv2v_reg <= tag_mem_data_lo[13];
      tag_v_r_12_sv2v_reg <= tag_mem_data_lo[12];
      tag_v_r_11_sv2v_reg <= tag_mem_data_lo[11];
      tag_v_r_10_sv2v_reg <= tag_mem_data_lo[10];
      tag_v_r_9_sv2v_reg <= tag_mem_data_lo[9];
      tag_v_r_8_sv2v_reg <= tag_mem_data_lo[8];
      tag_v_r_7_sv2v_reg <= tag_mem_data_lo[7];
      tag_v_r_6_sv2v_reg <= tag_mem_data_lo[6];
      tag_v_r_5_sv2v_reg <= tag_mem_data_lo[5];
      tag_v_r_4_sv2v_reg <= tag_mem_data_lo[4];
      tag_v_r_3_sv2v_reg <= tag_mem_data_lo[3];
      tag_v_r_2_sv2v_reg <= tag_mem_data_lo[2];
      tag_v_r_1_sv2v_reg <= tag_mem_data_lo[1];
      tag_v_r_0_sv2v_reg <= tag_mem_data_lo[0];
    end 
    if(reset_i) begin
      mask_v_r_11_sv2v_reg <= 1'b0;
      tag_v_r_134_sv2v_reg <= 1'b0;
      tag_v_r_133_sv2v_reg <= 1'b0;
      tag_v_r_132_sv2v_reg <= 1'b0;
      tag_v_r_131_sv2v_reg <= 1'b0;
      tag_v_r_130_sv2v_reg <= 1'b0;
      tag_v_r_129_sv2v_reg <= 1'b0;
      tag_v_r_128_sv2v_reg <= 1'b0;
      tag_v_r_127_sv2v_reg <= 1'b0;
      tag_v_r_126_sv2v_reg <= 1'b0;
      tag_v_r_125_sv2v_reg <= 1'b0;
      tag_v_r_124_sv2v_reg <= 1'b0;
      tag_v_r_123_sv2v_reg <= 1'b0;
      tag_v_r_122_sv2v_reg <= 1'b0;
      tag_v_r_121_sv2v_reg <= 1'b0;
      tag_v_r_120_sv2v_reg <= 1'b0;
      tag_v_r_119_sv2v_reg <= 1'b0;
      tag_v_r_118_sv2v_reg <= 1'b0;
      tag_v_r_117_sv2v_reg <= 1'b0;
      tag_v_r_116_sv2v_reg <= 1'b0;
      tag_v_r_115_sv2v_reg <= 1'b0;
      tag_v_r_114_sv2v_reg <= 1'b0;
      tag_v_r_113_sv2v_reg <= 1'b0;
      tag_v_r_112_sv2v_reg <= 1'b0;
      tag_v_r_111_sv2v_reg <= 1'b0;
      tag_v_r_110_sv2v_reg <= 1'b0;
      tag_v_r_109_sv2v_reg <= 1'b0;
      tag_v_r_108_sv2v_reg <= 1'b0;
      tag_v_r_107_sv2v_reg <= 1'b0;
      tag_v_r_106_sv2v_reg <= 1'b0;
      tag_v_r_105_sv2v_reg <= 1'b0;
      tag_v_r_104_sv2v_reg <= 1'b0;
      tag_v_r_103_sv2v_reg <= 1'b0;
      tag_v_r_102_sv2v_reg <= 1'b0;
      tag_v_r_101_sv2v_reg <= 1'b0;
      tag_v_r_100_sv2v_reg <= 1'b0;
      tag_v_r_99_sv2v_reg <= 1'b0;
      tag_v_r_98_sv2v_reg <= 1'b0;
      tag_v_r_97_sv2v_reg <= 1'b0;
      tag_v_r_96_sv2v_reg <= 1'b0;
      tag_v_r_95_sv2v_reg <= 1'b0;
      tag_v_r_94_sv2v_reg <= 1'b0;
      tag_v_r_93_sv2v_reg <= 1'b0;
      tag_v_r_92_sv2v_reg <= 1'b0;
      tag_v_r_91_sv2v_reg <= 1'b0;
      tag_v_r_90_sv2v_reg <= 1'b0;
      tag_v_r_89_sv2v_reg <= 1'b0;
      tag_v_r_88_sv2v_reg <= 1'b0;
      tag_v_r_87_sv2v_reg <= 1'b0;
      tag_v_r_86_sv2v_reg <= 1'b0;
      tag_v_r_85_sv2v_reg <= 1'b0;
      tag_v_r_84_sv2v_reg <= 1'b0;
      tag_v_r_83_sv2v_reg <= 1'b0;
      tag_v_r_82_sv2v_reg <= 1'b0;
      tag_v_r_81_sv2v_reg <= 1'b0;
      tag_v_r_80_sv2v_reg <= 1'b0;
      tag_v_r_79_sv2v_reg <= 1'b0;
      tag_v_r_78_sv2v_reg <= 1'b0;
      tag_v_r_77_sv2v_reg <= 1'b0;
      tag_v_r_76_sv2v_reg <= 1'b0;
      tag_v_r_75_sv2v_reg <= 1'b0;
      tag_v_r_74_sv2v_reg <= 1'b0;
      tag_v_r_73_sv2v_reg <= 1'b0;
      tag_v_r_72_sv2v_reg <= 1'b0;
      tag_v_r_71_sv2v_reg <= 1'b0;
      tag_v_r_70_sv2v_reg <= 1'b0;
      tag_v_r_69_sv2v_reg <= 1'b0;
      tag_v_r_68_sv2v_reg <= 1'b0;
      tag_v_r_67_sv2v_reg <= 1'b0;
      tag_v_r_66_sv2v_reg <= 1'b0;
      tag_v_r_65_sv2v_reg <= 1'b0;
      tag_v_r_64_sv2v_reg <= 1'b0;
      tag_v_r_63_sv2v_reg <= 1'b0;
      tag_v_r_62_sv2v_reg <= 1'b0;
      tag_v_r_61_sv2v_reg <= 1'b0;
      tag_v_r_60_sv2v_reg <= 1'b0;
      tag_v_r_59_sv2v_reg <= 1'b0;
      tag_v_r_58_sv2v_reg <= 1'b0;
      tag_v_r_57_sv2v_reg <= 1'b0;
      tag_v_r_56_sv2v_reg <= 1'b0;
      tag_v_r_55_sv2v_reg <= 1'b0;
      tag_v_r_54_sv2v_reg <= 1'b0;
      tag_v_r_53_sv2v_reg <= 1'b0;
      tag_v_r_52_sv2v_reg <= 1'b0;
      tag_v_r_51_sv2v_reg <= 1'b0;
      tag_v_r_50_sv2v_reg <= 1'b0;
      tag_v_r_49_sv2v_reg <= 1'b0;
      tag_v_r_48_sv2v_reg <= 1'b0;
      tag_v_r_47_sv2v_reg <= 1'b0;
      tag_v_r_46_sv2v_reg <= 1'b0;
      tag_v_r_45_sv2v_reg <= 1'b0;
      tag_v_r_44_sv2v_reg <= 1'b0;
      tag_v_r_43_sv2v_reg <= 1'b0;
      tag_v_r_42_sv2v_reg <= 1'b0;
      tag_v_r_41_sv2v_reg <= 1'b0;
      tag_v_r_40_sv2v_reg <= 1'b0;
      tag_v_r_39_sv2v_reg <= 1'b0;
      tag_v_r_38_sv2v_reg <= 1'b0;
      tag_v_r_37_sv2v_reg <= 1'b0;
      tag_v_r_36_sv2v_reg <= 1'b0;
    end else if(N100) begin
      mask_v_r_11_sv2v_reg <= mask_tl_r[11];
      tag_v_r_134_sv2v_reg <= tag_mem_data_lo[146];
      tag_v_r_133_sv2v_reg <= tag_mem_data_lo[145];
      tag_v_r_132_sv2v_reg <= tag_mem_data_lo[144];
      tag_v_r_131_sv2v_reg <= tag_mem_data_lo[143];
      tag_v_r_130_sv2v_reg <= tag_mem_data_lo[142];
      tag_v_r_129_sv2v_reg <= tag_mem_data_lo[141];
      tag_v_r_128_sv2v_reg <= tag_mem_data_lo[140];
      tag_v_r_127_sv2v_reg <= tag_mem_data_lo[139];
      tag_v_r_126_sv2v_reg <= tag_mem_data_lo[138];
      tag_v_r_125_sv2v_reg <= tag_mem_data_lo[137];
      tag_v_r_124_sv2v_reg <= tag_mem_data_lo[136];
      tag_v_r_123_sv2v_reg <= tag_mem_data_lo[135];
      tag_v_r_122_sv2v_reg <= tag_mem_data_lo[134];
      tag_v_r_121_sv2v_reg <= tag_mem_data_lo[133];
      tag_v_r_120_sv2v_reg <= tag_mem_data_lo[132];
      tag_v_r_119_sv2v_reg <= tag_mem_data_lo[129];
      tag_v_r_118_sv2v_reg <= tag_mem_data_lo[128];
      tag_v_r_117_sv2v_reg <= tag_mem_data_lo[127];
      tag_v_r_116_sv2v_reg <= tag_mem_data_lo[126];
      tag_v_r_115_sv2v_reg <= tag_mem_data_lo[125];
      tag_v_r_114_sv2v_reg <= tag_mem_data_lo[124];
      tag_v_r_113_sv2v_reg <= tag_mem_data_lo[123];
      tag_v_r_112_sv2v_reg <= tag_mem_data_lo[122];
      tag_v_r_111_sv2v_reg <= tag_mem_data_lo[121];
      tag_v_r_110_sv2v_reg <= tag_mem_data_lo[120];
      tag_v_r_109_sv2v_reg <= tag_mem_data_lo[119];
      tag_v_r_108_sv2v_reg <= tag_mem_data_lo[118];
      tag_v_r_107_sv2v_reg <= tag_mem_data_lo[117];
      tag_v_r_106_sv2v_reg <= tag_mem_data_lo[116];
      tag_v_r_105_sv2v_reg <= tag_mem_data_lo[115];
      tag_v_r_104_sv2v_reg <= tag_mem_data_lo[114];
      tag_v_r_103_sv2v_reg <= tag_mem_data_lo[113];
      tag_v_r_102_sv2v_reg <= tag_mem_data_lo[112];
      tag_v_r_101_sv2v_reg <= tag_mem_data_lo[111];
      tag_v_r_100_sv2v_reg <= tag_mem_data_lo[110];
      tag_v_r_99_sv2v_reg <= tag_mem_data_lo[107];
      tag_v_r_98_sv2v_reg <= tag_mem_data_lo[106];
      tag_v_r_97_sv2v_reg <= tag_mem_data_lo[105];
      tag_v_r_96_sv2v_reg <= tag_mem_data_lo[104];
      tag_v_r_95_sv2v_reg <= tag_mem_data_lo[103];
      tag_v_r_94_sv2v_reg <= tag_mem_data_lo[102];
      tag_v_r_93_sv2v_reg <= tag_mem_data_lo[101];
      tag_v_r_92_sv2v_reg <= tag_mem_data_lo[100];
      tag_v_r_91_sv2v_reg <= tag_mem_data_lo[99];
      tag_v_r_90_sv2v_reg <= tag_mem_data_lo[98];
      tag_v_r_89_sv2v_reg <= tag_mem_data_lo[97];
      tag_v_r_88_sv2v_reg <= tag_mem_data_lo[96];
      tag_v_r_87_sv2v_reg <= tag_mem_data_lo[95];
      tag_v_r_86_sv2v_reg <= tag_mem_data_lo[94];
      tag_v_r_85_sv2v_reg <= tag_mem_data_lo[93];
      tag_v_r_84_sv2v_reg <= tag_mem_data_lo[92];
      tag_v_r_83_sv2v_reg <= tag_mem_data_lo[91];
      tag_v_r_82_sv2v_reg <= tag_mem_data_lo[90];
      tag_v_r_81_sv2v_reg <= tag_mem_data_lo[89];
      tag_v_r_80_sv2v_reg <= tag_mem_data_lo[88];
      tag_v_r_79_sv2v_reg <= tag_mem_data_lo[85];
      tag_v_r_78_sv2v_reg <= tag_mem_data_lo[84];
      tag_v_r_77_sv2v_reg <= tag_mem_data_lo[83];
      tag_v_r_76_sv2v_reg <= tag_mem_data_lo[82];
      tag_v_r_75_sv2v_reg <= tag_mem_data_lo[81];
      tag_v_r_74_sv2v_reg <= tag_mem_data_lo[80];
      tag_v_r_73_sv2v_reg <= tag_mem_data_lo[79];
      tag_v_r_72_sv2v_reg <= tag_mem_data_lo[78];
      tag_v_r_71_sv2v_reg <= tag_mem_data_lo[77];
      tag_v_r_70_sv2v_reg <= tag_mem_data_lo[76];
      tag_v_r_69_sv2v_reg <= tag_mem_data_lo[75];
      tag_v_r_68_sv2v_reg <= tag_mem_data_lo[74];
      tag_v_r_67_sv2v_reg <= tag_mem_data_lo[73];
      tag_v_r_66_sv2v_reg <= tag_mem_data_lo[72];
      tag_v_r_65_sv2v_reg <= tag_mem_data_lo[71];
      tag_v_r_64_sv2v_reg <= tag_mem_data_lo[70];
      tag_v_r_63_sv2v_reg <= tag_mem_data_lo[69];
      tag_v_r_62_sv2v_reg <= tag_mem_data_lo[68];
      tag_v_r_61_sv2v_reg <= tag_mem_data_lo[67];
      tag_v_r_60_sv2v_reg <= tag_mem_data_lo[66];
      tag_v_r_59_sv2v_reg <= tag_mem_data_lo[63];
      tag_v_r_58_sv2v_reg <= tag_mem_data_lo[62];
      tag_v_r_57_sv2v_reg <= tag_mem_data_lo[61];
      tag_v_r_56_sv2v_reg <= tag_mem_data_lo[60];
      tag_v_r_55_sv2v_reg <= tag_mem_data_lo[59];
      tag_v_r_54_sv2v_reg <= tag_mem_data_lo[58];
      tag_v_r_53_sv2v_reg <= tag_mem_data_lo[57];
      tag_v_r_52_sv2v_reg <= tag_mem_data_lo[56];
      tag_v_r_51_sv2v_reg <= tag_mem_data_lo[55];
      tag_v_r_50_sv2v_reg <= tag_mem_data_lo[54];
      tag_v_r_49_sv2v_reg <= tag_mem_data_lo[53];
      tag_v_r_48_sv2v_reg <= tag_mem_data_lo[52];
      tag_v_r_47_sv2v_reg <= tag_mem_data_lo[51];
      tag_v_r_46_sv2v_reg <= tag_mem_data_lo[50];
      tag_v_r_45_sv2v_reg <= tag_mem_data_lo[49];
      tag_v_r_44_sv2v_reg <= tag_mem_data_lo[48];
      tag_v_r_43_sv2v_reg <= tag_mem_data_lo[47];
      tag_v_r_42_sv2v_reg <= tag_mem_data_lo[46];
      tag_v_r_41_sv2v_reg <= tag_mem_data_lo[45];
      tag_v_r_40_sv2v_reg <= tag_mem_data_lo[44];
      tag_v_r_39_sv2v_reg <= tag_mem_data_lo[41];
      tag_v_r_38_sv2v_reg <= tag_mem_data_lo[40];
      tag_v_r_37_sv2v_reg <= tag_mem_data_lo[39];
      tag_v_r_36_sv2v_reg <= tag_mem_data_lo[38];
    end 
    if(reset_i) begin
      mask_v_r_10_sv2v_reg <= 1'b0;
      lock_v_r_7_sv2v_reg <= 1'b0;
      lock_v_r_6_sv2v_reg <= 1'b0;
      lock_v_r_5_sv2v_reg <= 1'b0;
      lock_v_r_4_sv2v_reg <= 1'b0;
      lock_v_r_3_sv2v_reg <= 1'b0;
      lock_v_r_2_sv2v_reg <= 1'b0;
      lock_v_r_1_sv2v_reg <= 1'b0;
      lock_v_r_0_sv2v_reg <= 1'b0;
      tag_v_r_159_sv2v_reg <= 1'b0;
      tag_v_r_158_sv2v_reg <= 1'b0;
      tag_v_r_157_sv2v_reg <= 1'b0;
      tag_v_r_156_sv2v_reg <= 1'b0;
      tag_v_r_155_sv2v_reg <= 1'b0;
      tag_v_r_154_sv2v_reg <= 1'b0;
      tag_v_r_153_sv2v_reg <= 1'b0;
      tag_v_r_152_sv2v_reg <= 1'b0;
      tag_v_r_151_sv2v_reg <= 1'b0;
      tag_v_r_150_sv2v_reg <= 1'b0;
      tag_v_r_149_sv2v_reg <= 1'b0;
      tag_v_r_148_sv2v_reg <= 1'b0;
      tag_v_r_147_sv2v_reg <= 1'b0;
      tag_v_r_146_sv2v_reg <= 1'b0;
      tag_v_r_145_sv2v_reg <= 1'b0;
      tag_v_r_144_sv2v_reg <= 1'b0;
      tag_v_r_143_sv2v_reg <= 1'b0;
      tag_v_r_142_sv2v_reg <= 1'b0;
      tag_v_r_141_sv2v_reg <= 1'b0;
      tag_v_r_140_sv2v_reg <= 1'b0;
      tag_v_r_139_sv2v_reg <= 1'b0;
      tag_v_r_138_sv2v_reg <= 1'b0;
      tag_v_r_137_sv2v_reg <= 1'b0;
      tag_v_r_136_sv2v_reg <= 1'b0;
      tag_v_r_135_sv2v_reg <= 1'b0;
    end else if(N99) begin
      mask_v_r_10_sv2v_reg <= mask_tl_r[10];
      lock_v_r_7_sv2v_reg <= tag_mem_data_lo[174];
      lock_v_r_6_sv2v_reg <= tag_mem_data_lo[152];
      lock_v_r_5_sv2v_reg <= tag_mem_data_lo[130];
      lock_v_r_4_sv2v_reg <= tag_mem_data_lo[108];
      lock_v_r_3_sv2v_reg <= tag_mem_data_lo[86];
      lock_v_r_2_sv2v_reg <= tag_mem_data_lo[64];
      lock_v_r_1_sv2v_reg <= tag_mem_data_lo[42];
      lock_v_r_0_sv2v_reg <= tag_mem_data_lo[20];
      tag_v_r_159_sv2v_reg <= tag_mem_data_lo[173];
      tag_v_r_158_sv2v_reg <= tag_mem_data_lo[172];
      tag_v_r_157_sv2v_reg <= tag_mem_data_lo[171];
      tag_v_r_156_sv2v_reg <= tag_mem_data_lo[170];
      tag_v_r_155_sv2v_reg <= tag_mem_data_lo[169];
      tag_v_r_154_sv2v_reg <= tag_mem_data_lo[168];
      tag_v_r_153_sv2v_reg <= tag_mem_data_lo[167];
      tag_v_r_152_sv2v_reg <= tag_mem_data_lo[166];
      tag_v_r_151_sv2v_reg <= tag_mem_data_lo[165];
      tag_v_r_150_sv2v_reg <= tag_mem_data_lo[164];
      tag_v_r_149_sv2v_reg <= tag_mem_data_lo[163];
      tag_v_r_148_sv2v_reg <= tag_mem_data_lo[162];
      tag_v_r_147_sv2v_reg <= tag_mem_data_lo[161];
      tag_v_r_146_sv2v_reg <= tag_mem_data_lo[160];
      tag_v_r_145_sv2v_reg <= tag_mem_data_lo[159];
      tag_v_r_144_sv2v_reg <= tag_mem_data_lo[158];
      tag_v_r_143_sv2v_reg <= tag_mem_data_lo[157];
      tag_v_r_142_sv2v_reg <= tag_mem_data_lo[156];
      tag_v_r_141_sv2v_reg <= tag_mem_data_lo[155];
      tag_v_r_140_sv2v_reg <= tag_mem_data_lo[154];
      tag_v_r_139_sv2v_reg <= tag_mem_data_lo[151];
      tag_v_r_138_sv2v_reg <= tag_mem_data_lo[150];
      tag_v_r_137_sv2v_reg <= tag_mem_data_lo[149];
      tag_v_r_136_sv2v_reg <= tag_mem_data_lo[148];
      tag_v_r_135_sv2v_reg <= tag_mem_data_lo[147];
    end 
    if(reset_i) begin
      mask_v_r_9_sv2v_reg <= 1'b0;
    end else if(N98) begin
      mask_v_r_9_sv2v_reg <= mask_tl_r[9];
    end 
    if(reset_i) begin
      mask_v_r_8_sv2v_reg <= 1'b0;
    end else if(N97) begin
      mask_v_r_8_sv2v_reg <= mask_tl_r[8];
    end 
    if(reset_i) begin
      mask_v_r_7_sv2v_reg <= 1'b0;
    end else if(N96) begin
      mask_v_r_7_sv2v_reg <= mask_tl_r[7];
    end 
    if(reset_i) begin
      mask_v_r_6_sv2v_reg <= 1'b0;
    end else if(N95) begin
      mask_v_r_6_sv2v_reg <= mask_tl_r[6];
    end 
    if(reset_i) begin
      mask_v_r_5_sv2v_reg <= 1'b0;
    end else if(N94) begin
      mask_v_r_5_sv2v_reg <= mask_tl_r[5];
    end 
    if(reset_i) begin
      mask_v_r_4_sv2v_reg <= 1'b0;
    end else if(N93) begin
      mask_v_r_4_sv2v_reg <= mask_tl_r[4];
    end 
    if(reset_i) begin
      mask_v_r_3_sv2v_reg <= 1'b0;
    end else if(N92) begin
      mask_v_r_3_sv2v_reg <= mask_tl_r[3];
    end 
    if(reset_i) begin
      mask_v_r_2_sv2v_reg <= 1'b0;
    end else if(N91) begin
      mask_v_r_2_sv2v_reg <= mask_tl_r[2];
    end 
    if(reset_i) begin
      mask_v_r_1_sv2v_reg <= 1'b0;
    end else if(N90) begin
      mask_v_r_1_sv2v_reg <= mask_tl_r[1];
    end 
  end


endmodule



module bp_me_dram_hash_decode_00
(
  daddr_i,
  daddr_o
);

  input [32:0] daddr_i;
  output [32:0] daddr_o;
  wire [32:0] daddr_o;
  assign daddr_o[32] = daddr_i[32];
  assign daddr_o[31] = daddr_i[31];
  assign daddr_o[30] = daddr_i[30];
  assign daddr_o[29] = daddr_i[29];
  assign daddr_o[28] = daddr_i[28];
  assign daddr_o[27] = daddr_i[27];
  assign daddr_o[26] = daddr_i[26];
  assign daddr_o[25] = daddr_i[25];
  assign daddr_o[24] = daddr_i[24];
  assign daddr_o[23] = daddr_i[23];
  assign daddr_o[22] = daddr_i[22];
  assign daddr_o[21] = daddr_i[21];
  assign daddr_o[20] = daddr_i[20];
  assign daddr_o[19] = daddr_i[19];
  assign daddr_o[18] = daddr_i[18];
  assign daddr_o[17] = daddr_i[17];
  assign daddr_o[16] = daddr_i[16];
  assign daddr_o[15] = daddr_i[15];
  assign daddr_o[14] = daddr_i[14];
  assign daddr_o[13] = daddr_i[13];
  assign daddr_o[12] = daddr_i[12];
  assign daddr_o[11] = daddr_i[11];
  assign daddr_o[10] = daddr_i[10];
  assign daddr_o[9] = daddr_i[9];
  assign daddr_o[8] = daddr_i[8];
  assign daddr_o[7] = daddr_i[7];
  assign daddr_o[6] = daddr_i[6];
  assign daddr_o[5] = daddr_i[5];
  assign daddr_o[4] = daddr_i[4];
  assign daddr_o[3] = daddr_i[3];
  assign daddr_o[2] = daddr_i[2];
  assign daddr_o[1] = daddr_i[1];
  assign daddr_o[0] = daddr_i[0];

endmodule



module bp_me_cache_slice
(
  clk_i,
  reset_i,
  mem_fwd_header_i,
  mem_fwd_data_i,
  mem_fwd_v_i,
  mem_fwd_ready_and_o,
  mem_rev_header_o,
  mem_rev_data_o,
  mem_rev_v_o,
  mem_rev_ready_and_i,
  dma_pkt_o,
  dma_pkt_v_o,
  dma_pkt_ready_and_i,
  dma_data_i,
  dma_data_v_i,
  dma_data_ready_and_o,
  dma_data_o,
  dma_data_v_o,
  dma_data_ready_and_i
);

  input [64:0] mem_fwd_header_i;
  input [127:0] mem_fwd_data_i;
  output [64:0] mem_rev_header_o;
  output [127:0] mem_rev_data_o;
  output [75:0] dma_pkt_o;
  output [1:0] dma_pkt_v_o;
  input [1:0] dma_pkt_ready_and_i;
  input [255:0] dma_data_i;
  input [1:0] dma_data_v_i;
  output [1:0] dma_data_ready_and_o;
  output [255:0] dma_data_o;
  output [1:0] dma_data_v_o;
  input [1:0] dma_data_ready_and_i;
  input clk_i;
  input reset_i;
  input mem_fwd_v_i;
  input mem_rev_ready_and_i;
  output mem_fwd_ready_and_o;
  output mem_rev_v_o;
  wire [64:0] mem_rev_header_o,mem_fwd_header_li;
  wire [127:0] mem_rev_data_o,mem_fwd_data_li;
  wire [75:0] dma_pkt_o;
  wire [1:0] dma_pkt_v_o,dma_data_ready_and_o,dma_data_v_o,cache_pkt_v_li,cache_pkt_yumi_lo,
  cache_data_v_lo,cache_data_yumi_li;
  wire [255:0] dma_data_o,cache_data_lo;
  wire mem_fwd_ready_and_o,mem_rev_v_o,mem_fwd_v_li,_2_net_,mem_fwd_ready_and_lo,
  dma_pkt_lo_1__addr__32_,dma_pkt_lo_1__addr__31_,dma_pkt_lo_1__addr__30_,
  dma_pkt_lo_1__addr__29_,dma_pkt_lo_1__addr__28_,dma_pkt_lo_1__addr__27_,
  dma_pkt_lo_1__addr__26_,dma_pkt_lo_1__addr__25_,dma_pkt_lo_1__addr__24_,dma_pkt_lo_1__addr__23_,
  dma_pkt_lo_1__addr__22_,dma_pkt_lo_1__addr__21_,dma_pkt_lo_1__addr__20_,
  dma_pkt_lo_1__addr__19_,dma_pkt_lo_1__addr__18_,dma_pkt_lo_1__addr__17_,
  dma_pkt_lo_1__addr__16_,dma_pkt_lo_1__addr__15_,dma_pkt_lo_1__addr__14_,dma_pkt_lo_1__addr__13_,
  dma_pkt_lo_1__addr__12_,dma_pkt_lo_1__addr__11_,dma_pkt_lo_1__addr__10_,
  dma_pkt_lo_1__addr__9_,dma_pkt_lo_1__addr__8_,dma_pkt_lo_1__addr__7_,dma_pkt_lo_1__addr__6_,
  dma_pkt_lo_1__addr__5_,dma_pkt_lo_1__addr__4_,dma_pkt_lo_1__addr__3_,
  dma_pkt_lo_1__addr__2_,dma_pkt_lo_1__addr__1_,dma_pkt_lo_1__addr__0_,dma_pkt_lo_0__addr__32_,
  dma_pkt_lo_0__addr__31_,dma_pkt_lo_0__addr__30_,dma_pkt_lo_0__addr__29_,
  dma_pkt_lo_0__addr__28_,dma_pkt_lo_0__addr__27_,dma_pkt_lo_0__addr__26_,
  dma_pkt_lo_0__addr__25_,dma_pkt_lo_0__addr__24_,dma_pkt_lo_0__addr__23_,dma_pkt_lo_0__addr__22_,
  dma_pkt_lo_0__addr__21_,dma_pkt_lo_0__addr__20_,dma_pkt_lo_0__addr__19_,
  dma_pkt_lo_0__addr__18_,dma_pkt_lo_0__addr__17_,dma_pkt_lo_0__addr__16_,
  dma_pkt_lo_0__addr__15_,dma_pkt_lo_0__addr__14_,dma_pkt_lo_0__addr__13_,dma_pkt_lo_0__addr__12_,
  dma_pkt_lo_0__addr__11_,dma_pkt_lo_0__addr__10_,dma_pkt_lo_0__addr__9_,
  dma_pkt_lo_0__addr__8_,dma_pkt_lo_0__addr__7_,dma_pkt_lo_0__addr__6_,
  dma_pkt_lo_0__addr__5_,dma_pkt_lo_0__addr__4_,dma_pkt_lo_0__addr__3_,dma_pkt_lo_0__addr__2_,
  dma_pkt_lo_0__addr__1_,dma_pkt_lo_0__addr__0_,_3_net_,_4_net_,_7_net_,_8_net_;
  wire [365:0] cache_pkt_li;

  bsg_fifo_1r1w_small_000000c1_00000004
  fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(mem_fwd_v_i),
    .ready_param_o(mem_fwd_ready_and_o),
    .data_i({ mem_fwd_data_i, mem_fwd_header_i }),
    .v_o(mem_fwd_v_li),
    .data_o({ mem_fwd_data_li, mem_fwd_header_li }),
    .yumi_i(_2_net_)
  );


  bp_me_cache_controller_00
  cache_controller
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .mem_fwd_header_i(mem_fwd_header_li),
    .mem_fwd_data_i(mem_fwd_data_li),
    .mem_fwd_v_i(mem_fwd_v_li),
    .mem_fwd_ready_and_o(mem_fwd_ready_and_lo),
    .mem_rev_header_o(mem_rev_header_o),
    .mem_rev_data_o(mem_rev_data_o),
    .mem_rev_v_o(mem_rev_v_o),
    .mem_rev_ready_and_i(mem_rev_ready_and_i),
    .cache_pkt_o(cache_pkt_li),
    .cache_pkt_v_o(cache_pkt_v_li),
    .cache_pkt_yumi_i(cache_pkt_yumi_lo),
    .cache_data_i(cache_data_lo),
    .cache_data_v_i(cache_data_v_lo),
    .cache_data_yumi_o(cache_data_yumi_li)
  );


  bsg_cache_00000021_00000080_00000004_00000080_00000008_1_1_00000080
  \bank_0_.cache 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .cache_pkt_i(cache_pkt_li[182:0]),
    .v_i(cache_pkt_v_li[0]),
    .yumi_o(cache_pkt_yumi_lo[0]),
    .data_o(cache_data_lo[127:0]),
    .v_o(cache_data_v_lo[0]),
    .yumi_i(cache_data_yumi_li[0]),
    .dma_pkt_o({ dma_pkt_o[37:37], dma_pkt_lo_0__addr__32_, dma_pkt_lo_0__addr__31_, dma_pkt_lo_0__addr__30_, dma_pkt_lo_0__addr__29_, dma_pkt_lo_0__addr__28_, dma_pkt_lo_0__addr__27_, dma_pkt_lo_0__addr__26_, dma_pkt_lo_0__addr__25_, dma_pkt_lo_0__addr__24_, dma_pkt_lo_0__addr__23_, dma_pkt_lo_0__addr__22_, dma_pkt_lo_0__addr__21_, dma_pkt_lo_0__addr__20_, dma_pkt_lo_0__addr__19_, dma_pkt_lo_0__addr__18_, dma_pkt_lo_0__addr__17_, dma_pkt_lo_0__addr__16_, dma_pkt_lo_0__addr__15_, dma_pkt_lo_0__addr__14_, dma_pkt_lo_0__addr__13_, dma_pkt_lo_0__addr__12_, dma_pkt_lo_0__addr__11_, dma_pkt_lo_0__addr__10_, dma_pkt_lo_0__addr__9_, dma_pkt_lo_0__addr__8_, dma_pkt_lo_0__addr__7_, dma_pkt_lo_0__addr__6_, dma_pkt_lo_0__addr__5_, dma_pkt_lo_0__addr__4_, dma_pkt_lo_0__addr__3_, dma_pkt_lo_0__addr__2_, dma_pkt_lo_0__addr__1_, dma_pkt_lo_0__addr__0_, dma_pkt_o[3:0] }),
    .dma_pkt_v_o(dma_pkt_v_o[0]),
    .dma_pkt_yumi_i(_3_net_),
    .dma_data_i(dma_data_i[127:0]),
    .dma_data_v_i(dma_data_v_i[0]),
    .dma_data_ready_and_o(dma_data_ready_and_o[0]),
    .dma_data_o(dma_data_o[127:0]),
    .dma_data_v_o(dma_data_v_o[0]),
    .dma_data_yumi_i(_4_net_)
  );


  bp_me_dram_hash_decode_00
  \bank_0_.dma_addr_hash_decode 
  (
    .daddr_i({ dma_pkt_lo_0__addr__32_, dma_pkt_lo_0__addr__31_, dma_pkt_lo_0__addr__30_, dma_pkt_lo_0__addr__29_, dma_pkt_lo_0__addr__28_, dma_pkt_lo_0__addr__27_, dma_pkt_lo_0__addr__26_, dma_pkt_lo_0__addr__25_, dma_pkt_lo_0__addr__24_, dma_pkt_lo_0__addr__23_, dma_pkt_lo_0__addr__22_, dma_pkt_lo_0__addr__21_, dma_pkt_lo_0__addr__20_, dma_pkt_lo_0__addr__19_, dma_pkt_lo_0__addr__18_, dma_pkt_lo_0__addr__17_, dma_pkt_lo_0__addr__16_, dma_pkt_lo_0__addr__15_, dma_pkt_lo_0__addr__14_, dma_pkt_lo_0__addr__13_, dma_pkt_lo_0__addr__12_, dma_pkt_lo_0__addr__11_, dma_pkt_lo_0__addr__10_, dma_pkt_lo_0__addr__9_, dma_pkt_lo_0__addr__8_, dma_pkt_lo_0__addr__7_, dma_pkt_lo_0__addr__6_, dma_pkt_lo_0__addr__5_, dma_pkt_lo_0__addr__4_, dma_pkt_lo_0__addr__3_, dma_pkt_lo_0__addr__2_, dma_pkt_lo_0__addr__1_, dma_pkt_lo_0__addr__0_ }),
    .daddr_o(dma_pkt_o[36:4])
  );


  bsg_cache_00000021_00000080_00000004_00000080_00000008_1_1_00000080
  \bank_1_.cache 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .cache_pkt_i(cache_pkt_li[365:183]),
    .v_i(cache_pkt_v_li[1]),
    .yumi_o(cache_pkt_yumi_lo[1]),
    .data_o(cache_data_lo[255:128]),
    .v_o(cache_data_v_lo[1]),
    .yumi_i(cache_data_yumi_li[1]),
    .dma_pkt_o({ dma_pkt_o[75:75], dma_pkt_lo_1__addr__32_, dma_pkt_lo_1__addr__31_, dma_pkt_lo_1__addr__30_, dma_pkt_lo_1__addr__29_, dma_pkt_lo_1__addr__28_, dma_pkt_lo_1__addr__27_, dma_pkt_lo_1__addr__26_, dma_pkt_lo_1__addr__25_, dma_pkt_lo_1__addr__24_, dma_pkt_lo_1__addr__23_, dma_pkt_lo_1__addr__22_, dma_pkt_lo_1__addr__21_, dma_pkt_lo_1__addr__20_, dma_pkt_lo_1__addr__19_, dma_pkt_lo_1__addr__18_, dma_pkt_lo_1__addr__17_, dma_pkt_lo_1__addr__16_, dma_pkt_lo_1__addr__15_, dma_pkt_lo_1__addr__14_, dma_pkt_lo_1__addr__13_, dma_pkt_lo_1__addr__12_, dma_pkt_lo_1__addr__11_, dma_pkt_lo_1__addr__10_, dma_pkt_lo_1__addr__9_, dma_pkt_lo_1__addr__8_, dma_pkt_lo_1__addr__7_, dma_pkt_lo_1__addr__6_, dma_pkt_lo_1__addr__5_, dma_pkt_lo_1__addr__4_, dma_pkt_lo_1__addr__3_, dma_pkt_lo_1__addr__2_, dma_pkt_lo_1__addr__1_, dma_pkt_lo_1__addr__0_, dma_pkt_o[41:38] }),
    .dma_pkt_v_o(dma_pkt_v_o[1]),
    .dma_pkt_yumi_i(_7_net_),
    .dma_data_i(dma_data_i[255:128]),
    .dma_data_v_i(dma_data_v_i[1]),
    .dma_data_ready_and_o(dma_data_ready_and_o[1]),
    .dma_data_o(dma_data_o[255:128]),
    .dma_data_v_o(dma_data_v_o[1]),
    .dma_data_yumi_i(_8_net_)
  );


  bp_me_dram_hash_decode_00
  \bank_1_.dma_addr_hash_decode 
  (
    .daddr_i({ dma_pkt_lo_1__addr__32_, dma_pkt_lo_1__addr__31_, dma_pkt_lo_1__addr__30_, dma_pkt_lo_1__addr__29_, dma_pkt_lo_1__addr__28_, dma_pkt_lo_1__addr__27_, dma_pkt_lo_1__addr__26_, dma_pkt_lo_1__addr__25_, dma_pkt_lo_1__addr__24_, dma_pkt_lo_1__addr__23_, dma_pkt_lo_1__addr__22_, dma_pkt_lo_1__addr__21_, dma_pkt_lo_1__addr__20_, dma_pkt_lo_1__addr__19_, dma_pkt_lo_1__addr__18_, dma_pkt_lo_1__addr__17_, dma_pkt_lo_1__addr__16_, dma_pkt_lo_1__addr__15_, dma_pkt_lo_1__addr__14_, dma_pkt_lo_1__addr__13_, dma_pkt_lo_1__addr__12_, dma_pkt_lo_1__addr__11_, dma_pkt_lo_1__addr__10_, dma_pkt_lo_1__addr__9_, dma_pkt_lo_1__addr__8_, dma_pkt_lo_1__addr__7_, dma_pkt_lo_1__addr__6_, dma_pkt_lo_1__addr__5_, dma_pkt_lo_1__addr__4_, dma_pkt_lo_1__addr__3_, dma_pkt_lo_1__addr__2_, dma_pkt_lo_1__addr__1_, dma_pkt_lo_1__addr__0_ }),
    .daddr_o(dma_pkt_o[74:42])
  );

  assign _2_net_ = mem_fwd_ready_and_lo & mem_fwd_v_li;
  assign _4_net_ = dma_data_ready_and_i[0] & dma_data_v_o[0];
  assign _3_net_ = dma_pkt_ready_and_i[0] & dma_pkt_v_o[0];
  assign _8_net_ = dma_data_ready_and_i[1] & dma_data_v_o[1];
  assign _7_net_ = dma_pkt_ready_and_i[1] & dma_pkt_v_o[1];

endmodule

