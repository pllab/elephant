

module bsg_circular_ptr_slots_p128_max_add_p127
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [6:0] add_i;
  output [6:0] o;
  output [6:0] n_o;
  input clk;
  input reset_i;
  wire [6:0] o,n_o;
  reg o_6_sv2v_reg,o_5_sv2v_reg,o_4_sv2v_reg,o_3_sv2v_reg,o_2_sv2v_reg,o_1_sv2v_reg,
  o_0_sv2v_reg;
  assign o[6] = o_6_sv2v_reg;
  assign o[5] = o_5_sv2v_reg;
  assign o[4] = o_4_sv2v_reg;
  assign o[3] = o_3_sv2v_reg;
  assign o[2] = o_2_sv2v_reg;
  assign o[1] = o_1_sv2v_reg;
  assign o[0] = o_0_sv2v_reg;
  assign n_o = o + add_i;

  always @(posedge clk) begin
    if(reset_i) begin
      o_6_sv2v_reg <= 1'b0;
      o_5_sv2v_reg <= 1'b0;
      o_4_sv2v_reg <= 1'b0;
      o_3_sv2v_reg <= 1'b0;
      o_2_sv2v_reg <= 1'b0;
      o_1_sv2v_reg <= 1'b0;
      o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      o_6_sv2v_reg <= n_o[6];
      o_5_sv2v_reg <= n_o[5];
      o_4_sv2v_reg <= n_o[4];
      o_3_sv2v_reg <= n_o[3];
      o_2_sv2v_reg <= n_o[2];
      o_1_sv2v_reg <= n_o[1];
      o_0_sv2v_reg <= n_o[0];
    end 
  end


endmodule



module bsg_mem_1r1w_synth_00000050_00000008_0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [2:0] w_addr_i;
  input [79:0] w_data_i;
  input [2:0] r_addr_i;
  output [79:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [79:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45;
  wire [639:0] \nz.mem ;
  reg \nz.mem_639_sv2v_reg ,\nz.mem_638_sv2v_reg ,\nz.mem_637_sv2v_reg ,
  \nz.mem_636_sv2v_reg ,\nz.mem_635_sv2v_reg ,\nz.mem_634_sv2v_reg ,\nz.mem_633_sv2v_reg ,
  \nz.mem_632_sv2v_reg ,\nz.mem_631_sv2v_reg ,\nz.mem_630_sv2v_reg ,
  \nz.mem_629_sv2v_reg ,\nz.mem_628_sv2v_reg ,\nz.mem_627_sv2v_reg ,\nz.mem_626_sv2v_reg ,
  \nz.mem_625_sv2v_reg ,\nz.mem_624_sv2v_reg ,\nz.mem_623_sv2v_reg ,\nz.mem_622_sv2v_reg ,
  \nz.mem_621_sv2v_reg ,\nz.mem_620_sv2v_reg ,\nz.mem_619_sv2v_reg ,
  \nz.mem_618_sv2v_reg ,\nz.mem_617_sv2v_reg ,\nz.mem_616_sv2v_reg ,\nz.mem_615_sv2v_reg ,
  \nz.mem_614_sv2v_reg ,\nz.mem_613_sv2v_reg ,\nz.mem_612_sv2v_reg ,\nz.mem_611_sv2v_reg ,
  \nz.mem_610_sv2v_reg ,\nz.mem_609_sv2v_reg ,\nz.mem_608_sv2v_reg ,
  \nz.mem_607_sv2v_reg ,\nz.mem_606_sv2v_reg ,\nz.mem_605_sv2v_reg ,\nz.mem_604_sv2v_reg ,
  \nz.mem_603_sv2v_reg ,\nz.mem_602_sv2v_reg ,\nz.mem_601_sv2v_reg ,\nz.mem_600_sv2v_reg ,
  \nz.mem_599_sv2v_reg ,\nz.mem_598_sv2v_reg ,\nz.mem_597_sv2v_reg ,
  \nz.mem_596_sv2v_reg ,\nz.mem_595_sv2v_reg ,\nz.mem_594_sv2v_reg ,\nz.mem_593_sv2v_reg ,
  \nz.mem_592_sv2v_reg ,\nz.mem_591_sv2v_reg ,\nz.mem_590_sv2v_reg ,
  \nz.mem_589_sv2v_reg ,\nz.mem_588_sv2v_reg ,\nz.mem_587_sv2v_reg ,\nz.mem_586_sv2v_reg ,
  \nz.mem_585_sv2v_reg ,\nz.mem_584_sv2v_reg ,\nz.mem_583_sv2v_reg ,\nz.mem_582_sv2v_reg ,
  \nz.mem_581_sv2v_reg ,\nz.mem_580_sv2v_reg ,\nz.mem_579_sv2v_reg ,
  \nz.mem_578_sv2v_reg ,\nz.mem_577_sv2v_reg ,\nz.mem_576_sv2v_reg ,\nz.mem_575_sv2v_reg ,
  \nz.mem_574_sv2v_reg ,\nz.mem_573_sv2v_reg ,\nz.mem_572_sv2v_reg ,\nz.mem_571_sv2v_reg ,
  \nz.mem_570_sv2v_reg ,\nz.mem_569_sv2v_reg ,\nz.mem_568_sv2v_reg ,
  \nz.mem_567_sv2v_reg ,\nz.mem_566_sv2v_reg ,\nz.mem_565_sv2v_reg ,\nz.mem_564_sv2v_reg ,
  \nz.mem_563_sv2v_reg ,\nz.mem_562_sv2v_reg ,\nz.mem_561_sv2v_reg ,\nz.mem_560_sv2v_reg ,
  \nz.mem_559_sv2v_reg ,\nz.mem_558_sv2v_reg ,\nz.mem_557_sv2v_reg ,
  \nz.mem_556_sv2v_reg ,\nz.mem_555_sv2v_reg ,\nz.mem_554_sv2v_reg ,\nz.mem_553_sv2v_reg ,
  \nz.mem_552_sv2v_reg ,\nz.mem_551_sv2v_reg ,\nz.mem_550_sv2v_reg ,
  \nz.mem_549_sv2v_reg ,\nz.mem_548_sv2v_reg ,\nz.mem_547_sv2v_reg ,\nz.mem_546_sv2v_reg ,
  \nz.mem_545_sv2v_reg ,\nz.mem_544_sv2v_reg ,\nz.mem_543_sv2v_reg ,\nz.mem_542_sv2v_reg ,
  \nz.mem_541_sv2v_reg ,\nz.mem_540_sv2v_reg ,\nz.mem_539_sv2v_reg ,
  \nz.mem_538_sv2v_reg ,\nz.mem_537_sv2v_reg ,\nz.mem_536_sv2v_reg ,\nz.mem_535_sv2v_reg ,
  \nz.mem_534_sv2v_reg ,\nz.mem_533_sv2v_reg ,\nz.mem_532_sv2v_reg ,\nz.mem_531_sv2v_reg ,
  \nz.mem_530_sv2v_reg ,\nz.mem_529_sv2v_reg ,\nz.mem_528_sv2v_reg ,
  \nz.mem_527_sv2v_reg ,\nz.mem_526_sv2v_reg ,\nz.mem_525_sv2v_reg ,\nz.mem_524_sv2v_reg ,
  \nz.mem_523_sv2v_reg ,\nz.mem_522_sv2v_reg ,\nz.mem_521_sv2v_reg ,\nz.mem_520_sv2v_reg ,
  \nz.mem_519_sv2v_reg ,\nz.mem_518_sv2v_reg ,\nz.mem_517_sv2v_reg ,
  \nz.mem_516_sv2v_reg ,\nz.mem_515_sv2v_reg ,\nz.mem_514_sv2v_reg ,\nz.mem_513_sv2v_reg ,
  \nz.mem_512_sv2v_reg ,\nz.mem_511_sv2v_reg ,\nz.mem_510_sv2v_reg ,
  \nz.mem_509_sv2v_reg ,\nz.mem_508_sv2v_reg ,\nz.mem_507_sv2v_reg ,\nz.mem_506_sv2v_reg ,
  \nz.mem_505_sv2v_reg ,\nz.mem_504_sv2v_reg ,\nz.mem_503_sv2v_reg ,\nz.mem_502_sv2v_reg ,
  \nz.mem_501_sv2v_reg ,\nz.mem_500_sv2v_reg ,\nz.mem_499_sv2v_reg ,
  \nz.mem_498_sv2v_reg ,\nz.mem_497_sv2v_reg ,\nz.mem_496_sv2v_reg ,\nz.mem_495_sv2v_reg ,
  \nz.mem_494_sv2v_reg ,\nz.mem_493_sv2v_reg ,\nz.mem_492_sv2v_reg ,\nz.mem_491_sv2v_reg ,
  \nz.mem_490_sv2v_reg ,\nz.mem_489_sv2v_reg ,\nz.mem_488_sv2v_reg ,
  \nz.mem_487_sv2v_reg ,\nz.mem_486_sv2v_reg ,\nz.mem_485_sv2v_reg ,\nz.mem_484_sv2v_reg ,
  \nz.mem_483_sv2v_reg ,\nz.mem_482_sv2v_reg ,\nz.mem_481_sv2v_reg ,\nz.mem_480_sv2v_reg ,
  \nz.mem_479_sv2v_reg ,\nz.mem_478_sv2v_reg ,\nz.mem_477_sv2v_reg ,
  \nz.mem_476_sv2v_reg ,\nz.mem_475_sv2v_reg ,\nz.mem_474_sv2v_reg ,\nz.mem_473_sv2v_reg ,
  \nz.mem_472_sv2v_reg ,\nz.mem_471_sv2v_reg ,\nz.mem_470_sv2v_reg ,
  \nz.mem_469_sv2v_reg ,\nz.mem_468_sv2v_reg ,\nz.mem_467_sv2v_reg ,\nz.mem_466_sv2v_reg ,
  \nz.mem_465_sv2v_reg ,\nz.mem_464_sv2v_reg ,\nz.mem_463_sv2v_reg ,\nz.mem_462_sv2v_reg ,
  \nz.mem_461_sv2v_reg ,\nz.mem_460_sv2v_reg ,\nz.mem_459_sv2v_reg ,
  \nz.mem_458_sv2v_reg ,\nz.mem_457_sv2v_reg ,\nz.mem_456_sv2v_reg ,\nz.mem_455_sv2v_reg ,
  \nz.mem_454_sv2v_reg ,\nz.mem_453_sv2v_reg ,\nz.mem_452_sv2v_reg ,\nz.mem_451_sv2v_reg ,
  \nz.mem_450_sv2v_reg ,\nz.mem_449_sv2v_reg ,\nz.mem_448_sv2v_reg ,
  \nz.mem_447_sv2v_reg ,\nz.mem_446_sv2v_reg ,\nz.mem_445_sv2v_reg ,\nz.mem_444_sv2v_reg ,
  \nz.mem_443_sv2v_reg ,\nz.mem_442_sv2v_reg ,\nz.mem_441_sv2v_reg ,\nz.mem_440_sv2v_reg ,
  \nz.mem_439_sv2v_reg ,\nz.mem_438_sv2v_reg ,\nz.mem_437_sv2v_reg ,
  \nz.mem_436_sv2v_reg ,\nz.mem_435_sv2v_reg ,\nz.mem_434_sv2v_reg ,\nz.mem_433_sv2v_reg ,
  \nz.mem_432_sv2v_reg ,\nz.mem_431_sv2v_reg ,\nz.mem_430_sv2v_reg ,
  \nz.mem_429_sv2v_reg ,\nz.mem_428_sv2v_reg ,\nz.mem_427_sv2v_reg ,\nz.mem_426_sv2v_reg ,
  \nz.mem_425_sv2v_reg ,\nz.mem_424_sv2v_reg ,\nz.mem_423_sv2v_reg ,\nz.mem_422_sv2v_reg ,
  \nz.mem_421_sv2v_reg ,\nz.mem_420_sv2v_reg ,\nz.mem_419_sv2v_reg ,
  \nz.mem_418_sv2v_reg ,\nz.mem_417_sv2v_reg ,\nz.mem_416_sv2v_reg ,\nz.mem_415_sv2v_reg ,
  \nz.mem_414_sv2v_reg ,\nz.mem_413_sv2v_reg ,\nz.mem_412_sv2v_reg ,\nz.mem_411_sv2v_reg ,
  \nz.mem_410_sv2v_reg ,\nz.mem_409_sv2v_reg ,\nz.mem_408_sv2v_reg ,
  \nz.mem_407_sv2v_reg ,\nz.mem_406_sv2v_reg ,\nz.mem_405_sv2v_reg ,\nz.mem_404_sv2v_reg ,
  \nz.mem_403_sv2v_reg ,\nz.mem_402_sv2v_reg ,\nz.mem_401_sv2v_reg ,\nz.mem_400_sv2v_reg ,
  \nz.mem_399_sv2v_reg ,\nz.mem_398_sv2v_reg ,\nz.mem_397_sv2v_reg ,
  \nz.mem_396_sv2v_reg ,\nz.mem_395_sv2v_reg ,\nz.mem_394_sv2v_reg ,\nz.mem_393_sv2v_reg ,
  \nz.mem_392_sv2v_reg ,\nz.mem_391_sv2v_reg ,\nz.mem_390_sv2v_reg ,
  \nz.mem_389_sv2v_reg ,\nz.mem_388_sv2v_reg ,\nz.mem_387_sv2v_reg ,\nz.mem_386_sv2v_reg ,
  \nz.mem_385_sv2v_reg ,\nz.mem_384_sv2v_reg ,\nz.mem_383_sv2v_reg ,\nz.mem_382_sv2v_reg ,
  \nz.mem_381_sv2v_reg ,\nz.mem_380_sv2v_reg ,\nz.mem_379_sv2v_reg ,
  \nz.mem_378_sv2v_reg ,\nz.mem_377_sv2v_reg ,\nz.mem_376_sv2v_reg ,\nz.mem_375_sv2v_reg ,
  \nz.mem_374_sv2v_reg ,\nz.mem_373_sv2v_reg ,\nz.mem_372_sv2v_reg ,\nz.mem_371_sv2v_reg ,
  \nz.mem_370_sv2v_reg ,\nz.mem_369_sv2v_reg ,\nz.mem_368_sv2v_reg ,
  \nz.mem_367_sv2v_reg ,\nz.mem_366_sv2v_reg ,\nz.mem_365_sv2v_reg ,\nz.mem_364_sv2v_reg ,
  \nz.mem_363_sv2v_reg ,\nz.mem_362_sv2v_reg ,\nz.mem_361_sv2v_reg ,\nz.mem_360_sv2v_reg ,
  \nz.mem_359_sv2v_reg ,\nz.mem_358_sv2v_reg ,\nz.mem_357_sv2v_reg ,
  \nz.mem_356_sv2v_reg ,\nz.mem_355_sv2v_reg ,\nz.mem_354_sv2v_reg ,\nz.mem_353_sv2v_reg ,
  \nz.mem_352_sv2v_reg ,\nz.mem_351_sv2v_reg ,\nz.mem_350_sv2v_reg ,
  \nz.mem_349_sv2v_reg ,\nz.mem_348_sv2v_reg ,\nz.mem_347_sv2v_reg ,\nz.mem_346_sv2v_reg ,
  \nz.mem_345_sv2v_reg ,\nz.mem_344_sv2v_reg ,\nz.mem_343_sv2v_reg ,\nz.mem_342_sv2v_reg ,
  \nz.mem_341_sv2v_reg ,\nz.mem_340_sv2v_reg ,\nz.mem_339_sv2v_reg ,
  \nz.mem_338_sv2v_reg ,\nz.mem_337_sv2v_reg ,\nz.mem_336_sv2v_reg ,\nz.mem_335_sv2v_reg ,
  \nz.mem_334_sv2v_reg ,\nz.mem_333_sv2v_reg ,\nz.mem_332_sv2v_reg ,\nz.mem_331_sv2v_reg ,
  \nz.mem_330_sv2v_reg ,\nz.mem_329_sv2v_reg ,\nz.mem_328_sv2v_reg ,
  \nz.mem_327_sv2v_reg ,\nz.mem_326_sv2v_reg ,\nz.mem_325_sv2v_reg ,\nz.mem_324_sv2v_reg ,
  \nz.mem_323_sv2v_reg ,\nz.mem_322_sv2v_reg ,\nz.mem_321_sv2v_reg ,\nz.mem_320_sv2v_reg ,
  \nz.mem_319_sv2v_reg ,\nz.mem_318_sv2v_reg ,\nz.mem_317_sv2v_reg ,
  \nz.mem_316_sv2v_reg ,\nz.mem_315_sv2v_reg ,\nz.mem_314_sv2v_reg ,\nz.mem_313_sv2v_reg ,
  \nz.mem_312_sv2v_reg ,\nz.mem_311_sv2v_reg ,\nz.mem_310_sv2v_reg ,
  \nz.mem_309_sv2v_reg ,\nz.mem_308_sv2v_reg ,\nz.mem_307_sv2v_reg ,\nz.mem_306_sv2v_reg ,
  \nz.mem_305_sv2v_reg ,\nz.mem_304_sv2v_reg ,\nz.mem_303_sv2v_reg ,\nz.mem_302_sv2v_reg ,
  \nz.mem_301_sv2v_reg ,\nz.mem_300_sv2v_reg ,\nz.mem_299_sv2v_reg ,
  \nz.mem_298_sv2v_reg ,\nz.mem_297_sv2v_reg ,\nz.mem_296_sv2v_reg ,\nz.mem_295_sv2v_reg ,
  \nz.mem_294_sv2v_reg ,\nz.mem_293_sv2v_reg ,\nz.mem_292_sv2v_reg ,\nz.mem_291_sv2v_reg ,
  \nz.mem_290_sv2v_reg ,\nz.mem_289_sv2v_reg ,\nz.mem_288_sv2v_reg ,
  \nz.mem_287_sv2v_reg ,\nz.mem_286_sv2v_reg ,\nz.mem_285_sv2v_reg ,\nz.mem_284_sv2v_reg ,
  \nz.mem_283_sv2v_reg ,\nz.mem_282_sv2v_reg ,\nz.mem_281_sv2v_reg ,\nz.mem_280_sv2v_reg ,
  \nz.mem_279_sv2v_reg ,\nz.mem_278_sv2v_reg ,\nz.mem_277_sv2v_reg ,
  \nz.mem_276_sv2v_reg ,\nz.mem_275_sv2v_reg ,\nz.mem_274_sv2v_reg ,\nz.mem_273_sv2v_reg ,
  \nz.mem_272_sv2v_reg ,\nz.mem_271_sv2v_reg ,\nz.mem_270_sv2v_reg ,
  \nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,\nz.mem_267_sv2v_reg ,\nz.mem_266_sv2v_reg ,
  \nz.mem_265_sv2v_reg ,\nz.mem_264_sv2v_reg ,\nz.mem_263_sv2v_reg ,\nz.mem_262_sv2v_reg ,
  \nz.mem_261_sv2v_reg ,\nz.mem_260_sv2v_reg ,\nz.mem_259_sv2v_reg ,
  \nz.mem_258_sv2v_reg ,\nz.mem_257_sv2v_reg ,\nz.mem_256_sv2v_reg ,\nz.mem_255_sv2v_reg ,
  \nz.mem_254_sv2v_reg ,\nz.mem_253_sv2v_reg ,\nz.mem_252_sv2v_reg ,\nz.mem_251_sv2v_reg ,
  \nz.mem_250_sv2v_reg ,\nz.mem_249_sv2v_reg ,\nz.mem_248_sv2v_reg ,
  \nz.mem_247_sv2v_reg ,\nz.mem_246_sv2v_reg ,\nz.mem_245_sv2v_reg ,\nz.mem_244_sv2v_reg ,
  \nz.mem_243_sv2v_reg ,\nz.mem_242_sv2v_reg ,\nz.mem_241_sv2v_reg ,\nz.mem_240_sv2v_reg ,
  \nz.mem_239_sv2v_reg ,\nz.mem_238_sv2v_reg ,\nz.mem_237_sv2v_reg ,
  \nz.mem_236_sv2v_reg ,\nz.mem_235_sv2v_reg ,\nz.mem_234_sv2v_reg ,\nz.mem_233_sv2v_reg ,
  \nz.mem_232_sv2v_reg ,\nz.mem_231_sv2v_reg ,\nz.mem_230_sv2v_reg ,
  \nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,\nz.mem_227_sv2v_reg ,\nz.mem_226_sv2v_reg ,
  \nz.mem_225_sv2v_reg ,\nz.mem_224_sv2v_reg ,\nz.mem_223_sv2v_reg ,\nz.mem_222_sv2v_reg ,
  \nz.mem_221_sv2v_reg ,\nz.mem_220_sv2v_reg ,\nz.mem_219_sv2v_reg ,
  \nz.mem_218_sv2v_reg ,\nz.mem_217_sv2v_reg ,\nz.mem_216_sv2v_reg ,\nz.mem_215_sv2v_reg ,
  \nz.mem_214_sv2v_reg ,\nz.mem_213_sv2v_reg ,\nz.mem_212_sv2v_reg ,\nz.mem_211_sv2v_reg ,
  \nz.mem_210_sv2v_reg ,\nz.mem_209_sv2v_reg ,\nz.mem_208_sv2v_reg ,
  \nz.mem_207_sv2v_reg ,\nz.mem_206_sv2v_reg ,\nz.mem_205_sv2v_reg ,\nz.mem_204_sv2v_reg ,
  \nz.mem_203_sv2v_reg ,\nz.mem_202_sv2v_reg ,\nz.mem_201_sv2v_reg ,\nz.mem_200_sv2v_reg ,
  \nz.mem_199_sv2v_reg ,\nz.mem_198_sv2v_reg ,\nz.mem_197_sv2v_reg ,
  \nz.mem_196_sv2v_reg ,\nz.mem_195_sv2v_reg ,\nz.mem_194_sv2v_reg ,\nz.mem_193_sv2v_reg ,
  \nz.mem_192_sv2v_reg ,\nz.mem_191_sv2v_reg ,\nz.mem_190_sv2v_reg ,
  \nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,\nz.mem_187_sv2v_reg ,\nz.mem_186_sv2v_reg ,
  \nz.mem_185_sv2v_reg ,\nz.mem_184_sv2v_reg ,\nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,
  \nz.mem_181_sv2v_reg ,\nz.mem_180_sv2v_reg ,\nz.mem_179_sv2v_reg ,
  \nz.mem_178_sv2v_reg ,\nz.mem_177_sv2v_reg ,\nz.mem_176_sv2v_reg ,\nz.mem_175_sv2v_reg ,
  \nz.mem_174_sv2v_reg ,\nz.mem_173_sv2v_reg ,\nz.mem_172_sv2v_reg ,\nz.mem_171_sv2v_reg ,
  \nz.mem_170_sv2v_reg ,\nz.mem_169_sv2v_reg ,\nz.mem_168_sv2v_reg ,
  \nz.mem_167_sv2v_reg ,\nz.mem_166_sv2v_reg ,\nz.mem_165_sv2v_reg ,\nz.mem_164_sv2v_reg ,
  \nz.mem_163_sv2v_reg ,\nz.mem_162_sv2v_reg ,\nz.mem_161_sv2v_reg ,\nz.mem_160_sv2v_reg ,
  \nz.mem_159_sv2v_reg ,\nz.mem_158_sv2v_reg ,\nz.mem_157_sv2v_reg ,
  \nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,\nz.mem_154_sv2v_reg ,\nz.mem_153_sv2v_reg ,
  \nz.mem_152_sv2v_reg ,\nz.mem_151_sv2v_reg ,\nz.mem_150_sv2v_reg ,
  \nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,\nz.mem_147_sv2v_reg ,\nz.mem_146_sv2v_reg ,
  \nz.mem_145_sv2v_reg ,\nz.mem_144_sv2v_reg ,\nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,
  \nz.mem_141_sv2v_reg ,\nz.mem_140_sv2v_reg ,\nz.mem_139_sv2v_reg ,
  \nz.mem_138_sv2v_reg ,\nz.mem_137_sv2v_reg ,\nz.mem_136_sv2v_reg ,\nz.mem_135_sv2v_reg ,
  \nz.mem_134_sv2v_reg ,\nz.mem_133_sv2v_reg ,\nz.mem_132_sv2v_reg ,\nz.mem_131_sv2v_reg ,
  \nz.mem_130_sv2v_reg ,\nz.mem_129_sv2v_reg ,\nz.mem_128_sv2v_reg ,
  \nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,\nz.mem_125_sv2v_reg ,\nz.mem_124_sv2v_reg ,
  \nz.mem_123_sv2v_reg ,\nz.mem_122_sv2v_reg ,\nz.mem_121_sv2v_reg ,\nz.mem_120_sv2v_reg ,
  \nz.mem_119_sv2v_reg ,\nz.mem_118_sv2v_reg ,\nz.mem_117_sv2v_reg ,
  \nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,\nz.mem_114_sv2v_reg ,\nz.mem_113_sv2v_reg ,
  \nz.mem_112_sv2v_reg ,\nz.mem_111_sv2v_reg ,\nz.mem_110_sv2v_reg ,
  \nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,\nz.mem_107_sv2v_reg ,\nz.mem_106_sv2v_reg ,
  \nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,\nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,
  \nz.mem_101_sv2v_reg ,\nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,
  \nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,\nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,
  \nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,\nz.mem_92_sv2v_reg ,\nz.mem_91_sv2v_reg ,
  \nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,\nz.mem_88_sv2v_reg ,\nz.mem_87_sv2v_reg ,
  \nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,\nz.mem_83_sv2v_reg ,
  \nz.mem_82_sv2v_reg ,\nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,
  \nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,\nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,
  \nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,\nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,
  \nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,\nz.mem_69_sv2v_reg ,\nz.mem_68_sv2v_reg ,
  \nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,
  \nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,\nz.mem_60_sv2v_reg ,
  \nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,
  \nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,
  \nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,
  \nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,
  \nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,\nz.mem_41_sv2v_reg ,
  \nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,
  \nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,
  \nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,
  \nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,
  \nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,\nz.mem_22_sv2v_reg ,
  \nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,
  \nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,
  \nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,
  \nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,
  \nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,
  \nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.mem [639] = \nz.mem_639_sv2v_reg ;
  assign \nz.mem [638] = \nz.mem_638_sv2v_reg ;
  assign \nz.mem [637] = \nz.mem_637_sv2v_reg ;
  assign \nz.mem [636] = \nz.mem_636_sv2v_reg ;
  assign \nz.mem [635] = \nz.mem_635_sv2v_reg ;
  assign \nz.mem [634] = \nz.mem_634_sv2v_reg ;
  assign \nz.mem [633] = \nz.mem_633_sv2v_reg ;
  assign \nz.mem [632] = \nz.mem_632_sv2v_reg ;
  assign \nz.mem [631] = \nz.mem_631_sv2v_reg ;
  assign \nz.mem [630] = \nz.mem_630_sv2v_reg ;
  assign \nz.mem [629] = \nz.mem_629_sv2v_reg ;
  assign \nz.mem [628] = \nz.mem_628_sv2v_reg ;
  assign \nz.mem [627] = \nz.mem_627_sv2v_reg ;
  assign \nz.mem [626] = \nz.mem_626_sv2v_reg ;
  assign \nz.mem [625] = \nz.mem_625_sv2v_reg ;
  assign \nz.mem [624] = \nz.mem_624_sv2v_reg ;
  assign \nz.mem [623] = \nz.mem_623_sv2v_reg ;
  assign \nz.mem [622] = \nz.mem_622_sv2v_reg ;
  assign \nz.mem [621] = \nz.mem_621_sv2v_reg ;
  assign \nz.mem [620] = \nz.mem_620_sv2v_reg ;
  assign \nz.mem [619] = \nz.mem_619_sv2v_reg ;
  assign \nz.mem [618] = \nz.mem_618_sv2v_reg ;
  assign \nz.mem [617] = \nz.mem_617_sv2v_reg ;
  assign \nz.mem [616] = \nz.mem_616_sv2v_reg ;
  assign \nz.mem [615] = \nz.mem_615_sv2v_reg ;
  assign \nz.mem [614] = \nz.mem_614_sv2v_reg ;
  assign \nz.mem [613] = \nz.mem_613_sv2v_reg ;
  assign \nz.mem [612] = \nz.mem_612_sv2v_reg ;
  assign \nz.mem [611] = \nz.mem_611_sv2v_reg ;
  assign \nz.mem [610] = \nz.mem_610_sv2v_reg ;
  assign \nz.mem [609] = \nz.mem_609_sv2v_reg ;
  assign \nz.mem [608] = \nz.mem_608_sv2v_reg ;
  assign \nz.mem [607] = \nz.mem_607_sv2v_reg ;
  assign \nz.mem [606] = \nz.mem_606_sv2v_reg ;
  assign \nz.mem [605] = \nz.mem_605_sv2v_reg ;
  assign \nz.mem [604] = \nz.mem_604_sv2v_reg ;
  assign \nz.mem [603] = \nz.mem_603_sv2v_reg ;
  assign \nz.mem [602] = \nz.mem_602_sv2v_reg ;
  assign \nz.mem [601] = \nz.mem_601_sv2v_reg ;
  assign \nz.mem [600] = \nz.mem_600_sv2v_reg ;
  assign \nz.mem [599] = \nz.mem_599_sv2v_reg ;
  assign \nz.mem [598] = \nz.mem_598_sv2v_reg ;
  assign \nz.mem [597] = \nz.mem_597_sv2v_reg ;
  assign \nz.mem [596] = \nz.mem_596_sv2v_reg ;
  assign \nz.mem [595] = \nz.mem_595_sv2v_reg ;
  assign \nz.mem [594] = \nz.mem_594_sv2v_reg ;
  assign \nz.mem [593] = \nz.mem_593_sv2v_reg ;
  assign \nz.mem [592] = \nz.mem_592_sv2v_reg ;
  assign \nz.mem [591] = \nz.mem_591_sv2v_reg ;
  assign \nz.mem [590] = \nz.mem_590_sv2v_reg ;
  assign \nz.mem [589] = \nz.mem_589_sv2v_reg ;
  assign \nz.mem [588] = \nz.mem_588_sv2v_reg ;
  assign \nz.mem [587] = \nz.mem_587_sv2v_reg ;
  assign \nz.mem [586] = \nz.mem_586_sv2v_reg ;
  assign \nz.mem [585] = \nz.mem_585_sv2v_reg ;
  assign \nz.mem [584] = \nz.mem_584_sv2v_reg ;
  assign \nz.mem [583] = \nz.mem_583_sv2v_reg ;
  assign \nz.mem [582] = \nz.mem_582_sv2v_reg ;
  assign \nz.mem [581] = \nz.mem_581_sv2v_reg ;
  assign \nz.mem [580] = \nz.mem_580_sv2v_reg ;
  assign \nz.mem [579] = \nz.mem_579_sv2v_reg ;
  assign \nz.mem [578] = \nz.mem_578_sv2v_reg ;
  assign \nz.mem [577] = \nz.mem_577_sv2v_reg ;
  assign \nz.mem [576] = \nz.mem_576_sv2v_reg ;
  assign \nz.mem [575] = \nz.mem_575_sv2v_reg ;
  assign \nz.mem [574] = \nz.mem_574_sv2v_reg ;
  assign \nz.mem [573] = \nz.mem_573_sv2v_reg ;
  assign \nz.mem [572] = \nz.mem_572_sv2v_reg ;
  assign \nz.mem [571] = \nz.mem_571_sv2v_reg ;
  assign \nz.mem [570] = \nz.mem_570_sv2v_reg ;
  assign \nz.mem [569] = \nz.mem_569_sv2v_reg ;
  assign \nz.mem [568] = \nz.mem_568_sv2v_reg ;
  assign \nz.mem [567] = \nz.mem_567_sv2v_reg ;
  assign \nz.mem [566] = \nz.mem_566_sv2v_reg ;
  assign \nz.mem [565] = \nz.mem_565_sv2v_reg ;
  assign \nz.mem [564] = \nz.mem_564_sv2v_reg ;
  assign \nz.mem [563] = \nz.mem_563_sv2v_reg ;
  assign \nz.mem [562] = \nz.mem_562_sv2v_reg ;
  assign \nz.mem [561] = \nz.mem_561_sv2v_reg ;
  assign \nz.mem [560] = \nz.mem_560_sv2v_reg ;
  assign \nz.mem [559] = \nz.mem_559_sv2v_reg ;
  assign \nz.mem [558] = \nz.mem_558_sv2v_reg ;
  assign \nz.mem [557] = \nz.mem_557_sv2v_reg ;
  assign \nz.mem [556] = \nz.mem_556_sv2v_reg ;
  assign \nz.mem [555] = \nz.mem_555_sv2v_reg ;
  assign \nz.mem [554] = \nz.mem_554_sv2v_reg ;
  assign \nz.mem [553] = \nz.mem_553_sv2v_reg ;
  assign \nz.mem [552] = \nz.mem_552_sv2v_reg ;
  assign \nz.mem [551] = \nz.mem_551_sv2v_reg ;
  assign \nz.mem [550] = \nz.mem_550_sv2v_reg ;
  assign \nz.mem [549] = \nz.mem_549_sv2v_reg ;
  assign \nz.mem [548] = \nz.mem_548_sv2v_reg ;
  assign \nz.mem [547] = \nz.mem_547_sv2v_reg ;
  assign \nz.mem [546] = \nz.mem_546_sv2v_reg ;
  assign \nz.mem [545] = \nz.mem_545_sv2v_reg ;
  assign \nz.mem [544] = \nz.mem_544_sv2v_reg ;
  assign \nz.mem [543] = \nz.mem_543_sv2v_reg ;
  assign \nz.mem [542] = \nz.mem_542_sv2v_reg ;
  assign \nz.mem [541] = \nz.mem_541_sv2v_reg ;
  assign \nz.mem [540] = \nz.mem_540_sv2v_reg ;
  assign \nz.mem [539] = \nz.mem_539_sv2v_reg ;
  assign \nz.mem [538] = \nz.mem_538_sv2v_reg ;
  assign \nz.mem [537] = \nz.mem_537_sv2v_reg ;
  assign \nz.mem [536] = \nz.mem_536_sv2v_reg ;
  assign \nz.mem [535] = \nz.mem_535_sv2v_reg ;
  assign \nz.mem [534] = \nz.mem_534_sv2v_reg ;
  assign \nz.mem [533] = \nz.mem_533_sv2v_reg ;
  assign \nz.mem [532] = \nz.mem_532_sv2v_reg ;
  assign \nz.mem [531] = \nz.mem_531_sv2v_reg ;
  assign \nz.mem [530] = \nz.mem_530_sv2v_reg ;
  assign \nz.mem [529] = \nz.mem_529_sv2v_reg ;
  assign \nz.mem [528] = \nz.mem_528_sv2v_reg ;
  assign \nz.mem [527] = \nz.mem_527_sv2v_reg ;
  assign \nz.mem [526] = \nz.mem_526_sv2v_reg ;
  assign \nz.mem [525] = \nz.mem_525_sv2v_reg ;
  assign \nz.mem [524] = \nz.mem_524_sv2v_reg ;
  assign \nz.mem [523] = \nz.mem_523_sv2v_reg ;
  assign \nz.mem [522] = \nz.mem_522_sv2v_reg ;
  assign \nz.mem [521] = \nz.mem_521_sv2v_reg ;
  assign \nz.mem [520] = \nz.mem_520_sv2v_reg ;
  assign \nz.mem [519] = \nz.mem_519_sv2v_reg ;
  assign \nz.mem [518] = \nz.mem_518_sv2v_reg ;
  assign \nz.mem [517] = \nz.mem_517_sv2v_reg ;
  assign \nz.mem [516] = \nz.mem_516_sv2v_reg ;
  assign \nz.mem [515] = \nz.mem_515_sv2v_reg ;
  assign \nz.mem [514] = \nz.mem_514_sv2v_reg ;
  assign \nz.mem [513] = \nz.mem_513_sv2v_reg ;
  assign \nz.mem [512] = \nz.mem_512_sv2v_reg ;
  assign \nz.mem [511] = \nz.mem_511_sv2v_reg ;
  assign \nz.mem [510] = \nz.mem_510_sv2v_reg ;
  assign \nz.mem [509] = \nz.mem_509_sv2v_reg ;
  assign \nz.mem [508] = \nz.mem_508_sv2v_reg ;
  assign \nz.mem [507] = \nz.mem_507_sv2v_reg ;
  assign \nz.mem [506] = \nz.mem_506_sv2v_reg ;
  assign \nz.mem [505] = \nz.mem_505_sv2v_reg ;
  assign \nz.mem [504] = \nz.mem_504_sv2v_reg ;
  assign \nz.mem [503] = \nz.mem_503_sv2v_reg ;
  assign \nz.mem [502] = \nz.mem_502_sv2v_reg ;
  assign \nz.mem [501] = \nz.mem_501_sv2v_reg ;
  assign \nz.mem [500] = \nz.mem_500_sv2v_reg ;
  assign \nz.mem [499] = \nz.mem_499_sv2v_reg ;
  assign \nz.mem [498] = \nz.mem_498_sv2v_reg ;
  assign \nz.mem [497] = \nz.mem_497_sv2v_reg ;
  assign \nz.mem [496] = \nz.mem_496_sv2v_reg ;
  assign \nz.mem [495] = \nz.mem_495_sv2v_reg ;
  assign \nz.mem [494] = \nz.mem_494_sv2v_reg ;
  assign \nz.mem [493] = \nz.mem_493_sv2v_reg ;
  assign \nz.mem [492] = \nz.mem_492_sv2v_reg ;
  assign \nz.mem [491] = \nz.mem_491_sv2v_reg ;
  assign \nz.mem [490] = \nz.mem_490_sv2v_reg ;
  assign \nz.mem [489] = \nz.mem_489_sv2v_reg ;
  assign \nz.mem [488] = \nz.mem_488_sv2v_reg ;
  assign \nz.mem [487] = \nz.mem_487_sv2v_reg ;
  assign \nz.mem [486] = \nz.mem_486_sv2v_reg ;
  assign \nz.mem [485] = \nz.mem_485_sv2v_reg ;
  assign \nz.mem [484] = \nz.mem_484_sv2v_reg ;
  assign \nz.mem [483] = \nz.mem_483_sv2v_reg ;
  assign \nz.mem [482] = \nz.mem_482_sv2v_reg ;
  assign \nz.mem [481] = \nz.mem_481_sv2v_reg ;
  assign \nz.mem [480] = \nz.mem_480_sv2v_reg ;
  assign \nz.mem [479] = \nz.mem_479_sv2v_reg ;
  assign \nz.mem [478] = \nz.mem_478_sv2v_reg ;
  assign \nz.mem [477] = \nz.mem_477_sv2v_reg ;
  assign \nz.mem [476] = \nz.mem_476_sv2v_reg ;
  assign \nz.mem [475] = \nz.mem_475_sv2v_reg ;
  assign \nz.mem [474] = \nz.mem_474_sv2v_reg ;
  assign \nz.mem [473] = \nz.mem_473_sv2v_reg ;
  assign \nz.mem [472] = \nz.mem_472_sv2v_reg ;
  assign \nz.mem [471] = \nz.mem_471_sv2v_reg ;
  assign \nz.mem [470] = \nz.mem_470_sv2v_reg ;
  assign \nz.mem [469] = \nz.mem_469_sv2v_reg ;
  assign \nz.mem [468] = \nz.mem_468_sv2v_reg ;
  assign \nz.mem [467] = \nz.mem_467_sv2v_reg ;
  assign \nz.mem [466] = \nz.mem_466_sv2v_reg ;
  assign \nz.mem [465] = \nz.mem_465_sv2v_reg ;
  assign \nz.mem [464] = \nz.mem_464_sv2v_reg ;
  assign \nz.mem [463] = \nz.mem_463_sv2v_reg ;
  assign \nz.mem [462] = \nz.mem_462_sv2v_reg ;
  assign \nz.mem [461] = \nz.mem_461_sv2v_reg ;
  assign \nz.mem [460] = \nz.mem_460_sv2v_reg ;
  assign \nz.mem [459] = \nz.mem_459_sv2v_reg ;
  assign \nz.mem [458] = \nz.mem_458_sv2v_reg ;
  assign \nz.mem [457] = \nz.mem_457_sv2v_reg ;
  assign \nz.mem [456] = \nz.mem_456_sv2v_reg ;
  assign \nz.mem [455] = \nz.mem_455_sv2v_reg ;
  assign \nz.mem [454] = \nz.mem_454_sv2v_reg ;
  assign \nz.mem [453] = \nz.mem_453_sv2v_reg ;
  assign \nz.mem [452] = \nz.mem_452_sv2v_reg ;
  assign \nz.mem [451] = \nz.mem_451_sv2v_reg ;
  assign \nz.mem [450] = \nz.mem_450_sv2v_reg ;
  assign \nz.mem [449] = \nz.mem_449_sv2v_reg ;
  assign \nz.mem [448] = \nz.mem_448_sv2v_reg ;
  assign \nz.mem [447] = \nz.mem_447_sv2v_reg ;
  assign \nz.mem [446] = \nz.mem_446_sv2v_reg ;
  assign \nz.mem [445] = \nz.mem_445_sv2v_reg ;
  assign \nz.mem [444] = \nz.mem_444_sv2v_reg ;
  assign \nz.mem [443] = \nz.mem_443_sv2v_reg ;
  assign \nz.mem [442] = \nz.mem_442_sv2v_reg ;
  assign \nz.mem [441] = \nz.mem_441_sv2v_reg ;
  assign \nz.mem [440] = \nz.mem_440_sv2v_reg ;
  assign \nz.mem [439] = \nz.mem_439_sv2v_reg ;
  assign \nz.mem [438] = \nz.mem_438_sv2v_reg ;
  assign \nz.mem [437] = \nz.mem_437_sv2v_reg ;
  assign \nz.mem [436] = \nz.mem_436_sv2v_reg ;
  assign \nz.mem [435] = \nz.mem_435_sv2v_reg ;
  assign \nz.mem [434] = \nz.mem_434_sv2v_reg ;
  assign \nz.mem [433] = \nz.mem_433_sv2v_reg ;
  assign \nz.mem [432] = \nz.mem_432_sv2v_reg ;
  assign \nz.mem [431] = \nz.mem_431_sv2v_reg ;
  assign \nz.mem [430] = \nz.mem_430_sv2v_reg ;
  assign \nz.mem [429] = \nz.mem_429_sv2v_reg ;
  assign \nz.mem [428] = \nz.mem_428_sv2v_reg ;
  assign \nz.mem [427] = \nz.mem_427_sv2v_reg ;
  assign \nz.mem [426] = \nz.mem_426_sv2v_reg ;
  assign \nz.mem [425] = \nz.mem_425_sv2v_reg ;
  assign \nz.mem [424] = \nz.mem_424_sv2v_reg ;
  assign \nz.mem [423] = \nz.mem_423_sv2v_reg ;
  assign \nz.mem [422] = \nz.mem_422_sv2v_reg ;
  assign \nz.mem [421] = \nz.mem_421_sv2v_reg ;
  assign \nz.mem [420] = \nz.mem_420_sv2v_reg ;
  assign \nz.mem [419] = \nz.mem_419_sv2v_reg ;
  assign \nz.mem [418] = \nz.mem_418_sv2v_reg ;
  assign \nz.mem [417] = \nz.mem_417_sv2v_reg ;
  assign \nz.mem [416] = \nz.mem_416_sv2v_reg ;
  assign \nz.mem [415] = \nz.mem_415_sv2v_reg ;
  assign \nz.mem [414] = \nz.mem_414_sv2v_reg ;
  assign \nz.mem [413] = \nz.mem_413_sv2v_reg ;
  assign \nz.mem [412] = \nz.mem_412_sv2v_reg ;
  assign \nz.mem [411] = \nz.mem_411_sv2v_reg ;
  assign \nz.mem [410] = \nz.mem_410_sv2v_reg ;
  assign \nz.mem [409] = \nz.mem_409_sv2v_reg ;
  assign \nz.mem [408] = \nz.mem_408_sv2v_reg ;
  assign \nz.mem [407] = \nz.mem_407_sv2v_reg ;
  assign \nz.mem [406] = \nz.mem_406_sv2v_reg ;
  assign \nz.mem [405] = \nz.mem_405_sv2v_reg ;
  assign \nz.mem [404] = \nz.mem_404_sv2v_reg ;
  assign \nz.mem [403] = \nz.mem_403_sv2v_reg ;
  assign \nz.mem [402] = \nz.mem_402_sv2v_reg ;
  assign \nz.mem [401] = \nz.mem_401_sv2v_reg ;
  assign \nz.mem [400] = \nz.mem_400_sv2v_reg ;
  assign \nz.mem [399] = \nz.mem_399_sv2v_reg ;
  assign \nz.mem [398] = \nz.mem_398_sv2v_reg ;
  assign \nz.mem [397] = \nz.mem_397_sv2v_reg ;
  assign \nz.mem [396] = \nz.mem_396_sv2v_reg ;
  assign \nz.mem [395] = \nz.mem_395_sv2v_reg ;
  assign \nz.mem [394] = \nz.mem_394_sv2v_reg ;
  assign \nz.mem [393] = \nz.mem_393_sv2v_reg ;
  assign \nz.mem [392] = \nz.mem_392_sv2v_reg ;
  assign \nz.mem [391] = \nz.mem_391_sv2v_reg ;
  assign \nz.mem [390] = \nz.mem_390_sv2v_reg ;
  assign \nz.mem [389] = \nz.mem_389_sv2v_reg ;
  assign \nz.mem [388] = \nz.mem_388_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[79] = (N17)? \nz.mem [79] : 
                        (N19)? \nz.mem [159] : 
                        (N21)? \nz.mem [239] : 
                        (N23)? \nz.mem [319] : 
                        (N18)? \nz.mem [399] : 
                        (N20)? \nz.mem [479] : 
                        (N22)? \nz.mem [559] : 
                        (N24)? \nz.mem [639] : 1'b0;
  assign r_data_o[78] = (N17)? \nz.mem [78] : 
                        (N19)? \nz.mem [158] : 
                        (N21)? \nz.mem [238] : 
                        (N23)? \nz.mem [318] : 
                        (N18)? \nz.mem [398] : 
                        (N20)? \nz.mem [478] : 
                        (N22)? \nz.mem [558] : 
                        (N24)? \nz.mem [638] : 1'b0;
  assign r_data_o[77] = (N17)? \nz.mem [77] : 
                        (N19)? \nz.mem [157] : 
                        (N21)? \nz.mem [237] : 
                        (N23)? \nz.mem [317] : 
                        (N18)? \nz.mem [397] : 
                        (N20)? \nz.mem [477] : 
                        (N22)? \nz.mem [557] : 
                        (N24)? \nz.mem [637] : 1'b0;
  assign r_data_o[76] = (N17)? \nz.mem [76] : 
                        (N19)? \nz.mem [156] : 
                        (N21)? \nz.mem [236] : 
                        (N23)? \nz.mem [316] : 
                        (N18)? \nz.mem [396] : 
                        (N20)? \nz.mem [476] : 
                        (N22)? \nz.mem [556] : 
                        (N24)? \nz.mem [636] : 1'b0;
  assign r_data_o[75] = (N17)? \nz.mem [75] : 
                        (N19)? \nz.mem [155] : 
                        (N21)? \nz.mem [235] : 
                        (N23)? \nz.mem [315] : 
                        (N18)? \nz.mem [395] : 
                        (N20)? \nz.mem [475] : 
                        (N22)? \nz.mem [555] : 
                        (N24)? \nz.mem [635] : 1'b0;
  assign r_data_o[74] = (N17)? \nz.mem [74] : 
                        (N19)? \nz.mem [154] : 
                        (N21)? \nz.mem [234] : 
                        (N23)? \nz.mem [314] : 
                        (N18)? \nz.mem [394] : 
                        (N20)? \nz.mem [474] : 
                        (N22)? \nz.mem [554] : 
                        (N24)? \nz.mem [634] : 1'b0;
  assign r_data_o[73] = (N17)? \nz.mem [73] : 
                        (N19)? \nz.mem [153] : 
                        (N21)? \nz.mem [233] : 
                        (N23)? \nz.mem [313] : 
                        (N18)? \nz.mem [393] : 
                        (N20)? \nz.mem [473] : 
                        (N22)? \nz.mem [553] : 
                        (N24)? \nz.mem [633] : 1'b0;
  assign r_data_o[72] = (N17)? \nz.mem [72] : 
                        (N19)? \nz.mem [152] : 
                        (N21)? \nz.mem [232] : 
                        (N23)? \nz.mem [312] : 
                        (N18)? \nz.mem [392] : 
                        (N20)? \nz.mem [472] : 
                        (N22)? \nz.mem [552] : 
                        (N24)? \nz.mem [632] : 1'b0;
  assign r_data_o[71] = (N17)? \nz.mem [71] : 
                        (N19)? \nz.mem [151] : 
                        (N21)? \nz.mem [231] : 
                        (N23)? \nz.mem [311] : 
                        (N18)? \nz.mem [391] : 
                        (N20)? \nz.mem [471] : 
                        (N22)? \nz.mem [551] : 
                        (N24)? \nz.mem [631] : 1'b0;
  assign r_data_o[70] = (N17)? \nz.mem [70] : 
                        (N19)? \nz.mem [150] : 
                        (N21)? \nz.mem [230] : 
                        (N23)? \nz.mem [310] : 
                        (N18)? \nz.mem [390] : 
                        (N20)? \nz.mem [470] : 
                        (N22)? \nz.mem [550] : 
                        (N24)? \nz.mem [630] : 1'b0;
  assign r_data_o[69] = (N17)? \nz.mem [69] : 
                        (N19)? \nz.mem [149] : 
                        (N21)? \nz.mem [229] : 
                        (N23)? \nz.mem [309] : 
                        (N18)? \nz.mem [389] : 
                        (N20)? \nz.mem [469] : 
                        (N22)? \nz.mem [549] : 
                        (N24)? \nz.mem [629] : 1'b0;
  assign r_data_o[68] = (N17)? \nz.mem [68] : 
                        (N19)? \nz.mem [148] : 
                        (N21)? \nz.mem [228] : 
                        (N23)? \nz.mem [308] : 
                        (N18)? \nz.mem [388] : 
                        (N20)? \nz.mem [468] : 
                        (N22)? \nz.mem [548] : 
                        (N24)? \nz.mem [628] : 1'b0;
  assign r_data_o[67] = (N17)? \nz.mem [67] : 
                        (N19)? \nz.mem [147] : 
                        (N21)? \nz.mem [227] : 
                        (N23)? \nz.mem [307] : 
                        (N18)? \nz.mem [387] : 
                        (N20)? \nz.mem [467] : 
                        (N22)? \nz.mem [547] : 
                        (N24)? \nz.mem [627] : 1'b0;
  assign r_data_o[66] = (N17)? \nz.mem [66] : 
                        (N19)? \nz.mem [146] : 
                        (N21)? \nz.mem [226] : 
                        (N23)? \nz.mem [306] : 
                        (N18)? \nz.mem [386] : 
                        (N20)? \nz.mem [466] : 
                        (N22)? \nz.mem [546] : 
                        (N24)? \nz.mem [626] : 1'b0;
  assign r_data_o[65] = (N17)? \nz.mem [65] : 
                        (N19)? \nz.mem [145] : 
                        (N21)? \nz.mem [225] : 
                        (N23)? \nz.mem [305] : 
                        (N18)? \nz.mem [385] : 
                        (N20)? \nz.mem [465] : 
                        (N22)? \nz.mem [545] : 
                        (N24)? \nz.mem [625] : 1'b0;
  assign r_data_o[64] = (N17)? \nz.mem [64] : 
                        (N19)? \nz.mem [144] : 
                        (N21)? \nz.mem [224] : 
                        (N23)? \nz.mem [304] : 
                        (N18)? \nz.mem [384] : 
                        (N20)? \nz.mem [464] : 
                        (N22)? \nz.mem [544] : 
                        (N24)? \nz.mem [624] : 1'b0;
  assign r_data_o[63] = (N17)? \nz.mem [63] : 
                        (N19)? \nz.mem [143] : 
                        (N21)? \nz.mem [223] : 
                        (N23)? \nz.mem [303] : 
                        (N18)? \nz.mem [383] : 
                        (N20)? \nz.mem [463] : 
                        (N22)? \nz.mem [543] : 
                        (N24)? \nz.mem [623] : 1'b0;
  assign r_data_o[62] = (N17)? \nz.mem [62] : 
                        (N19)? \nz.mem [142] : 
                        (N21)? \nz.mem [222] : 
                        (N23)? \nz.mem [302] : 
                        (N18)? \nz.mem [382] : 
                        (N20)? \nz.mem [462] : 
                        (N22)? \nz.mem [542] : 
                        (N24)? \nz.mem [622] : 1'b0;
  assign r_data_o[61] = (N17)? \nz.mem [61] : 
                        (N19)? \nz.mem [141] : 
                        (N21)? \nz.mem [221] : 
                        (N23)? \nz.mem [301] : 
                        (N18)? \nz.mem [381] : 
                        (N20)? \nz.mem [461] : 
                        (N22)? \nz.mem [541] : 
                        (N24)? \nz.mem [621] : 1'b0;
  assign r_data_o[60] = (N17)? \nz.mem [60] : 
                        (N19)? \nz.mem [140] : 
                        (N21)? \nz.mem [220] : 
                        (N23)? \nz.mem [300] : 
                        (N18)? \nz.mem [380] : 
                        (N20)? \nz.mem [460] : 
                        (N22)? \nz.mem [540] : 
                        (N24)? \nz.mem [620] : 1'b0;
  assign r_data_o[59] = (N17)? \nz.mem [59] : 
                        (N19)? \nz.mem [139] : 
                        (N21)? \nz.mem [219] : 
                        (N23)? \nz.mem [299] : 
                        (N18)? \nz.mem [379] : 
                        (N20)? \nz.mem [459] : 
                        (N22)? \nz.mem [539] : 
                        (N24)? \nz.mem [619] : 1'b0;
  assign r_data_o[58] = (N17)? \nz.mem [58] : 
                        (N19)? \nz.mem [138] : 
                        (N21)? \nz.mem [218] : 
                        (N23)? \nz.mem [298] : 
                        (N18)? \nz.mem [378] : 
                        (N20)? \nz.mem [458] : 
                        (N22)? \nz.mem [538] : 
                        (N24)? \nz.mem [618] : 1'b0;
  assign r_data_o[57] = (N17)? \nz.mem [57] : 
                        (N19)? \nz.mem [137] : 
                        (N21)? \nz.mem [217] : 
                        (N23)? \nz.mem [297] : 
                        (N18)? \nz.mem [377] : 
                        (N20)? \nz.mem [457] : 
                        (N22)? \nz.mem [537] : 
                        (N24)? \nz.mem [617] : 1'b0;
  assign r_data_o[56] = (N17)? \nz.mem [56] : 
                        (N19)? \nz.mem [136] : 
                        (N21)? \nz.mem [216] : 
                        (N23)? \nz.mem [296] : 
                        (N18)? \nz.mem [376] : 
                        (N20)? \nz.mem [456] : 
                        (N22)? \nz.mem [536] : 
                        (N24)? \nz.mem [616] : 1'b0;
  assign r_data_o[55] = (N17)? \nz.mem [55] : 
                        (N19)? \nz.mem [135] : 
                        (N21)? \nz.mem [215] : 
                        (N23)? \nz.mem [295] : 
                        (N18)? \nz.mem [375] : 
                        (N20)? \nz.mem [455] : 
                        (N22)? \nz.mem [535] : 
                        (N24)? \nz.mem [615] : 1'b0;
  assign r_data_o[54] = (N17)? \nz.mem [54] : 
                        (N19)? \nz.mem [134] : 
                        (N21)? \nz.mem [214] : 
                        (N23)? \nz.mem [294] : 
                        (N18)? \nz.mem [374] : 
                        (N20)? \nz.mem [454] : 
                        (N22)? \nz.mem [534] : 
                        (N24)? \nz.mem [614] : 1'b0;
  assign r_data_o[53] = (N17)? \nz.mem [53] : 
                        (N19)? \nz.mem [133] : 
                        (N21)? \nz.mem [213] : 
                        (N23)? \nz.mem [293] : 
                        (N18)? \nz.mem [373] : 
                        (N20)? \nz.mem [453] : 
                        (N22)? \nz.mem [533] : 
                        (N24)? \nz.mem [613] : 1'b0;
  assign r_data_o[52] = (N17)? \nz.mem [52] : 
                        (N19)? \nz.mem [132] : 
                        (N21)? \nz.mem [212] : 
                        (N23)? \nz.mem [292] : 
                        (N18)? \nz.mem [372] : 
                        (N20)? \nz.mem [452] : 
                        (N22)? \nz.mem [532] : 
                        (N24)? \nz.mem [612] : 1'b0;
  assign r_data_o[51] = (N17)? \nz.mem [51] : 
                        (N19)? \nz.mem [131] : 
                        (N21)? \nz.mem [211] : 
                        (N23)? \nz.mem [291] : 
                        (N18)? \nz.mem [371] : 
                        (N20)? \nz.mem [451] : 
                        (N22)? \nz.mem [531] : 
                        (N24)? \nz.mem [611] : 1'b0;
  assign r_data_o[50] = (N17)? \nz.mem [50] : 
                        (N19)? \nz.mem [130] : 
                        (N21)? \nz.mem [210] : 
                        (N23)? \nz.mem [290] : 
                        (N18)? \nz.mem [370] : 
                        (N20)? \nz.mem [450] : 
                        (N22)? \nz.mem [530] : 
                        (N24)? \nz.mem [610] : 1'b0;
  assign r_data_o[49] = (N17)? \nz.mem [49] : 
                        (N19)? \nz.mem [129] : 
                        (N21)? \nz.mem [209] : 
                        (N23)? \nz.mem [289] : 
                        (N18)? \nz.mem [369] : 
                        (N20)? \nz.mem [449] : 
                        (N22)? \nz.mem [529] : 
                        (N24)? \nz.mem [609] : 1'b0;
  assign r_data_o[48] = (N17)? \nz.mem [48] : 
                        (N19)? \nz.mem [128] : 
                        (N21)? \nz.mem [208] : 
                        (N23)? \nz.mem [288] : 
                        (N18)? \nz.mem [368] : 
                        (N20)? \nz.mem [448] : 
                        (N22)? \nz.mem [528] : 
                        (N24)? \nz.mem [608] : 1'b0;
  assign r_data_o[47] = (N17)? \nz.mem [47] : 
                        (N19)? \nz.mem [127] : 
                        (N21)? \nz.mem [207] : 
                        (N23)? \nz.mem [287] : 
                        (N18)? \nz.mem [367] : 
                        (N20)? \nz.mem [447] : 
                        (N22)? \nz.mem [527] : 
                        (N24)? \nz.mem [607] : 1'b0;
  assign r_data_o[46] = (N17)? \nz.mem [46] : 
                        (N19)? \nz.mem [126] : 
                        (N21)? \nz.mem [206] : 
                        (N23)? \nz.mem [286] : 
                        (N18)? \nz.mem [366] : 
                        (N20)? \nz.mem [446] : 
                        (N22)? \nz.mem [526] : 
                        (N24)? \nz.mem [606] : 1'b0;
  assign r_data_o[45] = (N17)? \nz.mem [45] : 
                        (N19)? \nz.mem [125] : 
                        (N21)? \nz.mem [205] : 
                        (N23)? \nz.mem [285] : 
                        (N18)? \nz.mem [365] : 
                        (N20)? \nz.mem [445] : 
                        (N22)? \nz.mem [525] : 
                        (N24)? \nz.mem [605] : 1'b0;
  assign r_data_o[44] = (N17)? \nz.mem [44] : 
                        (N19)? \nz.mem [124] : 
                        (N21)? \nz.mem [204] : 
                        (N23)? \nz.mem [284] : 
                        (N18)? \nz.mem [364] : 
                        (N20)? \nz.mem [444] : 
                        (N22)? \nz.mem [524] : 
                        (N24)? \nz.mem [604] : 1'b0;
  assign r_data_o[43] = (N17)? \nz.mem [43] : 
                        (N19)? \nz.mem [123] : 
                        (N21)? \nz.mem [203] : 
                        (N23)? \nz.mem [283] : 
                        (N18)? \nz.mem [363] : 
                        (N20)? \nz.mem [443] : 
                        (N22)? \nz.mem [523] : 
                        (N24)? \nz.mem [603] : 1'b0;
  assign r_data_o[42] = (N17)? \nz.mem [42] : 
                        (N19)? \nz.mem [122] : 
                        (N21)? \nz.mem [202] : 
                        (N23)? \nz.mem [282] : 
                        (N18)? \nz.mem [362] : 
                        (N20)? \nz.mem [442] : 
                        (N22)? \nz.mem [522] : 
                        (N24)? \nz.mem [602] : 1'b0;
  assign r_data_o[41] = (N17)? \nz.mem [41] : 
                        (N19)? \nz.mem [121] : 
                        (N21)? \nz.mem [201] : 
                        (N23)? \nz.mem [281] : 
                        (N18)? \nz.mem [361] : 
                        (N20)? \nz.mem [441] : 
                        (N22)? \nz.mem [521] : 
                        (N24)? \nz.mem [601] : 1'b0;
  assign r_data_o[40] = (N17)? \nz.mem [40] : 
                        (N19)? \nz.mem [120] : 
                        (N21)? \nz.mem [200] : 
                        (N23)? \nz.mem [280] : 
                        (N18)? \nz.mem [360] : 
                        (N20)? \nz.mem [440] : 
                        (N22)? \nz.mem [520] : 
                        (N24)? \nz.mem [600] : 1'b0;
  assign r_data_o[39] = (N17)? \nz.mem [39] : 
                        (N19)? \nz.mem [119] : 
                        (N21)? \nz.mem [199] : 
                        (N23)? \nz.mem [279] : 
                        (N18)? \nz.mem [359] : 
                        (N20)? \nz.mem [439] : 
                        (N22)? \nz.mem [519] : 
                        (N24)? \nz.mem [599] : 1'b0;
  assign r_data_o[38] = (N17)? \nz.mem [38] : 
                        (N19)? \nz.mem [118] : 
                        (N21)? \nz.mem [198] : 
                        (N23)? \nz.mem [278] : 
                        (N18)? \nz.mem [358] : 
                        (N20)? \nz.mem [438] : 
                        (N22)? \nz.mem [518] : 
                        (N24)? \nz.mem [598] : 1'b0;
  assign r_data_o[37] = (N17)? \nz.mem [37] : 
                        (N19)? \nz.mem [117] : 
                        (N21)? \nz.mem [197] : 
                        (N23)? \nz.mem [277] : 
                        (N18)? \nz.mem [357] : 
                        (N20)? \nz.mem [437] : 
                        (N22)? \nz.mem [517] : 
                        (N24)? \nz.mem [597] : 1'b0;
  assign r_data_o[36] = (N17)? \nz.mem [36] : 
                        (N19)? \nz.mem [116] : 
                        (N21)? \nz.mem [196] : 
                        (N23)? \nz.mem [276] : 
                        (N18)? \nz.mem [356] : 
                        (N20)? \nz.mem [436] : 
                        (N22)? \nz.mem [516] : 
                        (N24)? \nz.mem [596] : 1'b0;
  assign r_data_o[35] = (N17)? \nz.mem [35] : 
                        (N19)? \nz.mem [115] : 
                        (N21)? \nz.mem [195] : 
                        (N23)? \nz.mem [275] : 
                        (N18)? \nz.mem [355] : 
                        (N20)? \nz.mem [435] : 
                        (N22)? \nz.mem [515] : 
                        (N24)? \nz.mem [595] : 1'b0;
  assign r_data_o[34] = (N17)? \nz.mem [34] : 
                        (N19)? \nz.mem [114] : 
                        (N21)? \nz.mem [194] : 
                        (N23)? \nz.mem [274] : 
                        (N18)? \nz.mem [354] : 
                        (N20)? \nz.mem [434] : 
                        (N22)? \nz.mem [514] : 
                        (N24)? \nz.mem [594] : 1'b0;
  assign r_data_o[33] = (N17)? \nz.mem [33] : 
                        (N19)? \nz.mem [113] : 
                        (N21)? \nz.mem [193] : 
                        (N23)? \nz.mem [273] : 
                        (N18)? \nz.mem [353] : 
                        (N20)? \nz.mem [433] : 
                        (N22)? \nz.mem [513] : 
                        (N24)? \nz.mem [593] : 1'b0;
  assign r_data_o[32] = (N17)? \nz.mem [32] : 
                        (N19)? \nz.mem [112] : 
                        (N21)? \nz.mem [192] : 
                        (N23)? \nz.mem [272] : 
                        (N18)? \nz.mem [352] : 
                        (N20)? \nz.mem [432] : 
                        (N22)? \nz.mem [512] : 
                        (N24)? \nz.mem [592] : 1'b0;
  assign r_data_o[31] = (N17)? \nz.mem [31] : 
                        (N19)? \nz.mem [111] : 
                        (N21)? \nz.mem [191] : 
                        (N23)? \nz.mem [271] : 
                        (N18)? \nz.mem [351] : 
                        (N20)? \nz.mem [431] : 
                        (N22)? \nz.mem [511] : 
                        (N24)? \nz.mem [591] : 1'b0;
  assign r_data_o[30] = (N17)? \nz.mem [30] : 
                        (N19)? \nz.mem [110] : 
                        (N21)? \nz.mem [190] : 
                        (N23)? \nz.mem [270] : 
                        (N18)? \nz.mem [350] : 
                        (N20)? \nz.mem [430] : 
                        (N22)? \nz.mem [510] : 
                        (N24)? \nz.mem [590] : 1'b0;
  assign r_data_o[29] = (N17)? \nz.mem [29] : 
                        (N19)? \nz.mem [109] : 
                        (N21)? \nz.mem [189] : 
                        (N23)? \nz.mem [269] : 
                        (N18)? \nz.mem [349] : 
                        (N20)? \nz.mem [429] : 
                        (N22)? \nz.mem [509] : 
                        (N24)? \nz.mem [589] : 1'b0;
  assign r_data_o[28] = (N17)? \nz.mem [28] : 
                        (N19)? \nz.mem [108] : 
                        (N21)? \nz.mem [188] : 
                        (N23)? \nz.mem [268] : 
                        (N18)? \nz.mem [348] : 
                        (N20)? \nz.mem [428] : 
                        (N22)? \nz.mem [508] : 
                        (N24)? \nz.mem [588] : 1'b0;
  assign r_data_o[27] = (N17)? \nz.mem [27] : 
                        (N19)? \nz.mem [107] : 
                        (N21)? \nz.mem [187] : 
                        (N23)? \nz.mem [267] : 
                        (N18)? \nz.mem [347] : 
                        (N20)? \nz.mem [427] : 
                        (N22)? \nz.mem [507] : 
                        (N24)? \nz.mem [587] : 1'b0;
  assign r_data_o[26] = (N17)? \nz.mem [26] : 
                        (N19)? \nz.mem [106] : 
                        (N21)? \nz.mem [186] : 
                        (N23)? \nz.mem [266] : 
                        (N18)? \nz.mem [346] : 
                        (N20)? \nz.mem [426] : 
                        (N22)? \nz.mem [506] : 
                        (N24)? \nz.mem [586] : 1'b0;
  assign r_data_o[25] = (N17)? \nz.mem [25] : 
                        (N19)? \nz.mem [105] : 
                        (N21)? \nz.mem [185] : 
                        (N23)? \nz.mem [265] : 
                        (N18)? \nz.mem [345] : 
                        (N20)? \nz.mem [425] : 
                        (N22)? \nz.mem [505] : 
                        (N24)? \nz.mem [585] : 1'b0;
  assign r_data_o[24] = (N17)? \nz.mem [24] : 
                        (N19)? \nz.mem [104] : 
                        (N21)? \nz.mem [184] : 
                        (N23)? \nz.mem [264] : 
                        (N18)? \nz.mem [344] : 
                        (N20)? \nz.mem [424] : 
                        (N22)? \nz.mem [504] : 
                        (N24)? \nz.mem [584] : 1'b0;
  assign r_data_o[23] = (N17)? \nz.mem [23] : 
                        (N19)? \nz.mem [103] : 
                        (N21)? \nz.mem [183] : 
                        (N23)? \nz.mem [263] : 
                        (N18)? \nz.mem [343] : 
                        (N20)? \nz.mem [423] : 
                        (N22)? \nz.mem [503] : 
                        (N24)? \nz.mem [583] : 1'b0;
  assign r_data_o[22] = (N17)? \nz.mem [22] : 
                        (N19)? \nz.mem [102] : 
                        (N21)? \nz.mem [182] : 
                        (N23)? \nz.mem [262] : 
                        (N18)? \nz.mem [342] : 
                        (N20)? \nz.mem [422] : 
                        (N22)? \nz.mem [502] : 
                        (N24)? \nz.mem [582] : 1'b0;
  assign r_data_o[21] = (N17)? \nz.mem [21] : 
                        (N19)? \nz.mem [101] : 
                        (N21)? \nz.mem [181] : 
                        (N23)? \nz.mem [261] : 
                        (N18)? \nz.mem [341] : 
                        (N20)? \nz.mem [421] : 
                        (N22)? \nz.mem [501] : 
                        (N24)? \nz.mem [581] : 1'b0;
  assign r_data_o[20] = (N17)? \nz.mem [20] : 
                        (N19)? \nz.mem [100] : 
                        (N21)? \nz.mem [180] : 
                        (N23)? \nz.mem [260] : 
                        (N18)? \nz.mem [340] : 
                        (N20)? \nz.mem [420] : 
                        (N22)? \nz.mem [500] : 
                        (N24)? \nz.mem [580] : 1'b0;
  assign r_data_o[19] = (N17)? \nz.mem [19] : 
                        (N19)? \nz.mem [99] : 
                        (N21)? \nz.mem [179] : 
                        (N23)? \nz.mem [259] : 
                        (N18)? \nz.mem [339] : 
                        (N20)? \nz.mem [419] : 
                        (N22)? \nz.mem [499] : 
                        (N24)? \nz.mem [579] : 1'b0;
  assign r_data_o[18] = (N17)? \nz.mem [18] : 
                        (N19)? \nz.mem [98] : 
                        (N21)? \nz.mem [178] : 
                        (N23)? \nz.mem [258] : 
                        (N18)? \nz.mem [338] : 
                        (N20)? \nz.mem [418] : 
                        (N22)? \nz.mem [498] : 
                        (N24)? \nz.mem [578] : 1'b0;
  assign r_data_o[17] = (N17)? \nz.mem [17] : 
                        (N19)? \nz.mem [97] : 
                        (N21)? \nz.mem [177] : 
                        (N23)? \nz.mem [257] : 
                        (N18)? \nz.mem [337] : 
                        (N20)? \nz.mem [417] : 
                        (N22)? \nz.mem [497] : 
                        (N24)? \nz.mem [577] : 1'b0;
  assign r_data_o[16] = (N17)? \nz.mem [16] : 
                        (N19)? \nz.mem [96] : 
                        (N21)? \nz.mem [176] : 
                        (N23)? \nz.mem [256] : 
                        (N18)? \nz.mem [336] : 
                        (N20)? \nz.mem [416] : 
                        (N22)? \nz.mem [496] : 
                        (N24)? \nz.mem [576] : 1'b0;
  assign r_data_o[15] = (N17)? \nz.mem [15] : 
                        (N19)? \nz.mem [95] : 
                        (N21)? \nz.mem [175] : 
                        (N23)? \nz.mem [255] : 
                        (N18)? \nz.mem [335] : 
                        (N20)? \nz.mem [415] : 
                        (N22)? \nz.mem [495] : 
                        (N24)? \nz.mem [575] : 1'b0;
  assign r_data_o[14] = (N17)? \nz.mem [14] : 
                        (N19)? \nz.mem [94] : 
                        (N21)? \nz.mem [174] : 
                        (N23)? \nz.mem [254] : 
                        (N18)? \nz.mem [334] : 
                        (N20)? \nz.mem [414] : 
                        (N22)? \nz.mem [494] : 
                        (N24)? \nz.mem [574] : 1'b0;
  assign r_data_o[13] = (N17)? \nz.mem [13] : 
                        (N19)? \nz.mem [93] : 
                        (N21)? \nz.mem [173] : 
                        (N23)? \nz.mem [253] : 
                        (N18)? \nz.mem [333] : 
                        (N20)? \nz.mem [413] : 
                        (N22)? \nz.mem [493] : 
                        (N24)? \nz.mem [573] : 1'b0;
  assign r_data_o[12] = (N17)? \nz.mem [12] : 
                        (N19)? \nz.mem [92] : 
                        (N21)? \nz.mem [172] : 
                        (N23)? \nz.mem [252] : 
                        (N18)? \nz.mem [332] : 
                        (N20)? \nz.mem [412] : 
                        (N22)? \nz.mem [492] : 
                        (N24)? \nz.mem [572] : 1'b0;
  assign r_data_o[11] = (N17)? \nz.mem [11] : 
                        (N19)? \nz.mem [91] : 
                        (N21)? \nz.mem [171] : 
                        (N23)? \nz.mem [251] : 
                        (N18)? \nz.mem [331] : 
                        (N20)? \nz.mem [411] : 
                        (N22)? \nz.mem [491] : 
                        (N24)? \nz.mem [571] : 1'b0;
  assign r_data_o[10] = (N17)? \nz.mem [10] : 
                        (N19)? \nz.mem [90] : 
                        (N21)? \nz.mem [170] : 
                        (N23)? \nz.mem [250] : 
                        (N18)? \nz.mem [330] : 
                        (N20)? \nz.mem [410] : 
                        (N22)? \nz.mem [490] : 
                        (N24)? \nz.mem [570] : 1'b0;
  assign r_data_o[9] = (N17)? \nz.mem [9] : 
                       (N19)? \nz.mem [89] : 
                       (N21)? \nz.mem [169] : 
                       (N23)? \nz.mem [249] : 
                       (N18)? \nz.mem [329] : 
                       (N20)? \nz.mem [409] : 
                       (N22)? \nz.mem [489] : 
                       (N24)? \nz.mem [569] : 1'b0;
  assign r_data_o[8] = (N17)? \nz.mem [8] : 
                       (N19)? \nz.mem [88] : 
                       (N21)? \nz.mem [168] : 
                       (N23)? \nz.mem [248] : 
                       (N18)? \nz.mem [328] : 
                       (N20)? \nz.mem [408] : 
                       (N22)? \nz.mem [488] : 
                       (N24)? \nz.mem [568] : 1'b0;
  assign r_data_o[7] = (N17)? \nz.mem [7] : 
                       (N19)? \nz.mem [87] : 
                       (N21)? \nz.mem [167] : 
                       (N23)? \nz.mem [247] : 
                       (N18)? \nz.mem [327] : 
                       (N20)? \nz.mem [407] : 
                       (N22)? \nz.mem [487] : 
                       (N24)? \nz.mem [567] : 1'b0;
  assign r_data_o[6] = (N17)? \nz.mem [6] : 
                       (N19)? \nz.mem [86] : 
                       (N21)? \nz.mem [166] : 
                       (N23)? \nz.mem [246] : 
                       (N18)? \nz.mem [326] : 
                       (N20)? \nz.mem [406] : 
                       (N22)? \nz.mem [486] : 
                       (N24)? \nz.mem [566] : 1'b0;
  assign r_data_o[5] = (N17)? \nz.mem [5] : 
                       (N19)? \nz.mem [85] : 
                       (N21)? \nz.mem [165] : 
                       (N23)? \nz.mem [245] : 
                       (N18)? \nz.mem [325] : 
                       (N20)? \nz.mem [405] : 
                       (N22)? \nz.mem [485] : 
                       (N24)? \nz.mem [565] : 1'b0;
  assign r_data_o[4] = (N17)? \nz.mem [4] : 
                       (N19)? \nz.mem [84] : 
                       (N21)? \nz.mem [164] : 
                       (N23)? \nz.mem [244] : 
                       (N18)? \nz.mem [324] : 
                       (N20)? \nz.mem [404] : 
                       (N22)? \nz.mem [484] : 
                       (N24)? \nz.mem [564] : 1'b0;
  assign r_data_o[3] = (N17)? \nz.mem [3] : 
                       (N19)? \nz.mem [83] : 
                       (N21)? \nz.mem [163] : 
                       (N23)? \nz.mem [243] : 
                       (N18)? \nz.mem [323] : 
                       (N20)? \nz.mem [403] : 
                       (N22)? \nz.mem [483] : 
                       (N24)? \nz.mem [563] : 1'b0;
  assign r_data_o[2] = (N17)? \nz.mem [2] : 
                       (N19)? \nz.mem [82] : 
                       (N21)? \nz.mem [162] : 
                       (N23)? \nz.mem [242] : 
                       (N18)? \nz.mem [322] : 
                       (N20)? \nz.mem [402] : 
                       (N22)? \nz.mem [482] : 
                       (N24)? \nz.mem [562] : 1'b0;
  assign r_data_o[1] = (N17)? \nz.mem [1] : 
                       (N19)? \nz.mem [81] : 
                       (N21)? \nz.mem [161] : 
                       (N23)? \nz.mem [241] : 
                       (N18)? \nz.mem [321] : 
                       (N20)? \nz.mem [401] : 
                       (N22)? \nz.mem [481] : 
                       (N24)? \nz.mem [561] : 1'b0;
  assign r_data_o[0] = (N17)? \nz.mem [0] : 
                       (N19)? \nz.mem [80] : 
                       (N21)? \nz.mem [160] : 
                       (N23)? \nz.mem [240] : 
                       (N18)? \nz.mem [320] : 
                       (N20)? \nz.mem [400] : 
                       (N22)? \nz.mem [480] : 
                       (N24)? \nz.mem [560] : 1'b0;
  assign N42 = w_addr_i[0] & w_addr_i[1];
  assign N33 = N42 & w_addr_i[2];
  assign N43 = N0 & w_addr_i[1];
  assign N0 = ~w_addr_i[0];
  assign N32 = N43 & w_addr_i[2];
  assign N44 = w_addr_i[0] & N1;
  assign N1 = ~w_addr_i[1];
  assign N31 = N44 & w_addr_i[2];
  assign N45 = N2 & N3;
  assign N2 = ~w_addr_i[0];
  assign N3 = ~w_addr_i[1];
  assign N30 = N45 & w_addr_i[2];
  assign N29 = N42 & N4;
  assign N4 = ~w_addr_i[2];
  assign N28 = N43 & N5;
  assign N5 = ~w_addr_i[2];
  assign N27 = N44 & N6;
  assign N6 = ~w_addr_i[2];
  assign N26 = N45 & N7;
  assign N7 = ~w_addr_i[2];
  assign { N41, N40, N39, N38, N37, N36, N35, N34 } = (N8)? { N33, N32, N31, N30, N29, N28, N27, N26 } : 
                                                      (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N25;
  assign N10 = ~r_addr_i[0];
  assign N11 = ~r_addr_i[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r_addr_i[1];
  assign N14 = r_addr_i[0] & N11;
  assign N15 = r_addr_i[0] & r_addr_i[1];
  assign N16 = ~r_addr_i[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r_addr_i[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r_addr_i[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r_addr_i[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r_addr_i[2];
  assign N25 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N41) begin
      \nz.mem_639_sv2v_reg  <= w_data_i[79];
      \nz.mem_638_sv2v_reg  <= w_data_i[78];
      \nz.mem_637_sv2v_reg  <= w_data_i[77];
      \nz.mem_636_sv2v_reg  <= w_data_i[76];
      \nz.mem_635_sv2v_reg  <= w_data_i[75];
      \nz.mem_634_sv2v_reg  <= w_data_i[74];
      \nz.mem_633_sv2v_reg  <= w_data_i[73];
      \nz.mem_632_sv2v_reg  <= w_data_i[72];
      \nz.mem_631_sv2v_reg  <= w_data_i[71];
      \nz.mem_630_sv2v_reg  <= w_data_i[70];
      \nz.mem_629_sv2v_reg  <= w_data_i[69];
      \nz.mem_628_sv2v_reg  <= w_data_i[68];
      \nz.mem_627_sv2v_reg  <= w_data_i[67];
      \nz.mem_626_sv2v_reg  <= w_data_i[66];
      \nz.mem_625_sv2v_reg  <= w_data_i[65];
      \nz.mem_624_sv2v_reg  <= w_data_i[64];
      \nz.mem_623_sv2v_reg  <= w_data_i[63];
      \nz.mem_622_sv2v_reg  <= w_data_i[62];
      \nz.mem_621_sv2v_reg  <= w_data_i[61];
      \nz.mem_620_sv2v_reg  <= w_data_i[60];
      \nz.mem_619_sv2v_reg  <= w_data_i[59];
      \nz.mem_618_sv2v_reg  <= w_data_i[58];
      \nz.mem_617_sv2v_reg  <= w_data_i[57];
      \nz.mem_616_sv2v_reg  <= w_data_i[56];
      \nz.mem_615_sv2v_reg  <= w_data_i[55];
      \nz.mem_614_sv2v_reg  <= w_data_i[54];
      \nz.mem_613_sv2v_reg  <= w_data_i[53];
      \nz.mem_612_sv2v_reg  <= w_data_i[52];
      \nz.mem_611_sv2v_reg  <= w_data_i[51];
      \nz.mem_610_sv2v_reg  <= w_data_i[50];
      \nz.mem_609_sv2v_reg  <= w_data_i[49];
      \nz.mem_608_sv2v_reg  <= w_data_i[48];
      \nz.mem_607_sv2v_reg  <= w_data_i[47];
      \nz.mem_606_sv2v_reg  <= w_data_i[46];
      \nz.mem_605_sv2v_reg  <= w_data_i[45];
      \nz.mem_604_sv2v_reg  <= w_data_i[44];
      \nz.mem_603_sv2v_reg  <= w_data_i[43];
      \nz.mem_602_sv2v_reg  <= w_data_i[42];
      \nz.mem_601_sv2v_reg  <= w_data_i[41];
      \nz.mem_600_sv2v_reg  <= w_data_i[40];
      \nz.mem_599_sv2v_reg  <= w_data_i[39];
      \nz.mem_598_sv2v_reg  <= w_data_i[38];
      \nz.mem_597_sv2v_reg  <= w_data_i[37];
      \nz.mem_596_sv2v_reg  <= w_data_i[36];
      \nz.mem_595_sv2v_reg  <= w_data_i[35];
      \nz.mem_594_sv2v_reg  <= w_data_i[34];
      \nz.mem_593_sv2v_reg  <= w_data_i[33];
      \nz.mem_592_sv2v_reg  <= w_data_i[32];
      \nz.mem_591_sv2v_reg  <= w_data_i[31];
      \nz.mem_590_sv2v_reg  <= w_data_i[30];
      \nz.mem_589_sv2v_reg  <= w_data_i[29];
      \nz.mem_588_sv2v_reg  <= w_data_i[28];
      \nz.mem_587_sv2v_reg  <= w_data_i[27];
      \nz.mem_586_sv2v_reg  <= w_data_i[26];
      \nz.mem_585_sv2v_reg  <= w_data_i[25];
      \nz.mem_584_sv2v_reg  <= w_data_i[24];
      \nz.mem_583_sv2v_reg  <= w_data_i[23];
      \nz.mem_582_sv2v_reg  <= w_data_i[22];
      \nz.mem_581_sv2v_reg  <= w_data_i[21];
      \nz.mem_580_sv2v_reg  <= w_data_i[20];
      \nz.mem_579_sv2v_reg  <= w_data_i[19];
      \nz.mem_578_sv2v_reg  <= w_data_i[18];
      \nz.mem_577_sv2v_reg  <= w_data_i[17];
      \nz.mem_576_sv2v_reg  <= w_data_i[16];
      \nz.mem_575_sv2v_reg  <= w_data_i[15];
      \nz.mem_574_sv2v_reg  <= w_data_i[14];
      \nz.mem_573_sv2v_reg  <= w_data_i[13];
      \nz.mem_572_sv2v_reg  <= w_data_i[12];
      \nz.mem_571_sv2v_reg  <= w_data_i[11];
      \nz.mem_570_sv2v_reg  <= w_data_i[10];
      \nz.mem_569_sv2v_reg  <= w_data_i[9];
      \nz.mem_568_sv2v_reg  <= w_data_i[8];
      \nz.mem_567_sv2v_reg  <= w_data_i[7];
      \nz.mem_566_sv2v_reg  <= w_data_i[6];
      \nz.mem_565_sv2v_reg  <= w_data_i[5];
      \nz.mem_564_sv2v_reg  <= w_data_i[4];
      \nz.mem_563_sv2v_reg  <= w_data_i[3];
      \nz.mem_562_sv2v_reg  <= w_data_i[2];
      \nz.mem_561_sv2v_reg  <= w_data_i[1];
      \nz.mem_560_sv2v_reg  <= w_data_i[0];
    end 
    if(N40) begin
      \nz.mem_559_sv2v_reg  <= w_data_i[79];
      \nz.mem_558_sv2v_reg  <= w_data_i[78];
      \nz.mem_557_sv2v_reg  <= w_data_i[77];
      \nz.mem_556_sv2v_reg  <= w_data_i[76];
      \nz.mem_555_sv2v_reg  <= w_data_i[75];
      \nz.mem_554_sv2v_reg  <= w_data_i[74];
      \nz.mem_553_sv2v_reg  <= w_data_i[73];
      \nz.mem_552_sv2v_reg  <= w_data_i[72];
      \nz.mem_551_sv2v_reg  <= w_data_i[71];
      \nz.mem_550_sv2v_reg  <= w_data_i[70];
      \nz.mem_549_sv2v_reg  <= w_data_i[69];
      \nz.mem_548_sv2v_reg  <= w_data_i[68];
      \nz.mem_547_sv2v_reg  <= w_data_i[67];
      \nz.mem_546_sv2v_reg  <= w_data_i[66];
      \nz.mem_545_sv2v_reg  <= w_data_i[65];
      \nz.mem_544_sv2v_reg  <= w_data_i[64];
      \nz.mem_543_sv2v_reg  <= w_data_i[63];
      \nz.mem_542_sv2v_reg  <= w_data_i[62];
      \nz.mem_541_sv2v_reg  <= w_data_i[61];
      \nz.mem_540_sv2v_reg  <= w_data_i[60];
      \nz.mem_539_sv2v_reg  <= w_data_i[59];
      \nz.mem_538_sv2v_reg  <= w_data_i[58];
      \nz.mem_537_sv2v_reg  <= w_data_i[57];
      \nz.mem_536_sv2v_reg  <= w_data_i[56];
      \nz.mem_535_sv2v_reg  <= w_data_i[55];
      \nz.mem_534_sv2v_reg  <= w_data_i[54];
      \nz.mem_533_sv2v_reg  <= w_data_i[53];
      \nz.mem_532_sv2v_reg  <= w_data_i[52];
      \nz.mem_531_sv2v_reg  <= w_data_i[51];
      \nz.mem_530_sv2v_reg  <= w_data_i[50];
      \nz.mem_529_sv2v_reg  <= w_data_i[49];
      \nz.mem_528_sv2v_reg  <= w_data_i[48];
      \nz.mem_527_sv2v_reg  <= w_data_i[47];
      \nz.mem_526_sv2v_reg  <= w_data_i[46];
      \nz.mem_525_sv2v_reg  <= w_data_i[45];
      \nz.mem_524_sv2v_reg  <= w_data_i[44];
      \nz.mem_523_sv2v_reg  <= w_data_i[43];
      \nz.mem_522_sv2v_reg  <= w_data_i[42];
      \nz.mem_521_sv2v_reg  <= w_data_i[41];
      \nz.mem_520_sv2v_reg  <= w_data_i[40];
      \nz.mem_519_sv2v_reg  <= w_data_i[39];
      \nz.mem_518_sv2v_reg  <= w_data_i[38];
      \nz.mem_517_sv2v_reg  <= w_data_i[37];
      \nz.mem_516_sv2v_reg  <= w_data_i[36];
      \nz.mem_515_sv2v_reg  <= w_data_i[35];
      \nz.mem_514_sv2v_reg  <= w_data_i[34];
      \nz.mem_513_sv2v_reg  <= w_data_i[33];
      \nz.mem_512_sv2v_reg  <= w_data_i[32];
      \nz.mem_511_sv2v_reg  <= w_data_i[31];
      \nz.mem_510_sv2v_reg  <= w_data_i[30];
      \nz.mem_509_sv2v_reg  <= w_data_i[29];
      \nz.mem_508_sv2v_reg  <= w_data_i[28];
      \nz.mem_507_sv2v_reg  <= w_data_i[27];
      \nz.mem_506_sv2v_reg  <= w_data_i[26];
      \nz.mem_505_sv2v_reg  <= w_data_i[25];
      \nz.mem_504_sv2v_reg  <= w_data_i[24];
      \nz.mem_503_sv2v_reg  <= w_data_i[23];
      \nz.mem_502_sv2v_reg  <= w_data_i[22];
      \nz.mem_501_sv2v_reg  <= w_data_i[21];
      \nz.mem_500_sv2v_reg  <= w_data_i[20];
      \nz.mem_499_sv2v_reg  <= w_data_i[19];
      \nz.mem_498_sv2v_reg  <= w_data_i[18];
      \nz.mem_497_sv2v_reg  <= w_data_i[17];
      \nz.mem_496_sv2v_reg  <= w_data_i[16];
      \nz.mem_495_sv2v_reg  <= w_data_i[15];
      \nz.mem_494_sv2v_reg  <= w_data_i[14];
      \nz.mem_493_sv2v_reg  <= w_data_i[13];
      \nz.mem_492_sv2v_reg  <= w_data_i[12];
      \nz.mem_491_sv2v_reg  <= w_data_i[11];
      \nz.mem_490_sv2v_reg  <= w_data_i[10];
      \nz.mem_489_sv2v_reg  <= w_data_i[9];
      \nz.mem_488_sv2v_reg  <= w_data_i[8];
      \nz.mem_487_sv2v_reg  <= w_data_i[7];
      \nz.mem_486_sv2v_reg  <= w_data_i[6];
      \nz.mem_485_sv2v_reg  <= w_data_i[5];
      \nz.mem_484_sv2v_reg  <= w_data_i[4];
      \nz.mem_483_sv2v_reg  <= w_data_i[3];
      \nz.mem_482_sv2v_reg  <= w_data_i[2];
      \nz.mem_481_sv2v_reg  <= w_data_i[1];
      \nz.mem_480_sv2v_reg  <= w_data_i[0];
    end 
    if(N39) begin
      \nz.mem_479_sv2v_reg  <= w_data_i[79];
      \nz.mem_478_sv2v_reg  <= w_data_i[78];
      \nz.mem_477_sv2v_reg  <= w_data_i[77];
      \nz.mem_476_sv2v_reg  <= w_data_i[76];
      \nz.mem_475_sv2v_reg  <= w_data_i[75];
      \nz.mem_474_sv2v_reg  <= w_data_i[74];
      \nz.mem_473_sv2v_reg  <= w_data_i[73];
      \nz.mem_472_sv2v_reg  <= w_data_i[72];
      \nz.mem_471_sv2v_reg  <= w_data_i[71];
      \nz.mem_470_sv2v_reg  <= w_data_i[70];
      \nz.mem_469_sv2v_reg  <= w_data_i[69];
      \nz.mem_468_sv2v_reg  <= w_data_i[68];
      \nz.mem_467_sv2v_reg  <= w_data_i[67];
      \nz.mem_466_sv2v_reg  <= w_data_i[66];
      \nz.mem_465_sv2v_reg  <= w_data_i[65];
      \nz.mem_464_sv2v_reg  <= w_data_i[64];
      \nz.mem_463_sv2v_reg  <= w_data_i[63];
      \nz.mem_462_sv2v_reg  <= w_data_i[62];
      \nz.mem_461_sv2v_reg  <= w_data_i[61];
      \nz.mem_460_sv2v_reg  <= w_data_i[60];
      \nz.mem_459_sv2v_reg  <= w_data_i[59];
      \nz.mem_458_sv2v_reg  <= w_data_i[58];
      \nz.mem_457_sv2v_reg  <= w_data_i[57];
      \nz.mem_456_sv2v_reg  <= w_data_i[56];
      \nz.mem_455_sv2v_reg  <= w_data_i[55];
      \nz.mem_454_sv2v_reg  <= w_data_i[54];
      \nz.mem_453_sv2v_reg  <= w_data_i[53];
      \nz.mem_452_sv2v_reg  <= w_data_i[52];
      \nz.mem_451_sv2v_reg  <= w_data_i[51];
      \nz.mem_450_sv2v_reg  <= w_data_i[50];
      \nz.mem_449_sv2v_reg  <= w_data_i[49];
      \nz.mem_448_sv2v_reg  <= w_data_i[48];
      \nz.mem_447_sv2v_reg  <= w_data_i[47];
      \nz.mem_446_sv2v_reg  <= w_data_i[46];
      \nz.mem_445_sv2v_reg  <= w_data_i[45];
      \nz.mem_444_sv2v_reg  <= w_data_i[44];
      \nz.mem_443_sv2v_reg  <= w_data_i[43];
      \nz.mem_442_sv2v_reg  <= w_data_i[42];
      \nz.mem_441_sv2v_reg  <= w_data_i[41];
      \nz.mem_440_sv2v_reg  <= w_data_i[40];
      \nz.mem_439_sv2v_reg  <= w_data_i[39];
      \nz.mem_438_sv2v_reg  <= w_data_i[38];
      \nz.mem_437_sv2v_reg  <= w_data_i[37];
      \nz.mem_436_sv2v_reg  <= w_data_i[36];
      \nz.mem_435_sv2v_reg  <= w_data_i[35];
      \nz.mem_434_sv2v_reg  <= w_data_i[34];
      \nz.mem_433_sv2v_reg  <= w_data_i[33];
      \nz.mem_432_sv2v_reg  <= w_data_i[32];
      \nz.mem_431_sv2v_reg  <= w_data_i[31];
      \nz.mem_430_sv2v_reg  <= w_data_i[30];
      \nz.mem_429_sv2v_reg  <= w_data_i[29];
      \nz.mem_428_sv2v_reg  <= w_data_i[28];
      \nz.mem_427_sv2v_reg  <= w_data_i[27];
      \nz.mem_426_sv2v_reg  <= w_data_i[26];
      \nz.mem_425_sv2v_reg  <= w_data_i[25];
      \nz.mem_424_sv2v_reg  <= w_data_i[24];
      \nz.mem_423_sv2v_reg  <= w_data_i[23];
      \nz.mem_422_sv2v_reg  <= w_data_i[22];
      \nz.mem_421_sv2v_reg  <= w_data_i[21];
      \nz.mem_420_sv2v_reg  <= w_data_i[20];
      \nz.mem_419_sv2v_reg  <= w_data_i[19];
      \nz.mem_418_sv2v_reg  <= w_data_i[18];
      \nz.mem_417_sv2v_reg  <= w_data_i[17];
      \nz.mem_416_sv2v_reg  <= w_data_i[16];
      \nz.mem_415_sv2v_reg  <= w_data_i[15];
      \nz.mem_414_sv2v_reg  <= w_data_i[14];
      \nz.mem_413_sv2v_reg  <= w_data_i[13];
      \nz.mem_412_sv2v_reg  <= w_data_i[12];
      \nz.mem_411_sv2v_reg  <= w_data_i[11];
      \nz.mem_410_sv2v_reg  <= w_data_i[10];
      \nz.mem_409_sv2v_reg  <= w_data_i[9];
      \nz.mem_408_sv2v_reg  <= w_data_i[8];
      \nz.mem_407_sv2v_reg  <= w_data_i[7];
      \nz.mem_406_sv2v_reg  <= w_data_i[6];
      \nz.mem_405_sv2v_reg  <= w_data_i[5];
      \nz.mem_404_sv2v_reg  <= w_data_i[4];
      \nz.mem_403_sv2v_reg  <= w_data_i[3];
      \nz.mem_402_sv2v_reg  <= w_data_i[2];
      \nz.mem_401_sv2v_reg  <= w_data_i[1];
      \nz.mem_400_sv2v_reg  <= w_data_i[0];
    end 
    if(N38) begin
      \nz.mem_399_sv2v_reg  <= w_data_i[79];
      \nz.mem_398_sv2v_reg  <= w_data_i[78];
      \nz.mem_397_sv2v_reg  <= w_data_i[77];
      \nz.mem_396_sv2v_reg  <= w_data_i[76];
      \nz.mem_395_sv2v_reg  <= w_data_i[75];
      \nz.mem_394_sv2v_reg  <= w_data_i[74];
      \nz.mem_393_sv2v_reg  <= w_data_i[73];
      \nz.mem_392_sv2v_reg  <= w_data_i[72];
      \nz.mem_391_sv2v_reg  <= w_data_i[71];
      \nz.mem_390_sv2v_reg  <= w_data_i[70];
      \nz.mem_389_sv2v_reg  <= w_data_i[69];
      \nz.mem_388_sv2v_reg  <= w_data_i[68];
      \nz.mem_387_sv2v_reg  <= w_data_i[67];
      \nz.mem_386_sv2v_reg  <= w_data_i[66];
      \nz.mem_385_sv2v_reg  <= w_data_i[65];
      \nz.mem_384_sv2v_reg  <= w_data_i[64];
      \nz.mem_383_sv2v_reg  <= w_data_i[63];
      \nz.mem_382_sv2v_reg  <= w_data_i[62];
      \nz.mem_381_sv2v_reg  <= w_data_i[61];
      \nz.mem_380_sv2v_reg  <= w_data_i[60];
      \nz.mem_379_sv2v_reg  <= w_data_i[59];
      \nz.mem_378_sv2v_reg  <= w_data_i[58];
      \nz.mem_377_sv2v_reg  <= w_data_i[57];
      \nz.mem_376_sv2v_reg  <= w_data_i[56];
      \nz.mem_375_sv2v_reg  <= w_data_i[55];
      \nz.mem_374_sv2v_reg  <= w_data_i[54];
      \nz.mem_373_sv2v_reg  <= w_data_i[53];
      \nz.mem_372_sv2v_reg  <= w_data_i[52];
      \nz.mem_371_sv2v_reg  <= w_data_i[51];
      \nz.mem_370_sv2v_reg  <= w_data_i[50];
      \nz.mem_369_sv2v_reg  <= w_data_i[49];
      \nz.mem_368_sv2v_reg  <= w_data_i[48];
      \nz.mem_367_sv2v_reg  <= w_data_i[47];
      \nz.mem_366_sv2v_reg  <= w_data_i[46];
      \nz.mem_365_sv2v_reg  <= w_data_i[45];
      \nz.mem_364_sv2v_reg  <= w_data_i[44];
      \nz.mem_363_sv2v_reg  <= w_data_i[43];
      \nz.mem_362_sv2v_reg  <= w_data_i[42];
      \nz.mem_361_sv2v_reg  <= w_data_i[41];
      \nz.mem_360_sv2v_reg  <= w_data_i[40];
      \nz.mem_359_sv2v_reg  <= w_data_i[39];
      \nz.mem_358_sv2v_reg  <= w_data_i[38];
      \nz.mem_357_sv2v_reg  <= w_data_i[37];
      \nz.mem_356_sv2v_reg  <= w_data_i[36];
      \nz.mem_355_sv2v_reg  <= w_data_i[35];
      \nz.mem_354_sv2v_reg  <= w_data_i[34];
      \nz.mem_353_sv2v_reg  <= w_data_i[33];
      \nz.mem_352_sv2v_reg  <= w_data_i[32];
      \nz.mem_351_sv2v_reg  <= w_data_i[31];
      \nz.mem_350_sv2v_reg  <= w_data_i[30];
      \nz.mem_349_sv2v_reg  <= w_data_i[29];
      \nz.mem_348_sv2v_reg  <= w_data_i[28];
      \nz.mem_347_sv2v_reg  <= w_data_i[27];
      \nz.mem_346_sv2v_reg  <= w_data_i[26];
      \nz.mem_345_sv2v_reg  <= w_data_i[25];
      \nz.mem_344_sv2v_reg  <= w_data_i[24];
      \nz.mem_343_sv2v_reg  <= w_data_i[23];
      \nz.mem_342_sv2v_reg  <= w_data_i[22];
      \nz.mem_341_sv2v_reg  <= w_data_i[21];
      \nz.mem_340_sv2v_reg  <= w_data_i[20];
      \nz.mem_339_sv2v_reg  <= w_data_i[19];
      \nz.mem_338_sv2v_reg  <= w_data_i[18];
      \nz.mem_337_sv2v_reg  <= w_data_i[17];
      \nz.mem_336_sv2v_reg  <= w_data_i[16];
      \nz.mem_335_sv2v_reg  <= w_data_i[15];
      \nz.mem_334_sv2v_reg  <= w_data_i[14];
      \nz.mem_333_sv2v_reg  <= w_data_i[13];
      \nz.mem_332_sv2v_reg  <= w_data_i[12];
      \nz.mem_331_sv2v_reg  <= w_data_i[11];
      \nz.mem_330_sv2v_reg  <= w_data_i[10];
      \nz.mem_329_sv2v_reg  <= w_data_i[9];
      \nz.mem_328_sv2v_reg  <= w_data_i[8];
      \nz.mem_327_sv2v_reg  <= w_data_i[7];
      \nz.mem_326_sv2v_reg  <= w_data_i[6];
      \nz.mem_325_sv2v_reg  <= w_data_i[5];
      \nz.mem_324_sv2v_reg  <= w_data_i[4];
      \nz.mem_323_sv2v_reg  <= w_data_i[3];
      \nz.mem_322_sv2v_reg  <= w_data_i[2];
      \nz.mem_321_sv2v_reg  <= w_data_i[1];
      \nz.mem_320_sv2v_reg  <= w_data_i[0];
    end 
    if(N37) begin
      \nz.mem_319_sv2v_reg  <= w_data_i[79];
      \nz.mem_318_sv2v_reg  <= w_data_i[78];
      \nz.mem_317_sv2v_reg  <= w_data_i[77];
      \nz.mem_316_sv2v_reg  <= w_data_i[76];
      \nz.mem_315_sv2v_reg  <= w_data_i[75];
      \nz.mem_314_sv2v_reg  <= w_data_i[74];
      \nz.mem_313_sv2v_reg  <= w_data_i[73];
      \nz.mem_312_sv2v_reg  <= w_data_i[72];
      \nz.mem_311_sv2v_reg  <= w_data_i[71];
      \nz.mem_310_sv2v_reg  <= w_data_i[70];
      \nz.mem_309_sv2v_reg  <= w_data_i[69];
      \nz.mem_308_sv2v_reg  <= w_data_i[68];
      \nz.mem_307_sv2v_reg  <= w_data_i[67];
      \nz.mem_306_sv2v_reg  <= w_data_i[66];
      \nz.mem_305_sv2v_reg  <= w_data_i[65];
      \nz.mem_304_sv2v_reg  <= w_data_i[64];
      \nz.mem_303_sv2v_reg  <= w_data_i[63];
      \nz.mem_302_sv2v_reg  <= w_data_i[62];
      \nz.mem_301_sv2v_reg  <= w_data_i[61];
      \nz.mem_300_sv2v_reg  <= w_data_i[60];
      \nz.mem_299_sv2v_reg  <= w_data_i[59];
      \nz.mem_298_sv2v_reg  <= w_data_i[58];
      \nz.mem_297_sv2v_reg  <= w_data_i[57];
      \nz.mem_296_sv2v_reg  <= w_data_i[56];
      \nz.mem_295_sv2v_reg  <= w_data_i[55];
      \nz.mem_294_sv2v_reg  <= w_data_i[54];
      \nz.mem_293_sv2v_reg  <= w_data_i[53];
      \nz.mem_292_sv2v_reg  <= w_data_i[52];
      \nz.mem_291_sv2v_reg  <= w_data_i[51];
      \nz.mem_290_sv2v_reg  <= w_data_i[50];
      \nz.mem_289_sv2v_reg  <= w_data_i[49];
      \nz.mem_288_sv2v_reg  <= w_data_i[48];
      \nz.mem_287_sv2v_reg  <= w_data_i[47];
      \nz.mem_286_sv2v_reg  <= w_data_i[46];
      \nz.mem_285_sv2v_reg  <= w_data_i[45];
      \nz.mem_284_sv2v_reg  <= w_data_i[44];
      \nz.mem_283_sv2v_reg  <= w_data_i[43];
      \nz.mem_282_sv2v_reg  <= w_data_i[42];
      \nz.mem_281_sv2v_reg  <= w_data_i[41];
      \nz.mem_280_sv2v_reg  <= w_data_i[40];
      \nz.mem_279_sv2v_reg  <= w_data_i[39];
      \nz.mem_278_sv2v_reg  <= w_data_i[38];
      \nz.mem_277_sv2v_reg  <= w_data_i[37];
      \nz.mem_276_sv2v_reg  <= w_data_i[36];
      \nz.mem_275_sv2v_reg  <= w_data_i[35];
      \nz.mem_274_sv2v_reg  <= w_data_i[34];
      \nz.mem_273_sv2v_reg  <= w_data_i[33];
      \nz.mem_272_sv2v_reg  <= w_data_i[32];
      \nz.mem_271_sv2v_reg  <= w_data_i[31];
      \nz.mem_270_sv2v_reg  <= w_data_i[30];
      \nz.mem_269_sv2v_reg  <= w_data_i[29];
      \nz.mem_268_sv2v_reg  <= w_data_i[28];
      \nz.mem_267_sv2v_reg  <= w_data_i[27];
      \nz.mem_266_sv2v_reg  <= w_data_i[26];
      \nz.mem_265_sv2v_reg  <= w_data_i[25];
      \nz.mem_264_sv2v_reg  <= w_data_i[24];
      \nz.mem_263_sv2v_reg  <= w_data_i[23];
      \nz.mem_262_sv2v_reg  <= w_data_i[22];
      \nz.mem_261_sv2v_reg  <= w_data_i[21];
      \nz.mem_260_sv2v_reg  <= w_data_i[20];
      \nz.mem_259_sv2v_reg  <= w_data_i[19];
      \nz.mem_258_sv2v_reg  <= w_data_i[18];
      \nz.mem_257_sv2v_reg  <= w_data_i[17];
      \nz.mem_256_sv2v_reg  <= w_data_i[16];
      \nz.mem_255_sv2v_reg  <= w_data_i[15];
      \nz.mem_254_sv2v_reg  <= w_data_i[14];
      \nz.mem_253_sv2v_reg  <= w_data_i[13];
      \nz.mem_252_sv2v_reg  <= w_data_i[12];
      \nz.mem_251_sv2v_reg  <= w_data_i[11];
      \nz.mem_250_sv2v_reg  <= w_data_i[10];
      \nz.mem_249_sv2v_reg  <= w_data_i[9];
      \nz.mem_248_sv2v_reg  <= w_data_i[8];
      \nz.mem_247_sv2v_reg  <= w_data_i[7];
      \nz.mem_246_sv2v_reg  <= w_data_i[6];
      \nz.mem_245_sv2v_reg  <= w_data_i[5];
      \nz.mem_244_sv2v_reg  <= w_data_i[4];
      \nz.mem_243_sv2v_reg  <= w_data_i[3];
      \nz.mem_242_sv2v_reg  <= w_data_i[2];
      \nz.mem_241_sv2v_reg  <= w_data_i[1];
      \nz.mem_240_sv2v_reg  <= w_data_i[0];
    end 
    if(N36) begin
      \nz.mem_239_sv2v_reg  <= w_data_i[79];
      \nz.mem_238_sv2v_reg  <= w_data_i[78];
      \nz.mem_237_sv2v_reg  <= w_data_i[77];
      \nz.mem_236_sv2v_reg  <= w_data_i[76];
      \nz.mem_235_sv2v_reg  <= w_data_i[75];
      \nz.mem_234_sv2v_reg  <= w_data_i[74];
      \nz.mem_233_sv2v_reg  <= w_data_i[73];
      \nz.mem_232_sv2v_reg  <= w_data_i[72];
      \nz.mem_231_sv2v_reg  <= w_data_i[71];
      \nz.mem_230_sv2v_reg  <= w_data_i[70];
      \nz.mem_229_sv2v_reg  <= w_data_i[69];
      \nz.mem_228_sv2v_reg  <= w_data_i[68];
      \nz.mem_227_sv2v_reg  <= w_data_i[67];
      \nz.mem_226_sv2v_reg  <= w_data_i[66];
      \nz.mem_225_sv2v_reg  <= w_data_i[65];
      \nz.mem_224_sv2v_reg  <= w_data_i[64];
      \nz.mem_223_sv2v_reg  <= w_data_i[63];
      \nz.mem_222_sv2v_reg  <= w_data_i[62];
      \nz.mem_221_sv2v_reg  <= w_data_i[61];
      \nz.mem_220_sv2v_reg  <= w_data_i[60];
      \nz.mem_219_sv2v_reg  <= w_data_i[59];
      \nz.mem_218_sv2v_reg  <= w_data_i[58];
      \nz.mem_217_sv2v_reg  <= w_data_i[57];
      \nz.mem_216_sv2v_reg  <= w_data_i[56];
      \nz.mem_215_sv2v_reg  <= w_data_i[55];
      \nz.mem_214_sv2v_reg  <= w_data_i[54];
      \nz.mem_213_sv2v_reg  <= w_data_i[53];
      \nz.mem_212_sv2v_reg  <= w_data_i[52];
      \nz.mem_211_sv2v_reg  <= w_data_i[51];
      \nz.mem_210_sv2v_reg  <= w_data_i[50];
      \nz.mem_209_sv2v_reg  <= w_data_i[49];
      \nz.mem_208_sv2v_reg  <= w_data_i[48];
      \nz.mem_207_sv2v_reg  <= w_data_i[47];
      \nz.mem_206_sv2v_reg  <= w_data_i[46];
      \nz.mem_205_sv2v_reg  <= w_data_i[45];
      \nz.mem_204_sv2v_reg  <= w_data_i[44];
      \nz.mem_203_sv2v_reg  <= w_data_i[43];
      \nz.mem_202_sv2v_reg  <= w_data_i[42];
      \nz.mem_201_sv2v_reg  <= w_data_i[41];
      \nz.mem_200_sv2v_reg  <= w_data_i[40];
      \nz.mem_199_sv2v_reg  <= w_data_i[39];
      \nz.mem_198_sv2v_reg  <= w_data_i[38];
      \nz.mem_197_sv2v_reg  <= w_data_i[37];
      \nz.mem_196_sv2v_reg  <= w_data_i[36];
      \nz.mem_195_sv2v_reg  <= w_data_i[35];
      \nz.mem_194_sv2v_reg  <= w_data_i[34];
      \nz.mem_193_sv2v_reg  <= w_data_i[33];
      \nz.mem_192_sv2v_reg  <= w_data_i[32];
      \nz.mem_191_sv2v_reg  <= w_data_i[31];
      \nz.mem_190_sv2v_reg  <= w_data_i[30];
      \nz.mem_189_sv2v_reg  <= w_data_i[29];
      \nz.mem_188_sv2v_reg  <= w_data_i[28];
      \nz.mem_187_sv2v_reg  <= w_data_i[27];
      \nz.mem_186_sv2v_reg  <= w_data_i[26];
      \nz.mem_185_sv2v_reg  <= w_data_i[25];
      \nz.mem_184_sv2v_reg  <= w_data_i[24];
      \nz.mem_183_sv2v_reg  <= w_data_i[23];
      \nz.mem_182_sv2v_reg  <= w_data_i[22];
      \nz.mem_181_sv2v_reg  <= w_data_i[21];
      \nz.mem_180_sv2v_reg  <= w_data_i[20];
      \nz.mem_179_sv2v_reg  <= w_data_i[19];
      \nz.mem_178_sv2v_reg  <= w_data_i[18];
      \nz.mem_177_sv2v_reg  <= w_data_i[17];
      \nz.mem_176_sv2v_reg  <= w_data_i[16];
      \nz.mem_175_sv2v_reg  <= w_data_i[15];
      \nz.mem_174_sv2v_reg  <= w_data_i[14];
      \nz.mem_173_sv2v_reg  <= w_data_i[13];
      \nz.mem_172_sv2v_reg  <= w_data_i[12];
      \nz.mem_171_sv2v_reg  <= w_data_i[11];
      \nz.mem_170_sv2v_reg  <= w_data_i[10];
      \nz.mem_169_sv2v_reg  <= w_data_i[9];
      \nz.mem_168_sv2v_reg  <= w_data_i[8];
      \nz.mem_167_sv2v_reg  <= w_data_i[7];
      \nz.mem_166_sv2v_reg  <= w_data_i[6];
      \nz.mem_165_sv2v_reg  <= w_data_i[5];
      \nz.mem_164_sv2v_reg  <= w_data_i[4];
      \nz.mem_163_sv2v_reg  <= w_data_i[3];
      \nz.mem_162_sv2v_reg  <= w_data_i[2];
      \nz.mem_161_sv2v_reg  <= w_data_i[1];
      \nz.mem_160_sv2v_reg  <= w_data_i[0];
    end 
    if(N35) begin
      \nz.mem_159_sv2v_reg  <= w_data_i[79];
      \nz.mem_158_sv2v_reg  <= w_data_i[78];
      \nz.mem_157_sv2v_reg  <= w_data_i[77];
      \nz.mem_156_sv2v_reg  <= w_data_i[76];
      \nz.mem_155_sv2v_reg  <= w_data_i[75];
      \nz.mem_154_sv2v_reg  <= w_data_i[74];
      \nz.mem_153_sv2v_reg  <= w_data_i[73];
      \nz.mem_152_sv2v_reg  <= w_data_i[72];
      \nz.mem_151_sv2v_reg  <= w_data_i[71];
      \nz.mem_150_sv2v_reg  <= w_data_i[70];
      \nz.mem_149_sv2v_reg  <= w_data_i[69];
      \nz.mem_148_sv2v_reg  <= w_data_i[68];
      \nz.mem_147_sv2v_reg  <= w_data_i[67];
      \nz.mem_146_sv2v_reg  <= w_data_i[66];
      \nz.mem_145_sv2v_reg  <= w_data_i[65];
      \nz.mem_144_sv2v_reg  <= w_data_i[64];
      \nz.mem_143_sv2v_reg  <= w_data_i[63];
      \nz.mem_142_sv2v_reg  <= w_data_i[62];
      \nz.mem_141_sv2v_reg  <= w_data_i[61];
      \nz.mem_140_sv2v_reg  <= w_data_i[60];
      \nz.mem_139_sv2v_reg  <= w_data_i[59];
      \nz.mem_138_sv2v_reg  <= w_data_i[58];
      \nz.mem_137_sv2v_reg  <= w_data_i[57];
      \nz.mem_136_sv2v_reg  <= w_data_i[56];
      \nz.mem_135_sv2v_reg  <= w_data_i[55];
      \nz.mem_134_sv2v_reg  <= w_data_i[54];
      \nz.mem_133_sv2v_reg  <= w_data_i[53];
      \nz.mem_132_sv2v_reg  <= w_data_i[52];
      \nz.mem_131_sv2v_reg  <= w_data_i[51];
      \nz.mem_130_sv2v_reg  <= w_data_i[50];
      \nz.mem_129_sv2v_reg  <= w_data_i[49];
      \nz.mem_128_sv2v_reg  <= w_data_i[48];
      \nz.mem_127_sv2v_reg  <= w_data_i[47];
      \nz.mem_126_sv2v_reg  <= w_data_i[46];
      \nz.mem_125_sv2v_reg  <= w_data_i[45];
      \nz.mem_124_sv2v_reg  <= w_data_i[44];
      \nz.mem_123_sv2v_reg  <= w_data_i[43];
      \nz.mem_122_sv2v_reg  <= w_data_i[42];
      \nz.mem_121_sv2v_reg  <= w_data_i[41];
      \nz.mem_120_sv2v_reg  <= w_data_i[40];
      \nz.mem_119_sv2v_reg  <= w_data_i[39];
      \nz.mem_118_sv2v_reg  <= w_data_i[38];
      \nz.mem_117_sv2v_reg  <= w_data_i[37];
      \nz.mem_116_sv2v_reg  <= w_data_i[36];
      \nz.mem_115_sv2v_reg  <= w_data_i[35];
      \nz.mem_114_sv2v_reg  <= w_data_i[34];
      \nz.mem_113_sv2v_reg  <= w_data_i[33];
      \nz.mem_112_sv2v_reg  <= w_data_i[32];
      \nz.mem_111_sv2v_reg  <= w_data_i[31];
      \nz.mem_110_sv2v_reg  <= w_data_i[30];
      \nz.mem_109_sv2v_reg  <= w_data_i[29];
      \nz.mem_108_sv2v_reg  <= w_data_i[28];
      \nz.mem_107_sv2v_reg  <= w_data_i[27];
      \nz.mem_106_sv2v_reg  <= w_data_i[26];
      \nz.mem_105_sv2v_reg  <= w_data_i[25];
      \nz.mem_104_sv2v_reg  <= w_data_i[24];
      \nz.mem_103_sv2v_reg  <= w_data_i[23];
      \nz.mem_102_sv2v_reg  <= w_data_i[22];
      \nz.mem_101_sv2v_reg  <= w_data_i[21];
      \nz.mem_100_sv2v_reg  <= w_data_i[20];
      \nz.mem_99_sv2v_reg  <= w_data_i[19];
      \nz.mem_98_sv2v_reg  <= w_data_i[18];
      \nz.mem_97_sv2v_reg  <= w_data_i[17];
      \nz.mem_96_sv2v_reg  <= w_data_i[16];
      \nz.mem_95_sv2v_reg  <= w_data_i[15];
      \nz.mem_94_sv2v_reg  <= w_data_i[14];
      \nz.mem_93_sv2v_reg  <= w_data_i[13];
      \nz.mem_92_sv2v_reg  <= w_data_i[12];
      \nz.mem_91_sv2v_reg  <= w_data_i[11];
      \nz.mem_90_sv2v_reg  <= w_data_i[10];
      \nz.mem_89_sv2v_reg  <= w_data_i[9];
      \nz.mem_88_sv2v_reg  <= w_data_i[8];
      \nz.mem_87_sv2v_reg  <= w_data_i[7];
      \nz.mem_86_sv2v_reg  <= w_data_i[6];
      \nz.mem_85_sv2v_reg  <= w_data_i[5];
      \nz.mem_84_sv2v_reg  <= w_data_i[4];
      \nz.mem_83_sv2v_reg  <= w_data_i[3];
      \nz.mem_82_sv2v_reg  <= w_data_i[2];
      \nz.mem_81_sv2v_reg  <= w_data_i[1];
      \nz.mem_80_sv2v_reg  <= w_data_i[0];
    end 
    if(N34) begin
      \nz.mem_79_sv2v_reg  <= w_data_i[79];
      \nz.mem_78_sv2v_reg  <= w_data_i[78];
      \nz.mem_77_sv2v_reg  <= w_data_i[77];
      \nz.mem_76_sv2v_reg  <= w_data_i[76];
      \nz.mem_75_sv2v_reg  <= w_data_i[75];
      \nz.mem_74_sv2v_reg  <= w_data_i[74];
      \nz.mem_73_sv2v_reg  <= w_data_i[73];
      \nz.mem_72_sv2v_reg  <= w_data_i[72];
      \nz.mem_71_sv2v_reg  <= w_data_i[71];
      \nz.mem_70_sv2v_reg  <= w_data_i[70];
      \nz.mem_69_sv2v_reg  <= w_data_i[69];
      \nz.mem_68_sv2v_reg  <= w_data_i[68];
      \nz.mem_67_sv2v_reg  <= w_data_i[67];
      \nz.mem_66_sv2v_reg  <= w_data_i[66];
      \nz.mem_65_sv2v_reg  <= w_data_i[65];
      \nz.mem_64_sv2v_reg  <= w_data_i[64];
      \nz.mem_63_sv2v_reg  <= w_data_i[63];
      \nz.mem_62_sv2v_reg  <= w_data_i[62];
      \nz.mem_61_sv2v_reg  <= w_data_i[61];
      \nz.mem_60_sv2v_reg  <= w_data_i[60];
      \nz.mem_59_sv2v_reg  <= w_data_i[59];
      \nz.mem_58_sv2v_reg  <= w_data_i[58];
      \nz.mem_57_sv2v_reg  <= w_data_i[57];
      \nz.mem_56_sv2v_reg  <= w_data_i[56];
      \nz.mem_55_sv2v_reg  <= w_data_i[55];
      \nz.mem_54_sv2v_reg  <= w_data_i[54];
      \nz.mem_53_sv2v_reg  <= w_data_i[53];
      \nz.mem_52_sv2v_reg  <= w_data_i[52];
      \nz.mem_51_sv2v_reg  <= w_data_i[51];
      \nz.mem_50_sv2v_reg  <= w_data_i[50];
      \nz.mem_49_sv2v_reg  <= w_data_i[49];
      \nz.mem_48_sv2v_reg  <= w_data_i[48];
      \nz.mem_47_sv2v_reg  <= w_data_i[47];
      \nz.mem_46_sv2v_reg  <= w_data_i[46];
      \nz.mem_45_sv2v_reg  <= w_data_i[45];
      \nz.mem_44_sv2v_reg  <= w_data_i[44];
      \nz.mem_43_sv2v_reg  <= w_data_i[43];
      \nz.mem_42_sv2v_reg  <= w_data_i[42];
      \nz.mem_41_sv2v_reg  <= w_data_i[41];
      \nz.mem_40_sv2v_reg  <= w_data_i[40];
      \nz.mem_39_sv2v_reg  <= w_data_i[39];
      \nz.mem_38_sv2v_reg  <= w_data_i[38];
      \nz.mem_37_sv2v_reg  <= w_data_i[37];
      \nz.mem_36_sv2v_reg  <= w_data_i[36];
      \nz.mem_35_sv2v_reg  <= w_data_i[35];
      \nz.mem_34_sv2v_reg  <= w_data_i[34];
      \nz.mem_33_sv2v_reg  <= w_data_i[33];
      \nz.mem_32_sv2v_reg  <= w_data_i[32];
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_00000050_00000008
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [2:0] w_addr_i;
  input [79:0] w_data_i;
  input [2:0] r_addr_i;
  output [79:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [79:0] r_data_o;

  bsg_mem_1r1w_synth_00000050_00000008_0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bp_be_expander
(
  cinstr_i,
  instr_o
);

  input [15:0] cinstr_i;
  output [31:0] instr_o;
  wire [31:0] instr_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511;
  wire [4:3] rs1,rs2;
  wire [4:0] rd;
  wire [63:0] imm;
  assign N9 = cinstr_i[1] & N209;
  assign N10 = N212 & cinstr_i[0];
  assign N11 = N210 & N191;
  assign N12 = N11 & cinstr_i[0];
  assign N13 = N190 & N211;
  assign N14 = N13 & cinstr_i[0];
  assign N16 = cinstr_i[1] | N209;
  assign N18 = N198 & N209;
  assign N20 = N210 & N185;
  assign N21 = N20 & N209;
  assign N23 = N40 & N182;
  assign N24 = N23 & N209;
  assign N25 = N140 & N185;
  assign N26 = N25 & N209;
  assign N27 = N40 & N185;
  assign N28 = N27 & N209;
  assign N30 = N13 & N209;
  assign N31 = N41 & N209;
  assign N33 = N11 & N209;
  assign N34 = N192 & N209;
  assign N35 = N38 & N209;
  assign N36 = N43 & N209;
  assign N38 = N140 & N191;
  assign N39 = N38 & cinstr_i[0];
  assign N40 = cinstr_i[15] & cinstr_i[14];
  assign N41 = N40 & N211;
  assign N42 = N41 & cinstr_i[0];
  assign N43 = N40 & N191;
  assign N44 = N43 & cinstr_i[0];
  assign N46 = cinstr_i[15] | cinstr_i[14];
  assign N47 = cinstr_i[13] | cinstr_i[12];
  assign N48 = cinstr_i[11] | cinstr_i[10];
  assign N49 = cinstr_i[9] | cinstr_i[8];
  assign N50 = cinstr_i[7] | cinstr_i[6];
  assign N51 = cinstr_i[5] | cinstr_i[4];
  assign N52 = cinstr_i[3] | cinstr_i[2];
  assign N53 = N46 | N47;
  assign N54 = N48 | N49;
  assign N55 = N50 | N51;
  assign N56 = N52 | N16;
  assign N57 = N53 | N54;
  assign N58 = N55 | N56;
  assign N59 = N57 | N58;
  assign N60 = N74 & N65;
  assign N62 = N210 & N182;
  assign N63 = N62 & N209;
  assign N64 = N195 & N198;
  assign N65 = N64 & cinstr_i[0];
  assign N66 = N70 & N65;
  assign N68 = N208 & N194;
  assign N69 = cinstr_i[10] & N198;
  assign N70 = N140 & N68;
  assign N71 = N69 & cinstr_i[0];
  assign N72 = N70 & N71;
  assign N73 = N208 & cinstr_i[11];
  assign N74 = N140 & N73;
  assign N75 = N74 & cinstr_i[10];
  assign N76 = N208 & N209;
  assign N77 = N140 & N76;
  assign N80 = N194 & N195;
  assign N81 = N196 & N79;
  assign N82 = N197 & N133;
  assign N83 = N134 & N103;
  assign N84 = N104 & N105;
  assign N85 = N210 & N125;
  assign N86 = N80 & N81;
  assign N87 = N82 & N83;
  assign N88 = N84 & N18;
  assign N89 = N85 & N86;
  assign N90 = N87 & N88;
  assign N91 = N89 & N90;
  assign N92 = N189 | cinstr_i[14];
  assign N93 = cinstr_i[13] | N124;
  assign N94 = N198 | cinstr_i[0];
  assign N95 = N92 | N93;
  assign N96 = N52 | N94;
  assign N97 = N95 | N54;
  assign N98 = N55 | N96;
  assign N99 = N97 | N98;
  assign N101 = N126 & N108;
  assign N102 = N101 & N109;
  assign N106 = N103 & N104;
  assign N107 = N105 & cinstr_i[1];
  assign N108 = N135 & N106;
  assign N109 = N107 & N209;
  assign N110 = N144 & N108;
  assign N111 = N110 & N109;
  assign N112 = N126 & N9;
  assign N113 = N144 & N9;
  assign N114 = cinstr_i[6] & cinstr_i[5];
  assign N115 = N142 & N114;
  assign N116 = N126 & N115;
  assign N117 = N116 & N202;
  assign N118 = cinstr_i[6] & N134;
  assign N119 = N142 & N118;
  assign N120 = N126 & N119;
  assign N121 = N120 & N202;
  assign N122 = N126 & N130;
  assign N123 = N122 & N202;
  assign N125 = N208 & N124;
  assign N126 = N140 & N125;
  assign N127 = N126 & N136;
  assign N128 = N127 & N202;
  assign N129 = N133 & cinstr_i[5];
  assign N130 = N142 & N129;
  assign N131 = N144 & N130;
  assign N132 = N131 & N202;
  assign N135 = N133 & N134;
  assign N136 = N142 & N135;
  assign N137 = N144 & N136;
  assign N138 = N137 & N202;
  assign N139 = cinstr_i[1] & cinstr_i[0];
  assign N140 = cinstr_i[15] & N207;
  assign N141 = N208 & cinstr_i[12];
  assign N142 = cinstr_i[11] & cinstr_i[10];
  assign N143 = cinstr_i[6] & cinstr_i[0];
  assign N144 = N140 & N141;
  assign N145 = N142 & N143;
  assign N146 = N144 & N145;
  assign N147 = N140 & N211;
  assign N148 = N147 & N209;
  assign N182 = N208 & cinstr_i[1];
  assign N183 = N190 & N182;
  assign N184 = N183 & N209;
  assign N185 = cinstr_i[13] & cinstr_i[1];
  assign N186 = N190 & N185;
  assign N187 = N186 & N209;
  assign N190 = N189 & cinstr_i[14];
  assign N191 = cinstr_i[13] & N198;
  assign N192 = N190 & N191;
  assign N193 = N192 & cinstr_i[0];
  assign N199 = cinstr_i[13] & N194;
  assign N200 = N195 & N196;
  assign N201 = cinstr_i[8] & N197;
  assign N202 = N198 & cinstr_i[0];
  assign N203 = N190 & N199;
  assign N204 = N200 & N201;
  assign N205 = N203 & N204;
  assign N206 = N205 & N202;
  assign N210 = N189 & N207;
  assign N211 = N208 & N198;
  assign N212 = N210 & N211;
  assign N213 = N212 & N209;
  assign rs1 = (N0)? cinstr_i[11:10] : 
               (N284)? { 1'b0, 1'b1 } : 
               (N286)? { 1'b0, 1'b1 } : 1'b0;
  assign N0 = N15;
  assign rs2 = (N0)? cinstr_i[6:5] : 
               (N284)? { 1'b0, 1'b1 } : 
               (N286)? { 1'b0, 1'b1 } : 1'b0;
  assign rd = (N0)? cinstr_i[11:7] : 
              (N284)? { 1'b0, 1'b1, cinstr_i[9:7] } : 
              (N286)? { 1'b0, 1'b1, cinstr_i[4:2] } : 1'b0;
  assign imm = (N1)? { cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[4:3], cinstr_i[5:5], cinstr_i[2:2], cinstr_i[6:6], 1'b0, 1'b0, 1'b0, 1'b0 } : 
               (N288)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[10:7], cinstr_i[12:11], cinstr_i[5:5], cinstr_i[6:6], 1'b0, 1'b0 } : 
               (N291)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[3:2], cinstr_i[12:12], cinstr_i[6:4], 1'b0, 1'b0 } : 
               (N294)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[4:2], cinstr_i[12:12], cinstr_i[6:5], 1'b0, 1'b0, 1'b0 } : 
               (N297)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[8:7], cinstr_i[12:9], 1'b0, 1'b0 } : 
               (N300)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[9:7], cinstr_i[12:10], 1'b0, 1'b0, 1'b0 } : 
               (N303)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[5:5], cinstr_i[12:10], cinstr_i[6:6], 1'b0, 1'b0 } : 
               (N306)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[6:5], cinstr_i[12:10], 1'b0, 1'b0, 1'b0 } : 
               (N309)? { cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[8:8], cinstr_i[10:9], cinstr_i[6:6], cinstr_i[7:7], cinstr_i[2:2], cinstr_i[11:11], cinstr_i[5:3], 1'b0 } : 
               (N312)? { cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[6:5], cinstr_i[2:2], cinstr_i[11:10], cinstr_i[4:3], 1'b0 } : 
               (N315)? { cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[6:2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
               (N318)? { cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[12:12], cinstr_i[6:2] } : 
               (N321)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[12:12], cinstr_i[6:2] } : 
               (N324)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i[12:12], cinstr_i[6:2] } : 
               (N327)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = N206;
  assign { N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150 } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N329)? { imm[11:0], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N331)? { imm[11:0], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N333)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N335)? { imm[11:0], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, rd, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N337)? { imm[11:0], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, rd, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N340)? { imm[11:5], rs2, cinstr_i[4:2], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, imm[4:0], 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N342)? { imm[11:5], rs2, cinstr_i[4:2], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, imm[4:0], 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N345)? { imm[11:0], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, rd, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N348)? { imm[11:5], rs2, cinstr_i[4:2], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, imm[4:0], 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N351)? { imm[11:0], rs1, cinstr_i[9:7], 1'b0, 1'b1, 1'b0, rd, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N354)? { imm[11:0], rs1, cinstr_i[9:7], 1'b0, 1'b1, 1'b1, rd, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N357)? { imm[11:5], rs2, cinstr_i[4:2], rs1, cinstr_i[9:7], 1'b0, 1'b1, 1'b0, imm[4:0], 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N360)? { imm[11:5], rs2, cinstr_i[4:2], rs1, cinstr_i[9:7], 1'b0, 1'b1, 1'b1, imm[4:0], 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N363)? { imm[11:0], rs1, cinstr_i[9:7], 1'b0, 1'b1, 1'b1, rd, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N366)? { imm[11:5], rs2, cinstr_i[4:2], rs1, cinstr_i[9:7], 1'b0, 1'b1, 1'b1, imm[4:0], 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N369)? { imm[20:20], imm[10:1], imm[11:11], imm[19:12], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N371)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs1, cinstr_i[9:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N374)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs1, cinstr_i[9:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N377)? { imm[12:12], imm[10:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs1, cinstr_i[9:7], 1'b0, 1'b0, 1'b0, imm[4:1], imm[11:11], 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N380)? { imm[12:12], imm[10:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs1, cinstr_i[9:7], 1'b0, 1'b0, 1'b1, imm[4:1], imm[11:11], 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N383)? { imm[11:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N386)? { imm[31:12], rd, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N388)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N390)? { imm[11:0], rd, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N393)? { imm[11:0], rd, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N396)? { imm[11:0], rd, 1'b0, 1'b0, 1'b1, rd, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N399)? { imm[11:0], rd, 1'b1, 1'b0, 1'b1, rd, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N402)? { imm[11:0], rd, 1'b1, 1'b0, 1'b1, rd, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N404)? { imm[11:0], rd, 1'b1, 1'b1, 1'b1, rd, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N407)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs2, cinstr_i[4:2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N410)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs2, cinstr_i[4:2], rd, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N413)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs2, cinstr_i[4:2], rd, 1'b1, 1'b1, 1'b1, rd, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N416)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs2, cinstr_i[4:2], rd, 1'b1, 1'b1, 1'b0, rd, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N419)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs2, cinstr_i[4:2], rd, 1'b1, 1'b0, 1'b0, rd, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N422)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs2, cinstr_i[4:2], rd, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N425)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs2, cinstr_i[4:2], rd, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N428)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rs2, cinstr_i[4:2], rd, 1'b0, 1'b0, 1'b0, rd, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N431)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cinstr_i } : 1'b0;
  assign N2 = N91;
  assign { N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218 } = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N4)? { N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150 } : 1'b0;
  assign N3 = N217;
  assign N4 = N448;
  assign { N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N6)? { N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150 } : 1'b0;
  assign N5 = N250;
  assign N6 = N511;
  assign instr_o = (N7)? { N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218 } : 
                   (N8)? { N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251 } : 
                   (N216)? { N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150 } : 1'b0;
  assign N7 = N188;
  assign N8 = N214;
  assign N15 = N435 | N193;
  assign N435 = N434 | N206;
  assign N434 = N433 | N14;
  assign N433 = N432 | N12;
  assign N432 = N9 | N10;
  assign N17 = ~N16;
  assign N19 = N139 | N18;
  assign N22 = N21 | N187;
  assign N29 = N26 | N28;
  assign N32 = N30 | N31;
  assign N37 = N437 | N36;
  assign N437 = N436 | N35;
  assign N436 = N33 | N34;
  assign N45 = N42 | N44;
  assign N61 = N441 | N60;
  assign N441 = N440 | N14;
  assign N440 = N439 | N12;
  assign N439 = N438 | N10;
  assign N438 = ~N59;
  assign N67 = N63 | N66;
  assign N78 = N139 | N442;
  assign N442 = N75 | N77;
  assign N79 = ~cinstr_i[8];
  assign N100 = ~N99;
  assign N103 = ~cinstr_i[4];
  assign N104 = ~cinstr_i[3];
  assign N105 = ~cinstr_i[2];
  assign N124 = ~cinstr_i[12];
  assign N133 = ~cinstr_i[6];
  assign N134 = ~cinstr_i[5];
  assign N149 = N139 | N443;
  assign N443 = N146 | N148;
  assign N188 = N184 | N187;
  assign N189 = ~cinstr_i[15];
  assign N194 = ~cinstr_i[11];
  assign N195 = ~cinstr_i[10];
  assign N196 = ~cinstr_i[9];
  assign N197 = ~cinstr_i[7];
  assign N198 = ~cinstr_i[1];
  assign N207 = ~cinstr_i[14];
  assign N208 = ~cinstr_i[13];
  assign N209 = ~cinstr_i[0];
  assign N214 = N444 | N213;
  assign N444 = N193 | N206;
  assign N215 = N214 | N188;
  assign N216 = ~N215;
  assign N217 = ~N448;
  assign N448 = N447 | cinstr_i[7];
  assign N447 = N446 | cinstr_i[8];
  assign N446 = N445 | cinstr_i[9];
  assign N445 = cinstr_i[11] | cinstr_i[10];
  assign N250 = ~N511;
  assign N511 = N510 | imm[0];
  assign N510 = N509 | imm[1];
  assign N509 = N508 | imm[2];
  assign N508 = N507 | imm[3];
  assign N507 = N506 | imm[4];
  assign N506 = N505 | imm[5];
  assign N505 = N504 | imm[6];
  assign N504 = N503 | imm[7];
  assign N503 = N502 | imm[8];
  assign N502 = N501 | imm[9];
  assign N501 = N500 | imm[10];
  assign N500 = N499 | imm[11];
  assign N499 = N498 | imm[12];
  assign N498 = N497 | imm[13];
  assign N497 = N496 | imm[14];
  assign N496 = N495 | imm[15];
  assign N495 = N494 | imm[16];
  assign N494 = N493 | imm[17];
  assign N493 = N492 | imm[18];
  assign N492 = N491 | imm[19];
  assign N491 = N490 | imm[20];
  assign N490 = N489 | imm[21];
  assign N489 = N488 | imm[22];
  assign N488 = N487 | imm[23];
  assign N487 = N486 | imm[24];
  assign N486 = N485 | imm[25];
  assign N485 = N484 | imm[26];
  assign N484 = N483 | imm[27];
  assign N483 = N482 | imm[28];
  assign N482 = N481 | imm[29];
  assign N481 = N480 | imm[30];
  assign N480 = N479 | imm[31];
  assign N479 = N478 | imm[32];
  assign N478 = N477 | imm[33];
  assign N477 = N476 | imm[34];
  assign N476 = N475 | imm[35];
  assign N475 = N474 | imm[36];
  assign N474 = N473 | imm[37];
  assign N473 = N472 | imm[38];
  assign N472 = N471 | imm[39];
  assign N471 = N470 | imm[40];
  assign N470 = N469 | imm[41];
  assign N469 = N468 | imm[42];
  assign N468 = N467 | imm[43];
  assign N467 = N466 | imm[44];
  assign N466 = N465 | imm[45];
  assign N465 = N464 | imm[46];
  assign N464 = N463 | imm[47];
  assign N463 = N462 | imm[48];
  assign N462 = N461 | imm[49];
  assign N461 = N460 | imm[50];
  assign N460 = N459 | imm[51];
  assign N459 = N458 | imm[52];
  assign N458 = N457 | imm[53];
  assign N457 = N456 | imm[54];
  assign N456 = N455 | imm[55];
  assign N455 = N454 | imm[56];
  assign N454 = N453 | imm[57];
  assign N453 = N452 | imm[58];
  assign N452 = N451 | imm[59];
  assign N451 = N450 | imm[60];
  assign N450 = N449 | imm[61];
  assign N449 = imm[63] | imm[62];
  assign N283 = ~N15;
  assign N284 = N17 & N283;
  assign N285 = N283 & N16;
  assign N286 = N19 & N285;
  assign N287 = ~N206;
  assign N288 = N213 & N287;
  assign N289 = ~N213;
  assign N290 = N287 & N289;
  assign N291 = N184 & N290;
  assign N292 = ~N184;
  assign N293 = N290 & N292;
  assign N294 = N22 & N293;
  assign N295 = ~N22;
  assign N296 = N293 & N295;
  assign N297 = N24 & N296;
  assign N298 = ~N24;
  assign N299 = N296 & N298;
  assign N300 = N29 & N299;
  assign N301 = ~N29;
  assign N302 = N299 & N301;
  assign N303 = N32 & N302;
  assign N304 = ~N32;
  assign N305 = N302 & N304;
  assign N306 = N37 & N305;
  assign N307 = ~N37;
  assign N308 = N305 & N307;
  assign N309 = N39 & N308;
  assign N310 = ~N39;
  assign N311 = N308 & N310;
  assign N312 = N45 & N311;
  assign N313 = ~N45;
  assign N314 = N311 & N313;
  assign N315 = N193 & N314;
  assign N316 = ~N193;
  assign N317 = N314 & N316;
  assign N318 = N61 & N317;
  assign N319 = ~N61;
  assign N320 = N317 & N319;
  assign N321 = N67 & N320;
  assign N322 = ~N67;
  assign N323 = N320 & N322;
  assign N324 = N72 & N323;
  assign N325 = ~N72;
  assign N326 = N323 & N325;
  assign N327 = N78 & N326;
  assign N328 = ~N91;
  assign N329 = N213 & N328;
  assign N330 = N328 & N289;
  assign N331 = N206 & N330;
  assign N332 = N330 & N287;
  assign N333 = N100 & N332;
  assign N334 = N332 & N99;
  assign N335 = N184 & N334;
  assign N336 = N334 & N292;
  assign N337 = N187 & N336;
  assign N338 = ~N187;
  assign N339 = N336 & N338;
  assign N340 = N24 & N339;
  assign N341 = N339 & N298;
  assign N342 = N28 & N341;
  assign N343 = ~N28;
  assign N344 = N341 & N343;
  assign N345 = N21 & N344;
  assign N346 = ~N21;
  assign N347 = N344 & N346;
  assign N348 = N26 & N347;
  assign N349 = ~N26;
  assign N350 = N347 & N349;
  assign N351 = N30 & N350;
  assign N352 = ~N30;
  assign N353 = N350 & N352;
  assign N354 = N34 & N353;
  assign N355 = ~N34;
  assign N356 = N353 & N355;
  assign N357 = N31 & N356;
  assign N358 = ~N31;
  assign N359 = N356 & N358;
  assign N360 = N36 & N359;
  assign N361 = ~N36;
  assign N362 = N359 & N361;
  assign N363 = N33 & N362;
  assign N364 = ~N33;
  assign N365 = N362 & N364;
  assign N366 = N35 & N365;
  assign N367 = ~N35;
  assign N368 = N365 & N367;
  assign N369 = N39 & N368;
  assign N370 = N368 & N310;
  assign N371 = N102 & N370;
  assign N372 = ~N102;
  assign N373 = N370 & N372;
  assign N374 = N111 & N373;
  assign N375 = ~N111;
  assign N376 = N373 & N375;
  assign N377 = N42 & N376;
  assign N378 = ~N42;
  assign N379 = N376 & N378;
  assign N380 = N44 & N379;
  assign N381 = ~N44;
  assign N382 = N379 & N381;
  assign N383 = N14 & N382;
  assign N384 = ~N14;
  assign N385 = N382 & N384;
  assign N386 = N193 & N385;
  assign N387 = N385 & N316;
  assign N388 = N438 & N387;
  assign N389 = N387 & N59;
  assign N390 = N10 & N389;
  assign N391 = ~N10;
  assign N392 = N389 & N391;
  assign N393 = N12 & N392;
  assign N394 = ~N12;
  assign N395 = N392 & N394;
  assign N396 = N63 & N395;
  assign N397 = ~N63;
  assign N398 = N395 & N397;
  assign N399 = N66 & N398;
  assign N400 = ~N66;
  assign N401 = N398 & N400;
  assign N402 = N72 & N401;
  assign N403 = N401 & N325;
  assign N404 = N60 & N403;
  assign N405 = ~N60;
  assign N406 = N403 & N405;
  assign N407 = N112 & N406;
  assign N408 = ~N112;
  assign N409 = N406 & N408;
  assign N410 = N113 & N409;
  assign N411 = ~N113;
  assign N412 = N409 & N411;
  assign N413 = N117 & N412;
  assign N414 = ~N117;
  assign N415 = N412 & N414;
  assign N416 = N121 & N415;
  assign N417 = ~N121;
  assign N418 = N415 & N417;
  assign N419 = N123 & N418;
  assign N420 = ~N123;
  assign N421 = N418 & N420;
  assign N422 = N128 & N421;
  assign N423 = ~N128;
  assign N424 = N421 & N423;
  assign N425 = N132 & N424;
  assign N426 = ~N132;
  assign N427 = N424 & N426;
  assign N428 = N138 & N427;
  assign N429 = ~N138;
  assign N430 = N427 & N429;
  assign N431 = N149 & N430;

endmodule



module bsg_dff_reset_en_width_p39
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [38:0] data_i;
  output [38:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [38:0] data_o;
  wire N0,N1,N2;
  reg data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,
  data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,
  data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,
  data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,
  data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,
  data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_synth_000000ae_00000008_0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [2:0] w_addr_i;
  input [173:0] w_data_i;
  input [2:0] r_addr_i;
  output [173:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [173:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53;
  wire [1391:0] \nz.mem ;
  reg \nz.mem_1391_sv2v_reg ,\nz.mem_1390_sv2v_reg ,\nz.mem_1389_sv2v_reg ,
  \nz.mem_1388_sv2v_reg ,\nz.mem_1387_sv2v_reg ,\nz.mem_1386_sv2v_reg ,
  \nz.mem_1385_sv2v_reg ,\nz.mem_1384_sv2v_reg ,\nz.mem_1383_sv2v_reg ,\nz.mem_1382_sv2v_reg ,
  \nz.mem_1381_sv2v_reg ,\nz.mem_1380_sv2v_reg ,\nz.mem_1379_sv2v_reg ,
  \nz.mem_1378_sv2v_reg ,\nz.mem_1377_sv2v_reg ,\nz.mem_1376_sv2v_reg ,\nz.mem_1375_sv2v_reg ,
  \nz.mem_1374_sv2v_reg ,\nz.mem_1373_sv2v_reg ,\nz.mem_1372_sv2v_reg ,
  \nz.mem_1371_sv2v_reg ,\nz.mem_1370_sv2v_reg ,\nz.mem_1369_sv2v_reg ,\nz.mem_1368_sv2v_reg ,
  \nz.mem_1367_sv2v_reg ,\nz.mem_1366_sv2v_reg ,\nz.mem_1365_sv2v_reg ,
  \nz.mem_1364_sv2v_reg ,\nz.mem_1363_sv2v_reg ,\nz.mem_1362_sv2v_reg ,\nz.mem_1361_sv2v_reg ,
  \nz.mem_1360_sv2v_reg ,\nz.mem_1359_sv2v_reg ,\nz.mem_1358_sv2v_reg ,
  \nz.mem_1357_sv2v_reg ,\nz.mem_1356_sv2v_reg ,\nz.mem_1355_sv2v_reg ,\nz.mem_1354_sv2v_reg ,
  \nz.mem_1353_sv2v_reg ,\nz.mem_1352_sv2v_reg ,\nz.mem_1351_sv2v_reg ,
  \nz.mem_1350_sv2v_reg ,\nz.mem_1349_sv2v_reg ,\nz.mem_1348_sv2v_reg ,\nz.mem_1347_sv2v_reg ,
  \nz.mem_1346_sv2v_reg ,\nz.mem_1345_sv2v_reg ,\nz.mem_1344_sv2v_reg ,
  \nz.mem_1343_sv2v_reg ,\nz.mem_1342_sv2v_reg ,\nz.mem_1341_sv2v_reg ,\nz.mem_1340_sv2v_reg ,
  \nz.mem_1339_sv2v_reg ,\nz.mem_1338_sv2v_reg ,\nz.mem_1337_sv2v_reg ,
  \nz.mem_1336_sv2v_reg ,\nz.mem_1335_sv2v_reg ,\nz.mem_1334_sv2v_reg ,\nz.mem_1333_sv2v_reg ,
  \nz.mem_1332_sv2v_reg ,\nz.mem_1331_sv2v_reg ,\nz.mem_1330_sv2v_reg ,
  \nz.mem_1329_sv2v_reg ,\nz.mem_1328_sv2v_reg ,\nz.mem_1327_sv2v_reg ,\nz.mem_1326_sv2v_reg ,
  \nz.mem_1325_sv2v_reg ,\nz.mem_1324_sv2v_reg ,\nz.mem_1323_sv2v_reg ,
  \nz.mem_1322_sv2v_reg ,\nz.mem_1321_sv2v_reg ,\nz.mem_1320_sv2v_reg ,\nz.mem_1319_sv2v_reg ,
  \nz.mem_1318_sv2v_reg ,\nz.mem_1317_sv2v_reg ,\nz.mem_1316_sv2v_reg ,
  \nz.mem_1315_sv2v_reg ,\nz.mem_1314_sv2v_reg ,\nz.mem_1313_sv2v_reg ,\nz.mem_1312_sv2v_reg ,
  \nz.mem_1311_sv2v_reg ,\nz.mem_1310_sv2v_reg ,\nz.mem_1309_sv2v_reg ,
  \nz.mem_1308_sv2v_reg ,\nz.mem_1307_sv2v_reg ,\nz.mem_1306_sv2v_reg ,
  \nz.mem_1305_sv2v_reg ,\nz.mem_1304_sv2v_reg ,\nz.mem_1303_sv2v_reg ,\nz.mem_1302_sv2v_reg ,
  \nz.mem_1301_sv2v_reg ,\nz.mem_1300_sv2v_reg ,\nz.mem_1299_sv2v_reg ,
  \nz.mem_1298_sv2v_reg ,\nz.mem_1297_sv2v_reg ,\nz.mem_1296_sv2v_reg ,\nz.mem_1295_sv2v_reg ,
  \nz.mem_1294_sv2v_reg ,\nz.mem_1293_sv2v_reg ,\nz.mem_1292_sv2v_reg ,
  \nz.mem_1291_sv2v_reg ,\nz.mem_1290_sv2v_reg ,\nz.mem_1289_sv2v_reg ,\nz.mem_1288_sv2v_reg ,
  \nz.mem_1287_sv2v_reg ,\nz.mem_1286_sv2v_reg ,\nz.mem_1285_sv2v_reg ,
  \nz.mem_1284_sv2v_reg ,\nz.mem_1283_sv2v_reg ,\nz.mem_1282_sv2v_reg ,\nz.mem_1281_sv2v_reg ,
  \nz.mem_1280_sv2v_reg ,\nz.mem_1279_sv2v_reg ,\nz.mem_1278_sv2v_reg ,
  \nz.mem_1277_sv2v_reg ,\nz.mem_1276_sv2v_reg ,\nz.mem_1275_sv2v_reg ,\nz.mem_1274_sv2v_reg ,
  \nz.mem_1273_sv2v_reg ,\nz.mem_1272_sv2v_reg ,\nz.mem_1271_sv2v_reg ,
  \nz.mem_1270_sv2v_reg ,\nz.mem_1269_sv2v_reg ,\nz.mem_1268_sv2v_reg ,\nz.mem_1267_sv2v_reg ,
  \nz.mem_1266_sv2v_reg ,\nz.mem_1265_sv2v_reg ,\nz.mem_1264_sv2v_reg ,
  \nz.mem_1263_sv2v_reg ,\nz.mem_1262_sv2v_reg ,\nz.mem_1261_sv2v_reg ,\nz.mem_1260_sv2v_reg ,
  \nz.mem_1259_sv2v_reg ,\nz.mem_1258_sv2v_reg ,\nz.mem_1257_sv2v_reg ,
  \nz.mem_1256_sv2v_reg ,\nz.mem_1255_sv2v_reg ,\nz.mem_1254_sv2v_reg ,\nz.mem_1253_sv2v_reg ,
  \nz.mem_1252_sv2v_reg ,\nz.mem_1251_sv2v_reg ,\nz.mem_1250_sv2v_reg ,
  \nz.mem_1249_sv2v_reg ,\nz.mem_1248_sv2v_reg ,\nz.mem_1247_sv2v_reg ,\nz.mem_1246_sv2v_reg ,
  \nz.mem_1245_sv2v_reg ,\nz.mem_1244_sv2v_reg ,\nz.mem_1243_sv2v_reg ,
  \nz.mem_1242_sv2v_reg ,\nz.mem_1241_sv2v_reg ,\nz.mem_1240_sv2v_reg ,\nz.mem_1239_sv2v_reg ,
  \nz.mem_1238_sv2v_reg ,\nz.mem_1237_sv2v_reg ,\nz.mem_1236_sv2v_reg ,
  \nz.mem_1235_sv2v_reg ,\nz.mem_1234_sv2v_reg ,\nz.mem_1233_sv2v_reg ,\nz.mem_1232_sv2v_reg ,
  \nz.mem_1231_sv2v_reg ,\nz.mem_1230_sv2v_reg ,\nz.mem_1229_sv2v_reg ,
  \nz.mem_1228_sv2v_reg ,\nz.mem_1227_sv2v_reg ,\nz.mem_1226_sv2v_reg ,
  \nz.mem_1225_sv2v_reg ,\nz.mem_1224_sv2v_reg ,\nz.mem_1223_sv2v_reg ,\nz.mem_1222_sv2v_reg ,
  \nz.mem_1221_sv2v_reg ,\nz.mem_1220_sv2v_reg ,\nz.mem_1219_sv2v_reg ,
  \nz.mem_1218_sv2v_reg ,\nz.mem_1217_sv2v_reg ,\nz.mem_1216_sv2v_reg ,\nz.mem_1215_sv2v_reg ,
  \nz.mem_1214_sv2v_reg ,\nz.mem_1213_sv2v_reg ,\nz.mem_1212_sv2v_reg ,
  \nz.mem_1211_sv2v_reg ,\nz.mem_1210_sv2v_reg ,\nz.mem_1209_sv2v_reg ,\nz.mem_1208_sv2v_reg ,
  \nz.mem_1207_sv2v_reg ,\nz.mem_1206_sv2v_reg ,\nz.mem_1205_sv2v_reg ,
  \nz.mem_1204_sv2v_reg ,\nz.mem_1203_sv2v_reg ,\nz.mem_1202_sv2v_reg ,\nz.mem_1201_sv2v_reg ,
  \nz.mem_1200_sv2v_reg ,\nz.mem_1199_sv2v_reg ,\nz.mem_1198_sv2v_reg ,
  \nz.mem_1197_sv2v_reg ,\nz.mem_1196_sv2v_reg ,\nz.mem_1195_sv2v_reg ,\nz.mem_1194_sv2v_reg ,
  \nz.mem_1193_sv2v_reg ,\nz.mem_1192_sv2v_reg ,\nz.mem_1191_sv2v_reg ,
  \nz.mem_1190_sv2v_reg ,\nz.mem_1189_sv2v_reg ,\nz.mem_1188_sv2v_reg ,\nz.mem_1187_sv2v_reg ,
  \nz.mem_1186_sv2v_reg ,\nz.mem_1185_sv2v_reg ,\nz.mem_1184_sv2v_reg ,
  \nz.mem_1183_sv2v_reg ,\nz.mem_1182_sv2v_reg ,\nz.mem_1181_sv2v_reg ,\nz.mem_1180_sv2v_reg ,
  \nz.mem_1179_sv2v_reg ,\nz.mem_1178_sv2v_reg ,\nz.mem_1177_sv2v_reg ,
  \nz.mem_1176_sv2v_reg ,\nz.mem_1175_sv2v_reg ,\nz.mem_1174_sv2v_reg ,\nz.mem_1173_sv2v_reg ,
  \nz.mem_1172_sv2v_reg ,\nz.mem_1171_sv2v_reg ,\nz.mem_1170_sv2v_reg ,
  \nz.mem_1169_sv2v_reg ,\nz.mem_1168_sv2v_reg ,\nz.mem_1167_sv2v_reg ,\nz.mem_1166_sv2v_reg ,
  \nz.mem_1165_sv2v_reg ,\nz.mem_1164_sv2v_reg ,\nz.mem_1163_sv2v_reg ,
  \nz.mem_1162_sv2v_reg ,\nz.mem_1161_sv2v_reg ,\nz.mem_1160_sv2v_reg ,\nz.mem_1159_sv2v_reg ,
  \nz.mem_1158_sv2v_reg ,\nz.mem_1157_sv2v_reg ,\nz.mem_1156_sv2v_reg ,
  \nz.mem_1155_sv2v_reg ,\nz.mem_1154_sv2v_reg ,\nz.mem_1153_sv2v_reg ,\nz.mem_1152_sv2v_reg ,
  \nz.mem_1151_sv2v_reg ,\nz.mem_1150_sv2v_reg ,\nz.mem_1149_sv2v_reg ,
  \nz.mem_1148_sv2v_reg ,\nz.mem_1147_sv2v_reg ,\nz.mem_1146_sv2v_reg ,
  \nz.mem_1145_sv2v_reg ,\nz.mem_1144_sv2v_reg ,\nz.mem_1143_sv2v_reg ,\nz.mem_1142_sv2v_reg ,
  \nz.mem_1141_sv2v_reg ,\nz.mem_1140_sv2v_reg ,\nz.mem_1139_sv2v_reg ,
  \nz.mem_1138_sv2v_reg ,\nz.mem_1137_sv2v_reg ,\nz.mem_1136_sv2v_reg ,\nz.mem_1135_sv2v_reg ,
  \nz.mem_1134_sv2v_reg ,\nz.mem_1133_sv2v_reg ,\nz.mem_1132_sv2v_reg ,
  \nz.mem_1131_sv2v_reg ,\nz.mem_1130_sv2v_reg ,\nz.mem_1129_sv2v_reg ,\nz.mem_1128_sv2v_reg ,
  \nz.mem_1127_sv2v_reg ,\nz.mem_1126_sv2v_reg ,\nz.mem_1125_sv2v_reg ,
  \nz.mem_1124_sv2v_reg ,\nz.mem_1123_sv2v_reg ,\nz.mem_1122_sv2v_reg ,\nz.mem_1121_sv2v_reg ,
  \nz.mem_1120_sv2v_reg ,\nz.mem_1119_sv2v_reg ,\nz.mem_1118_sv2v_reg ,
  \nz.mem_1117_sv2v_reg ,\nz.mem_1116_sv2v_reg ,\nz.mem_1115_sv2v_reg ,\nz.mem_1114_sv2v_reg ,
  \nz.mem_1113_sv2v_reg ,\nz.mem_1112_sv2v_reg ,\nz.mem_1111_sv2v_reg ,
  \nz.mem_1110_sv2v_reg ,\nz.mem_1109_sv2v_reg ,\nz.mem_1108_sv2v_reg ,\nz.mem_1107_sv2v_reg ,
  \nz.mem_1106_sv2v_reg ,\nz.mem_1105_sv2v_reg ,\nz.mem_1104_sv2v_reg ,
  \nz.mem_1103_sv2v_reg ,\nz.mem_1102_sv2v_reg ,\nz.mem_1101_sv2v_reg ,\nz.mem_1100_sv2v_reg ,
  \nz.mem_1099_sv2v_reg ,\nz.mem_1098_sv2v_reg ,\nz.mem_1097_sv2v_reg ,
  \nz.mem_1096_sv2v_reg ,\nz.mem_1095_sv2v_reg ,\nz.mem_1094_sv2v_reg ,\nz.mem_1093_sv2v_reg ,
  \nz.mem_1092_sv2v_reg ,\nz.mem_1091_sv2v_reg ,\nz.mem_1090_sv2v_reg ,
  \nz.mem_1089_sv2v_reg ,\nz.mem_1088_sv2v_reg ,\nz.mem_1087_sv2v_reg ,\nz.mem_1086_sv2v_reg ,
  \nz.mem_1085_sv2v_reg ,\nz.mem_1084_sv2v_reg ,\nz.mem_1083_sv2v_reg ,
  \nz.mem_1082_sv2v_reg ,\nz.mem_1081_sv2v_reg ,\nz.mem_1080_sv2v_reg ,\nz.mem_1079_sv2v_reg ,
  \nz.mem_1078_sv2v_reg ,\nz.mem_1077_sv2v_reg ,\nz.mem_1076_sv2v_reg ,
  \nz.mem_1075_sv2v_reg ,\nz.mem_1074_sv2v_reg ,\nz.mem_1073_sv2v_reg ,\nz.mem_1072_sv2v_reg ,
  \nz.mem_1071_sv2v_reg ,\nz.mem_1070_sv2v_reg ,\nz.mem_1069_sv2v_reg ,
  \nz.mem_1068_sv2v_reg ,\nz.mem_1067_sv2v_reg ,\nz.mem_1066_sv2v_reg ,
  \nz.mem_1065_sv2v_reg ,\nz.mem_1064_sv2v_reg ,\nz.mem_1063_sv2v_reg ,\nz.mem_1062_sv2v_reg ,
  \nz.mem_1061_sv2v_reg ,\nz.mem_1060_sv2v_reg ,\nz.mem_1059_sv2v_reg ,
  \nz.mem_1058_sv2v_reg ,\nz.mem_1057_sv2v_reg ,\nz.mem_1056_sv2v_reg ,\nz.mem_1055_sv2v_reg ,
  \nz.mem_1054_sv2v_reg ,\nz.mem_1053_sv2v_reg ,\nz.mem_1052_sv2v_reg ,
  \nz.mem_1051_sv2v_reg ,\nz.mem_1050_sv2v_reg ,\nz.mem_1049_sv2v_reg ,\nz.mem_1048_sv2v_reg ,
  \nz.mem_1047_sv2v_reg ,\nz.mem_1046_sv2v_reg ,\nz.mem_1045_sv2v_reg ,
  \nz.mem_1044_sv2v_reg ,\nz.mem_1043_sv2v_reg ,\nz.mem_1042_sv2v_reg ,\nz.mem_1041_sv2v_reg ,
  \nz.mem_1040_sv2v_reg ,\nz.mem_1039_sv2v_reg ,\nz.mem_1038_sv2v_reg ,
  \nz.mem_1037_sv2v_reg ,\nz.mem_1036_sv2v_reg ,\nz.mem_1035_sv2v_reg ,\nz.mem_1034_sv2v_reg ,
  \nz.mem_1033_sv2v_reg ,\nz.mem_1032_sv2v_reg ,\nz.mem_1031_sv2v_reg ,
  \nz.mem_1030_sv2v_reg ,\nz.mem_1029_sv2v_reg ,\nz.mem_1028_sv2v_reg ,\nz.mem_1027_sv2v_reg ,
  \nz.mem_1026_sv2v_reg ,\nz.mem_1025_sv2v_reg ,\nz.mem_1024_sv2v_reg ,
  \nz.mem_1023_sv2v_reg ,\nz.mem_1022_sv2v_reg ,\nz.mem_1021_sv2v_reg ,\nz.mem_1020_sv2v_reg ,
  \nz.mem_1019_sv2v_reg ,\nz.mem_1018_sv2v_reg ,\nz.mem_1017_sv2v_reg ,
  \nz.mem_1016_sv2v_reg ,\nz.mem_1015_sv2v_reg ,\nz.mem_1014_sv2v_reg ,\nz.mem_1013_sv2v_reg ,
  \nz.mem_1012_sv2v_reg ,\nz.mem_1011_sv2v_reg ,\nz.mem_1010_sv2v_reg ,
  \nz.mem_1009_sv2v_reg ,\nz.mem_1008_sv2v_reg ,\nz.mem_1007_sv2v_reg ,\nz.mem_1006_sv2v_reg ,
  \nz.mem_1005_sv2v_reg ,\nz.mem_1004_sv2v_reg ,\nz.mem_1003_sv2v_reg ,
  \nz.mem_1002_sv2v_reg ,\nz.mem_1001_sv2v_reg ,\nz.mem_1000_sv2v_reg ,\nz.mem_999_sv2v_reg ,
  \nz.mem_998_sv2v_reg ,\nz.mem_997_sv2v_reg ,\nz.mem_996_sv2v_reg ,
  \nz.mem_995_sv2v_reg ,\nz.mem_994_sv2v_reg ,\nz.mem_993_sv2v_reg ,\nz.mem_992_sv2v_reg ,
  \nz.mem_991_sv2v_reg ,\nz.mem_990_sv2v_reg ,\nz.mem_989_sv2v_reg ,\nz.mem_988_sv2v_reg ,
  \nz.mem_987_sv2v_reg ,\nz.mem_986_sv2v_reg ,\nz.mem_985_sv2v_reg ,
  \nz.mem_984_sv2v_reg ,\nz.mem_983_sv2v_reg ,\nz.mem_982_sv2v_reg ,\nz.mem_981_sv2v_reg ,
  \nz.mem_980_sv2v_reg ,\nz.mem_979_sv2v_reg ,\nz.mem_978_sv2v_reg ,
  \nz.mem_977_sv2v_reg ,\nz.mem_976_sv2v_reg ,\nz.mem_975_sv2v_reg ,\nz.mem_974_sv2v_reg ,
  \nz.mem_973_sv2v_reg ,\nz.mem_972_sv2v_reg ,\nz.mem_971_sv2v_reg ,\nz.mem_970_sv2v_reg ,
  \nz.mem_969_sv2v_reg ,\nz.mem_968_sv2v_reg ,\nz.mem_967_sv2v_reg ,
  \nz.mem_966_sv2v_reg ,\nz.mem_965_sv2v_reg ,\nz.mem_964_sv2v_reg ,\nz.mem_963_sv2v_reg ,
  \nz.mem_962_sv2v_reg ,\nz.mem_961_sv2v_reg ,\nz.mem_960_sv2v_reg ,\nz.mem_959_sv2v_reg ,
  \nz.mem_958_sv2v_reg ,\nz.mem_957_sv2v_reg ,\nz.mem_956_sv2v_reg ,
  \nz.mem_955_sv2v_reg ,\nz.mem_954_sv2v_reg ,\nz.mem_953_sv2v_reg ,\nz.mem_952_sv2v_reg ,
  \nz.mem_951_sv2v_reg ,\nz.mem_950_sv2v_reg ,\nz.mem_949_sv2v_reg ,\nz.mem_948_sv2v_reg ,
  \nz.mem_947_sv2v_reg ,\nz.mem_946_sv2v_reg ,\nz.mem_945_sv2v_reg ,
  \nz.mem_944_sv2v_reg ,\nz.mem_943_sv2v_reg ,\nz.mem_942_sv2v_reg ,\nz.mem_941_sv2v_reg ,
  \nz.mem_940_sv2v_reg ,\nz.mem_939_sv2v_reg ,\nz.mem_938_sv2v_reg ,
  \nz.mem_937_sv2v_reg ,\nz.mem_936_sv2v_reg ,\nz.mem_935_sv2v_reg ,\nz.mem_934_sv2v_reg ,
  \nz.mem_933_sv2v_reg ,\nz.mem_932_sv2v_reg ,\nz.mem_931_sv2v_reg ,\nz.mem_930_sv2v_reg ,
  \nz.mem_929_sv2v_reg ,\nz.mem_928_sv2v_reg ,\nz.mem_927_sv2v_reg ,
  \nz.mem_926_sv2v_reg ,\nz.mem_925_sv2v_reg ,\nz.mem_924_sv2v_reg ,\nz.mem_923_sv2v_reg ,
  \nz.mem_922_sv2v_reg ,\nz.mem_921_sv2v_reg ,\nz.mem_920_sv2v_reg ,\nz.mem_919_sv2v_reg ,
  \nz.mem_918_sv2v_reg ,\nz.mem_917_sv2v_reg ,\nz.mem_916_sv2v_reg ,
  \nz.mem_915_sv2v_reg ,\nz.mem_914_sv2v_reg ,\nz.mem_913_sv2v_reg ,\nz.mem_912_sv2v_reg ,
  \nz.mem_911_sv2v_reg ,\nz.mem_910_sv2v_reg ,\nz.mem_909_sv2v_reg ,\nz.mem_908_sv2v_reg ,
  \nz.mem_907_sv2v_reg ,\nz.mem_906_sv2v_reg ,\nz.mem_905_sv2v_reg ,
  \nz.mem_904_sv2v_reg ,\nz.mem_903_sv2v_reg ,\nz.mem_902_sv2v_reg ,\nz.mem_901_sv2v_reg ,
  \nz.mem_900_sv2v_reg ,\nz.mem_899_sv2v_reg ,\nz.mem_898_sv2v_reg ,
  \nz.mem_897_sv2v_reg ,\nz.mem_896_sv2v_reg ,\nz.mem_895_sv2v_reg ,\nz.mem_894_sv2v_reg ,
  \nz.mem_893_sv2v_reg ,\nz.mem_892_sv2v_reg ,\nz.mem_891_sv2v_reg ,\nz.mem_890_sv2v_reg ,
  \nz.mem_889_sv2v_reg ,\nz.mem_888_sv2v_reg ,\nz.mem_887_sv2v_reg ,
  \nz.mem_886_sv2v_reg ,\nz.mem_885_sv2v_reg ,\nz.mem_884_sv2v_reg ,\nz.mem_883_sv2v_reg ,
  \nz.mem_882_sv2v_reg ,\nz.mem_881_sv2v_reg ,\nz.mem_880_sv2v_reg ,\nz.mem_879_sv2v_reg ,
  \nz.mem_878_sv2v_reg ,\nz.mem_877_sv2v_reg ,\nz.mem_876_sv2v_reg ,
  \nz.mem_875_sv2v_reg ,\nz.mem_874_sv2v_reg ,\nz.mem_873_sv2v_reg ,\nz.mem_872_sv2v_reg ,
  \nz.mem_871_sv2v_reg ,\nz.mem_870_sv2v_reg ,\nz.mem_869_sv2v_reg ,\nz.mem_868_sv2v_reg ,
  \nz.mem_867_sv2v_reg ,\nz.mem_866_sv2v_reg ,\nz.mem_865_sv2v_reg ,
  \nz.mem_864_sv2v_reg ,\nz.mem_863_sv2v_reg ,\nz.mem_862_sv2v_reg ,\nz.mem_861_sv2v_reg ,
  \nz.mem_860_sv2v_reg ,\nz.mem_859_sv2v_reg ,\nz.mem_858_sv2v_reg ,
  \nz.mem_857_sv2v_reg ,\nz.mem_856_sv2v_reg ,\nz.mem_855_sv2v_reg ,\nz.mem_854_sv2v_reg ,
  \nz.mem_853_sv2v_reg ,\nz.mem_852_sv2v_reg ,\nz.mem_851_sv2v_reg ,\nz.mem_850_sv2v_reg ,
  \nz.mem_849_sv2v_reg ,\nz.mem_848_sv2v_reg ,\nz.mem_847_sv2v_reg ,
  \nz.mem_846_sv2v_reg ,\nz.mem_845_sv2v_reg ,\nz.mem_844_sv2v_reg ,\nz.mem_843_sv2v_reg ,
  \nz.mem_842_sv2v_reg ,\nz.mem_841_sv2v_reg ,\nz.mem_840_sv2v_reg ,\nz.mem_839_sv2v_reg ,
  \nz.mem_838_sv2v_reg ,\nz.mem_837_sv2v_reg ,\nz.mem_836_sv2v_reg ,
  \nz.mem_835_sv2v_reg ,\nz.mem_834_sv2v_reg ,\nz.mem_833_sv2v_reg ,\nz.mem_832_sv2v_reg ,
  \nz.mem_831_sv2v_reg ,\nz.mem_830_sv2v_reg ,\nz.mem_829_sv2v_reg ,\nz.mem_828_sv2v_reg ,
  \nz.mem_827_sv2v_reg ,\nz.mem_826_sv2v_reg ,\nz.mem_825_sv2v_reg ,
  \nz.mem_824_sv2v_reg ,\nz.mem_823_sv2v_reg ,\nz.mem_822_sv2v_reg ,\nz.mem_821_sv2v_reg ,
  \nz.mem_820_sv2v_reg ,\nz.mem_819_sv2v_reg ,\nz.mem_818_sv2v_reg ,
  \nz.mem_817_sv2v_reg ,\nz.mem_816_sv2v_reg ,\nz.mem_815_sv2v_reg ,\nz.mem_814_sv2v_reg ,
  \nz.mem_813_sv2v_reg ,\nz.mem_812_sv2v_reg ,\nz.mem_811_sv2v_reg ,\nz.mem_810_sv2v_reg ,
  \nz.mem_809_sv2v_reg ,\nz.mem_808_sv2v_reg ,\nz.mem_807_sv2v_reg ,
  \nz.mem_806_sv2v_reg ,\nz.mem_805_sv2v_reg ,\nz.mem_804_sv2v_reg ,\nz.mem_803_sv2v_reg ,
  \nz.mem_802_sv2v_reg ,\nz.mem_801_sv2v_reg ,\nz.mem_800_sv2v_reg ,\nz.mem_799_sv2v_reg ,
  \nz.mem_798_sv2v_reg ,\nz.mem_797_sv2v_reg ,\nz.mem_796_sv2v_reg ,
  \nz.mem_795_sv2v_reg ,\nz.mem_794_sv2v_reg ,\nz.mem_793_sv2v_reg ,\nz.mem_792_sv2v_reg ,
  \nz.mem_791_sv2v_reg ,\nz.mem_790_sv2v_reg ,\nz.mem_789_sv2v_reg ,\nz.mem_788_sv2v_reg ,
  \nz.mem_787_sv2v_reg ,\nz.mem_786_sv2v_reg ,\nz.mem_785_sv2v_reg ,
  \nz.mem_784_sv2v_reg ,\nz.mem_783_sv2v_reg ,\nz.mem_782_sv2v_reg ,\nz.mem_781_sv2v_reg ,
  \nz.mem_780_sv2v_reg ,\nz.mem_779_sv2v_reg ,\nz.mem_778_sv2v_reg ,
  \nz.mem_777_sv2v_reg ,\nz.mem_776_sv2v_reg ,\nz.mem_775_sv2v_reg ,\nz.mem_774_sv2v_reg ,
  \nz.mem_773_sv2v_reg ,\nz.mem_772_sv2v_reg ,\nz.mem_771_sv2v_reg ,\nz.mem_770_sv2v_reg ,
  \nz.mem_769_sv2v_reg ,\nz.mem_768_sv2v_reg ,\nz.mem_767_sv2v_reg ,
  \nz.mem_766_sv2v_reg ,\nz.mem_765_sv2v_reg ,\nz.mem_764_sv2v_reg ,\nz.mem_763_sv2v_reg ,
  \nz.mem_762_sv2v_reg ,\nz.mem_761_sv2v_reg ,\nz.mem_760_sv2v_reg ,\nz.mem_759_sv2v_reg ,
  \nz.mem_758_sv2v_reg ,\nz.mem_757_sv2v_reg ,\nz.mem_756_sv2v_reg ,
  \nz.mem_755_sv2v_reg ,\nz.mem_754_sv2v_reg ,\nz.mem_753_sv2v_reg ,\nz.mem_752_sv2v_reg ,
  \nz.mem_751_sv2v_reg ,\nz.mem_750_sv2v_reg ,\nz.mem_749_sv2v_reg ,\nz.mem_748_sv2v_reg ,
  \nz.mem_747_sv2v_reg ,\nz.mem_746_sv2v_reg ,\nz.mem_745_sv2v_reg ,
  \nz.mem_744_sv2v_reg ,\nz.mem_743_sv2v_reg ,\nz.mem_742_sv2v_reg ,\nz.mem_741_sv2v_reg ,
  \nz.mem_740_sv2v_reg ,\nz.mem_739_sv2v_reg ,\nz.mem_738_sv2v_reg ,
  \nz.mem_737_sv2v_reg ,\nz.mem_736_sv2v_reg ,\nz.mem_735_sv2v_reg ,\nz.mem_734_sv2v_reg ,
  \nz.mem_733_sv2v_reg ,\nz.mem_732_sv2v_reg ,\nz.mem_731_sv2v_reg ,\nz.mem_730_sv2v_reg ,
  \nz.mem_729_sv2v_reg ,\nz.mem_728_sv2v_reg ,\nz.mem_727_sv2v_reg ,
  \nz.mem_726_sv2v_reg ,\nz.mem_725_sv2v_reg ,\nz.mem_724_sv2v_reg ,\nz.mem_723_sv2v_reg ,
  \nz.mem_722_sv2v_reg ,\nz.mem_721_sv2v_reg ,\nz.mem_720_sv2v_reg ,\nz.mem_719_sv2v_reg ,
  \nz.mem_718_sv2v_reg ,\nz.mem_717_sv2v_reg ,\nz.mem_716_sv2v_reg ,
  \nz.mem_715_sv2v_reg ,\nz.mem_714_sv2v_reg ,\nz.mem_713_sv2v_reg ,\nz.mem_712_sv2v_reg ,
  \nz.mem_711_sv2v_reg ,\nz.mem_710_sv2v_reg ,\nz.mem_709_sv2v_reg ,\nz.mem_708_sv2v_reg ,
  \nz.mem_707_sv2v_reg ,\nz.mem_706_sv2v_reg ,\nz.mem_705_sv2v_reg ,
  \nz.mem_704_sv2v_reg ,\nz.mem_703_sv2v_reg ,\nz.mem_702_sv2v_reg ,\nz.mem_701_sv2v_reg ,
  \nz.mem_700_sv2v_reg ,\nz.mem_699_sv2v_reg ,\nz.mem_698_sv2v_reg ,
  \nz.mem_697_sv2v_reg ,\nz.mem_696_sv2v_reg ,\nz.mem_695_sv2v_reg ,\nz.mem_694_sv2v_reg ,
  \nz.mem_693_sv2v_reg ,\nz.mem_692_sv2v_reg ,\nz.mem_691_sv2v_reg ,\nz.mem_690_sv2v_reg ,
  \nz.mem_689_sv2v_reg ,\nz.mem_688_sv2v_reg ,\nz.mem_687_sv2v_reg ,
  \nz.mem_686_sv2v_reg ,\nz.mem_685_sv2v_reg ,\nz.mem_684_sv2v_reg ,\nz.mem_683_sv2v_reg ,
  \nz.mem_682_sv2v_reg ,\nz.mem_681_sv2v_reg ,\nz.mem_680_sv2v_reg ,\nz.mem_679_sv2v_reg ,
  \nz.mem_678_sv2v_reg ,\nz.mem_677_sv2v_reg ,\nz.mem_676_sv2v_reg ,
  \nz.mem_675_sv2v_reg ,\nz.mem_674_sv2v_reg ,\nz.mem_673_sv2v_reg ,\nz.mem_672_sv2v_reg ,
  \nz.mem_671_sv2v_reg ,\nz.mem_670_sv2v_reg ,\nz.mem_669_sv2v_reg ,\nz.mem_668_sv2v_reg ,
  \nz.mem_667_sv2v_reg ,\nz.mem_666_sv2v_reg ,\nz.mem_665_sv2v_reg ,
  \nz.mem_664_sv2v_reg ,\nz.mem_663_sv2v_reg ,\nz.mem_662_sv2v_reg ,\nz.mem_661_sv2v_reg ,
  \nz.mem_660_sv2v_reg ,\nz.mem_659_sv2v_reg ,\nz.mem_658_sv2v_reg ,
  \nz.mem_657_sv2v_reg ,\nz.mem_656_sv2v_reg ,\nz.mem_655_sv2v_reg ,\nz.mem_654_sv2v_reg ,
  \nz.mem_653_sv2v_reg ,\nz.mem_652_sv2v_reg ,\nz.mem_651_sv2v_reg ,\nz.mem_650_sv2v_reg ,
  \nz.mem_649_sv2v_reg ,\nz.mem_648_sv2v_reg ,\nz.mem_647_sv2v_reg ,
  \nz.mem_646_sv2v_reg ,\nz.mem_645_sv2v_reg ,\nz.mem_644_sv2v_reg ,\nz.mem_643_sv2v_reg ,
  \nz.mem_642_sv2v_reg ,\nz.mem_641_sv2v_reg ,\nz.mem_640_sv2v_reg ,\nz.mem_639_sv2v_reg ,
  \nz.mem_638_sv2v_reg ,\nz.mem_637_sv2v_reg ,\nz.mem_636_sv2v_reg ,
  \nz.mem_635_sv2v_reg ,\nz.mem_634_sv2v_reg ,\nz.mem_633_sv2v_reg ,\nz.mem_632_sv2v_reg ,
  \nz.mem_631_sv2v_reg ,\nz.mem_630_sv2v_reg ,\nz.mem_629_sv2v_reg ,\nz.mem_628_sv2v_reg ,
  \nz.mem_627_sv2v_reg ,\nz.mem_626_sv2v_reg ,\nz.mem_625_sv2v_reg ,
  \nz.mem_624_sv2v_reg ,\nz.mem_623_sv2v_reg ,\nz.mem_622_sv2v_reg ,\nz.mem_621_sv2v_reg ,
  \nz.mem_620_sv2v_reg ,\nz.mem_619_sv2v_reg ,\nz.mem_618_sv2v_reg ,
  \nz.mem_617_sv2v_reg ,\nz.mem_616_sv2v_reg ,\nz.mem_615_sv2v_reg ,\nz.mem_614_sv2v_reg ,
  \nz.mem_613_sv2v_reg ,\nz.mem_612_sv2v_reg ,\nz.mem_611_sv2v_reg ,\nz.mem_610_sv2v_reg ,
  \nz.mem_609_sv2v_reg ,\nz.mem_608_sv2v_reg ,\nz.mem_607_sv2v_reg ,
  \nz.mem_606_sv2v_reg ,\nz.mem_605_sv2v_reg ,\nz.mem_604_sv2v_reg ,\nz.mem_603_sv2v_reg ,
  \nz.mem_602_sv2v_reg ,\nz.mem_601_sv2v_reg ,\nz.mem_600_sv2v_reg ,\nz.mem_599_sv2v_reg ,
  \nz.mem_598_sv2v_reg ,\nz.mem_597_sv2v_reg ,\nz.mem_596_sv2v_reg ,
  \nz.mem_595_sv2v_reg ,\nz.mem_594_sv2v_reg ,\nz.mem_593_sv2v_reg ,\nz.mem_592_sv2v_reg ,
  \nz.mem_591_sv2v_reg ,\nz.mem_590_sv2v_reg ,\nz.mem_589_sv2v_reg ,\nz.mem_588_sv2v_reg ,
  \nz.mem_587_sv2v_reg ,\nz.mem_586_sv2v_reg ,\nz.mem_585_sv2v_reg ,
  \nz.mem_584_sv2v_reg ,\nz.mem_583_sv2v_reg ,\nz.mem_582_sv2v_reg ,\nz.mem_581_sv2v_reg ,
  \nz.mem_580_sv2v_reg ,\nz.mem_579_sv2v_reg ,\nz.mem_578_sv2v_reg ,
  \nz.mem_577_sv2v_reg ,\nz.mem_576_sv2v_reg ,\nz.mem_575_sv2v_reg ,\nz.mem_574_sv2v_reg ,
  \nz.mem_573_sv2v_reg ,\nz.mem_572_sv2v_reg ,\nz.mem_571_sv2v_reg ,\nz.mem_570_sv2v_reg ,
  \nz.mem_569_sv2v_reg ,\nz.mem_568_sv2v_reg ,\nz.mem_567_sv2v_reg ,
  \nz.mem_566_sv2v_reg ,\nz.mem_565_sv2v_reg ,\nz.mem_564_sv2v_reg ,\nz.mem_563_sv2v_reg ,
  \nz.mem_562_sv2v_reg ,\nz.mem_561_sv2v_reg ,\nz.mem_560_sv2v_reg ,\nz.mem_559_sv2v_reg ,
  \nz.mem_558_sv2v_reg ,\nz.mem_557_sv2v_reg ,\nz.mem_556_sv2v_reg ,
  \nz.mem_555_sv2v_reg ,\nz.mem_554_sv2v_reg ,\nz.mem_553_sv2v_reg ,\nz.mem_552_sv2v_reg ,
  \nz.mem_551_sv2v_reg ,\nz.mem_550_sv2v_reg ,\nz.mem_549_sv2v_reg ,\nz.mem_548_sv2v_reg ,
  \nz.mem_547_sv2v_reg ,\nz.mem_546_sv2v_reg ,\nz.mem_545_sv2v_reg ,
  \nz.mem_544_sv2v_reg ,\nz.mem_543_sv2v_reg ,\nz.mem_542_sv2v_reg ,\nz.mem_541_sv2v_reg ,
  \nz.mem_540_sv2v_reg ,\nz.mem_539_sv2v_reg ,\nz.mem_538_sv2v_reg ,
  \nz.mem_537_sv2v_reg ,\nz.mem_536_sv2v_reg ,\nz.mem_535_sv2v_reg ,\nz.mem_534_sv2v_reg ,
  \nz.mem_533_sv2v_reg ,\nz.mem_532_sv2v_reg ,\nz.mem_531_sv2v_reg ,\nz.mem_530_sv2v_reg ,
  \nz.mem_529_sv2v_reg ,\nz.mem_528_sv2v_reg ,\nz.mem_527_sv2v_reg ,
  \nz.mem_526_sv2v_reg ,\nz.mem_525_sv2v_reg ,\nz.mem_524_sv2v_reg ,\nz.mem_523_sv2v_reg ,
  \nz.mem_522_sv2v_reg ,\nz.mem_521_sv2v_reg ,\nz.mem_520_sv2v_reg ,\nz.mem_519_sv2v_reg ,
  \nz.mem_518_sv2v_reg ,\nz.mem_517_sv2v_reg ,\nz.mem_516_sv2v_reg ,
  \nz.mem_515_sv2v_reg ,\nz.mem_514_sv2v_reg ,\nz.mem_513_sv2v_reg ,\nz.mem_512_sv2v_reg ,
  \nz.mem_511_sv2v_reg ,\nz.mem_510_sv2v_reg ,\nz.mem_509_sv2v_reg ,\nz.mem_508_sv2v_reg ,
  \nz.mem_507_sv2v_reg ,\nz.mem_506_sv2v_reg ,\nz.mem_505_sv2v_reg ,
  \nz.mem_504_sv2v_reg ,\nz.mem_503_sv2v_reg ,\nz.mem_502_sv2v_reg ,\nz.mem_501_sv2v_reg ,
  \nz.mem_500_sv2v_reg ,\nz.mem_499_sv2v_reg ,\nz.mem_498_sv2v_reg ,
  \nz.mem_497_sv2v_reg ,\nz.mem_496_sv2v_reg ,\nz.mem_495_sv2v_reg ,\nz.mem_494_sv2v_reg ,
  \nz.mem_493_sv2v_reg ,\nz.mem_492_sv2v_reg ,\nz.mem_491_sv2v_reg ,\nz.mem_490_sv2v_reg ,
  \nz.mem_489_sv2v_reg ,\nz.mem_488_sv2v_reg ,\nz.mem_487_sv2v_reg ,
  \nz.mem_486_sv2v_reg ,\nz.mem_485_sv2v_reg ,\nz.mem_484_sv2v_reg ,\nz.mem_483_sv2v_reg ,
  \nz.mem_482_sv2v_reg ,\nz.mem_481_sv2v_reg ,\nz.mem_480_sv2v_reg ,\nz.mem_479_sv2v_reg ,
  \nz.mem_478_sv2v_reg ,\nz.mem_477_sv2v_reg ,\nz.mem_476_sv2v_reg ,
  \nz.mem_475_sv2v_reg ,\nz.mem_474_sv2v_reg ,\nz.mem_473_sv2v_reg ,\nz.mem_472_sv2v_reg ,
  \nz.mem_471_sv2v_reg ,\nz.mem_470_sv2v_reg ,\nz.mem_469_sv2v_reg ,\nz.mem_468_sv2v_reg ,
  \nz.mem_467_sv2v_reg ,\nz.mem_466_sv2v_reg ,\nz.mem_465_sv2v_reg ,
  \nz.mem_464_sv2v_reg ,\nz.mem_463_sv2v_reg ,\nz.mem_462_sv2v_reg ,\nz.mem_461_sv2v_reg ,
  \nz.mem_460_sv2v_reg ,\nz.mem_459_sv2v_reg ,\nz.mem_458_sv2v_reg ,
  \nz.mem_457_sv2v_reg ,\nz.mem_456_sv2v_reg ,\nz.mem_455_sv2v_reg ,\nz.mem_454_sv2v_reg ,
  \nz.mem_453_sv2v_reg ,\nz.mem_452_sv2v_reg ,\nz.mem_451_sv2v_reg ,\nz.mem_450_sv2v_reg ,
  \nz.mem_449_sv2v_reg ,\nz.mem_448_sv2v_reg ,\nz.mem_447_sv2v_reg ,
  \nz.mem_446_sv2v_reg ,\nz.mem_445_sv2v_reg ,\nz.mem_444_sv2v_reg ,\nz.mem_443_sv2v_reg ,
  \nz.mem_442_sv2v_reg ,\nz.mem_441_sv2v_reg ,\nz.mem_440_sv2v_reg ,\nz.mem_439_sv2v_reg ,
  \nz.mem_438_sv2v_reg ,\nz.mem_437_sv2v_reg ,\nz.mem_436_sv2v_reg ,
  \nz.mem_435_sv2v_reg ,\nz.mem_434_sv2v_reg ,\nz.mem_433_sv2v_reg ,\nz.mem_432_sv2v_reg ,
  \nz.mem_431_sv2v_reg ,\nz.mem_430_sv2v_reg ,\nz.mem_429_sv2v_reg ,\nz.mem_428_sv2v_reg ,
  \nz.mem_427_sv2v_reg ,\nz.mem_426_sv2v_reg ,\nz.mem_425_sv2v_reg ,
  \nz.mem_424_sv2v_reg ,\nz.mem_423_sv2v_reg ,\nz.mem_422_sv2v_reg ,\nz.mem_421_sv2v_reg ,
  \nz.mem_420_sv2v_reg ,\nz.mem_419_sv2v_reg ,\nz.mem_418_sv2v_reg ,
  \nz.mem_417_sv2v_reg ,\nz.mem_416_sv2v_reg ,\nz.mem_415_sv2v_reg ,\nz.mem_414_sv2v_reg ,
  \nz.mem_413_sv2v_reg ,\nz.mem_412_sv2v_reg ,\nz.mem_411_sv2v_reg ,\nz.mem_410_sv2v_reg ,
  \nz.mem_409_sv2v_reg ,\nz.mem_408_sv2v_reg ,\nz.mem_407_sv2v_reg ,
  \nz.mem_406_sv2v_reg ,\nz.mem_405_sv2v_reg ,\nz.mem_404_sv2v_reg ,\nz.mem_403_sv2v_reg ,
  \nz.mem_402_sv2v_reg ,\nz.mem_401_sv2v_reg ,\nz.mem_400_sv2v_reg ,\nz.mem_399_sv2v_reg ,
  \nz.mem_398_sv2v_reg ,\nz.mem_397_sv2v_reg ,\nz.mem_396_sv2v_reg ,
  \nz.mem_395_sv2v_reg ,\nz.mem_394_sv2v_reg ,\nz.mem_393_sv2v_reg ,\nz.mem_392_sv2v_reg ,
  \nz.mem_391_sv2v_reg ,\nz.mem_390_sv2v_reg ,\nz.mem_389_sv2v_reg ,\nz.mem_388_sv2v_reg ,
  \nz.mem_387_sv2v_reg ,\nz.mem_386_sv2v_reg ,\nz.mem_385_sv2v_reg ,
  \nz.mem_384_sv2v_reg ,\nz.mem_383_sv2v_reg ,\nz.mem_382_sv2v_reg ,\nz.mem_381_sv2v_reg ,
  \nz.mem_380_sv2v_reg ,\nz.mem_379_sv2v_reg ,\nz.mem_378_sv2v_reg ,
  \nz.mem_377_sv2v_reg ,\nz.mem_376_sv2v_reg ,\nz.mem_375_sv2v_reg ,\nz.mem_374_sv2v_reg ,
  \nz.mem_373_sv2v_reg ,\nz.mem_372_sv2v_reg ,\nz.mem_371_sv2v_reg ,\nz.mem_370_sv2v_reg ,
  \nz.mem_369_sv2v_reg ,\nz.mem_368_sv2v_reg ,\nz.mem_367_sv2v_reg ,
  \nz.mem_366_sv2v_reg ,\nz.mem_365_sv2v_reg ,\nz.mem_364_sv2v_reg ,\nz.mem_363_sv2v_reg ,
  \nz.mem_362_sv2v_reg ,\nz.mem_361_sv2v_reg ,\nz.mem_360_sv2v_reg ,\nz.mem_359_sv2v_reg ,
  \nz.mem_358_sv2v_reg ,\nz.mem_357_sv2v_reg ,\nz.mem_356_sv2v_reg ,
  \nz.mem_355_sv2v_reg ,\nz.mem_354_sv2v_reg ,\nz.mem_353_sv2v_reg ,\nz.mem_352_sv2v_reg ,
  \nz.mem_351_sv2v_reg ,\nz.mem_350_sv2v_reg ,\nz.mem_349_sv2v_reg ,\nz.mem_348_sv2v_reg ,
  \nz.mem_347_sv2v_reg ,\nz.mem_346_sv2v_reg ,\nz.mem_345_sv2v_reg ,
  \nz.mem_344_sv2v_reg ,\nz.mem_343_sv2v_reg ,\nz.mem_342_sv2v_reg ,\nz.mem_341_sv2v_reg ,
  \nz.mem_340_sv2v_reg ,\nz.mem_339_sv2v_reg ,\nz.mem_338_sv2v_reg ,
  \nz.mem_337_sv2v_reg ,\nz.mem_336_sv2v_reg ,\nz.mem_335_sv2v_reg ,\nz.mem_334_sv2v_reg ,
  \nz.mem_333_sv2v_reg ,\nz.mem_332_sv2v_reg ,\nz.mem_331_sv2v_reg ,\nz.mem_330_sv2v_reg ,
  \nz.mem_329_sv2v_reg ,\nz.mem_328_sv2v_reg ,\nz.mem_327_sv2v_reg ,
  \nz.mem_326_sv2v_reg ,\nz.mem_325_sv2v_reg ,\nz.mem_324_sv2v_reg ,\nz.mem_323_sv2v_reg ,
  \nz.mem_322_sv2v_reg ,\nz.mem_321_sv2v_reg ,\nz.mem_320_sv2v_reg ,\nz.mem_319_sv2v_reg ,
  \nz.mem_318_sv2v_reg ,\nz.mem_317_sv2v_reg ,\nz.mem_316_sv2v_reg ,
  \nz.mem_315_sv2v_reg ,\nz.mem_314_sv2v_reg ,\nz.mem_313_sv2v_reg ,\nz.mem_312_sv2v_reg ,
  \nz.mem_311_sv2v_reg ,\nz.mem_310_sv2v_reg ,\nz.mem_309_sv2v_reg ,\nz.mem_308_sv2v_reg ,
  \nz.mem_307_sv2v_reg ,\nz.mem_306_sv2v_reg ,\nz.mem_305_sv2v_reg ,
  \nz.mem_304_sv2v_reg ,\nz.mem_303_sv2v_reg ,\nz.mem_302_sv2v_reg ,\nz.mem_301_sv2v_reg ,
  \nz.mem_300_sv2v_reg ,\nz.mem_299_sv2v_reg ,\nz.mem_298_sv2v_reg ,
  \nz.mem_297_sv2v_reg ,\nz.mem_296_sv2v_reg ,\nz.mem_295_sv2v_reg ,\nz.mem_294_sv2v_reg ,
  \nz.mem_293_sv2v_reg ,\nz.mem_292_sv2v_reg ,\nz.mem_291_sv2v_reg ,\nz.mem_290_sv2v_reg ,
  \nz.mem_289_sv2v_reg ,\nz.mem_288_sv2v_reg ,\nz.mem_287_sv2v_reg ,
  \nz.mem_286_sv2v_reg ,\nz.mem_285_sv2v_reg ,\nz.mem_284_sv2v_reg ,\nz.mem_283_sv2v_reg ,
  \nz.mem_282_sv2v_reg ,\nz.mem_281_sv2v_reg ,\nz.mem_280_sv2v_reg ,\nz.mem_279_sv2v_reg ,
  \nz.mem_278_sv2v_reg ,\nz.mem_277_sv2v_reg ,\nz.mem_276_sv2v_reg ,
  \nz.mem_275_sv2v_reg ,\nz.mem_274_sv2v_reg ,\nz.mem_273_sv2v_reg ,\nz.mem_272_sv2v_reg ,
  \nz.mem_271_sv2v_reg ,\nz.mem_270_sv2v_reg ,\nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,
  \nz.mem_267_sv2v_reg ,\nz.mem_266_sv2v_reg ,\nz.mem_265_sv2v_reg ,
  \nz.mem_264_sv2v_reg ,\nz.mem_263_sv2v_reg ,\nz.mem_262_sv2v_reg ,\nz.mem_261_sv2v_reg ,
  \nz.mem_260_sv2v_reg ,\nz.mem_259_sv2v_reg ,\nz.mem_258_sv2v_reg ,
  \nz.mem_257_sv2v_reg ,\nz.mem_256_sv2v_reg ,\nz.mem_255_sv2v_reg ,\nz.mem_254_sv2v_reg ,
  \nz.mem_253_sv2v_reg ,\nz.mem_252_sv2v_reg ,\nz.mem_251_sv2v_reg ,\nz.mem_250_sv2v_reg ,
  \nz.mem_249_sv2v_reg ,\nz.mem_248_sv2v_reg ,\nz.mem_247_sv2v_reg ,
  \nz.mem_246_sv2v_reg ,\nz.mem_245_sv2v_reg ,\nz.mem_244_sv2v_reg ,\nz.mem_243_sv2v_reg ,
  \nz.mem_242_sv2v_reg ,\nz.mem_241_sv2v_reg ,\nz.mem_240_sv2v_reg ,\nz.mem_239_sv2v_reg ,
  \nz.mem_238_sv2v_reg ,\nz.mem_237_sv2v_reg ,\nz.mem_236_sv2v_reg ,
  \nz.mem_235_sv2v_reg ,\nz.mem_234_sv2v_reg ,\nz.mem_233_sv2v_reg ,\nz.mem_232_sv2v_reg ,
  \nz.mem_231_sv2v_reg ,\nz.mem_230_sv2v_reg ,\nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,
  \nz.mem_227_sv2v_reg ,\nz.mem_226_sv2v_reg ,\nz.mem_225_sv2v_reg ,
  \nz.mem_224_sv2v_reg ,\nz.mem_223_sv2v_reg ,\nz.mem_222_sv2v_reg ,\nz.mem_221_sv2v_reg ,
  \nz.mem_220_sv2v_reg ,\nz.mem_219_sv2v_reg ,\nz.mem_218_sv2v_reg ,
  \nz.mem_217_sv2v_reg ,\nz.mem_216_sv2v_reg ,\nz.mem_215_sv2v_reg ,\nz.mem_214_sv2v_reg ,
  \nz.mem_213_sv2v_reg ,\nz.mem_212_sv2v_reg ,\nz.mem_211_sv2v_reg ,\nz.mem_210_sv2v_reg ,
  \nz.mem_209_sv2v_reg ,\nz.mem_208_sv2v_reg ,\nz.mem_207_sv2v_reg ,
  \nz.mem_206_sv2v_reg ,\nz.mem_205_sv2v_reg ,\nz.mem_204_sv2v_reg ,\nz.mem_203_sv2v_reg ,
  \nz.mem_202_sv2v_reg ,\nz.mem_201_sv2v_reg ,\nz.mem_200_sv2v_reg ,\nz.mem_199_sv2v_reg ,
  \nz.mem_198_sv2v_reg ,\nz.mem_197_sv2v_reg ,\nz.mem_196_sv2v_reg ,
  \nz.mem_195_sv2v_reg ,\nz.mem_194_sv2v_reg ,\nz.mem_193_sv2v_reg ,\nz.mem_192_sv2v_reg ,
  \nz.mem_191_sv2v_reg ,\nz.mem_190_sv2v_reg ,\nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,
  \nz.mem_187_sv2v_reg ,\nz.mem_186_sv2v_reg ,\nz.mem_185_sv2v_reg ,
  \nz.mem_184_sv2v_reg ,\nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,\nz.mem_181_sv2v_reg ,
  \nz.mem_180_sv2v_reg ,\nz.mem_179_sv2v_reg ,\nz.mem_178_sv2v_reg ,
  \nz.mem_177_sv2v_reg ,\nz.mem_176_sv2v_reg ,\nz.mem_175_sv2v_reg ,\nz.mem_174_sv2v_reg ,
  \nz.mem_173_sv2v_reg ,\nz.mem_172_sv2v_reg ,\nz.mem_171_sv2v_reg ,\nz.mem_170_sv2v_reg ,
  \nz.mem_169_sv2v_reg ,\nz.mem_168_sv2v_reg ,\nz.mem_167_sv2v_reg ,
  \nz.mem_166_sv2v_reg ,\nz.mem_165_sv2v_reg ,\nz.mem_164_sv2v_reg ,\nz.mem_163_sv2v_reg ,
  \nz.mem_162_sv2v_reg ,\nz.mem_161_sv2v_reg ,\nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,
  \nz.mem_158_sv2v_reg ,\nz.mem_157_sv2v_reg ,\nz.mem_156_sv2v_reg ,
  \nz.mem_155_sv2v_reg ,\nz.mem_154_sv2v_reg ,\nz.mem_153_sv2v_reg ,\nz.mem_152_sv2v_reg ,
  \nz.mem_151_sv2v_reg ,\nz.mem_150_sv2v_reg ,\nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,
  \nz.mem_147_sv2v_reg ,\nz.mem_146_sv2v_reg ,\nz.mem_145_sv2v_reg ,
  \nz.mem_144_sv2v_reg ,\nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,\nz.mem_141_sv2v_reg ,
  \nz.mem_140_sv2v_reg ,\nz.mem_139_sv2v_reg ,\nz.mem_138_sv2v_reg ,
  \nz.mem_137_sv2v_reg ,\nz.mem_136_sv2v_reg ,\nz.mem_135_sv2v_reg ,\nz.mem_134_sv2v_reg ,
  \nz.mem_133_sv2v_reg ,\nz.mem_132_sv2v_reg ,\nz.mem_131_sv2v_reg ,\nz.mem_130_sv2v_reg ,
  \nz.mem_129_sv2v_reg ,\nz.mem_128_sv2v_reg ,\nz.mem_127_sv2v_reg ,
  \nz.mem_126_sv2v_reg ,\nz.mem_125_sv2v_reg ,\nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,
  \nz.mem_122_sv2v_reg ,\nz.mem_121_sv2v_reg ,\nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,
  \nz.mem_118_sv2v_reg ,\nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,
  \nz.mem_115_sv2v_reg ,\nz.mem_114_sv2v_reg ,\nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,
  \nz.mem_111_sv2v_reg ,\nz.mem_110_sv2v_reg ,\nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,
  \nz.mem_107_sv2v_reg ,\nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,
  \nz.mem_104_sv2v_reg ,\nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,
  \nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,\nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,
  \nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,
  \nz.mem_93_sv2v_reg ,\nz.mem_92_sv2v_reg ,\nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,
  \nz.mem_89_sv2v_reg ,\nz.mem_88_sv2v_reg ,\nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,
  \nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,\nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,
  \nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,\nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,
  \nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,\nz.mem_75_sv2v_reg ,
  \nz.mem_74_sv2v_reg ,\nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,
  \nz.mem_70_sv2v_reg ,\nz.mem_69_sv2v_reg ,\nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,
  \nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,
  \nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,\nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,
  \nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,\nz.mem_56_sv2v_reg ,
  \nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,
  \nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,
  \nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,
  \nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,\nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,
  \nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,\nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,
  \nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,
  \nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,
  \nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,
  \nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,\nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,
  \nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,\nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,
  \nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,
  \nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,
  \nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,
  \nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,
  \nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.mem [1391] = \nz.mem_1391_sv2v_reg ;
  assign \nz.mem [1390] = \nz.mem_1390_sv2v_reg ;
  assign \nz.mem [1389] = \nz.mem_1389_sv2v_reg ;
  assign \nz.mem [1388] = \nz.mem_1388_sv2v_reg ;
  assign \nz.mem [1387] = \nz.mem_1387_sv2v_reg ;
  assign \nz.mem [1386] = \nz.mem_1386_sv2v_reg ;
  assign \nz.mem [1385] = \nz.mem_1385_sv2v_reg ;
  assign \nz.mem [1384] = \nz.mem_1384_sv2v_reg ;
  assign \nz.mem [1383] = \nz.mem_1383_sv2v_reg ;
  assign \nz.mem [1382] = \nz.mem_1382_sv2v_reg ;
  assign \nz.mem [1381] = \nz.mem_1381_sv2v_reg ;
  assign \nz.mem [1380] = \nz.mem_1380_sv2v_reg ;
  assign \nz.mem [1379] = \nz.mem_1379_sv2v_reg ;
  assign \nz.mem [1378] = \nz.mem_1378_sv2v_reg ;
  assign \nz.mem [1377] = \nz.mem_1377_sv2v_reg ;
  assign \nz.mem [1376] = \nz.mem_1376_sv2v_reg ;
  assign \nz.mem [1375] = \nz.mem_1375_sv2v_reg ;
  assign \nz.mem [1374] = \nz.mem_1374_sv2v_reg ;
  assign \nz.mem [1373] = \nz.mem_1373_sv2v_reg ;
  assign \nz.mem [1372] = \nz.mem_1372_sv2v_reg ;
  assign \nz.mem [1371] = \nz.mem_1371_sv2v_reg ;
  assign \nz.mem [1370] = \nz.mem_1370_sv2v_reg ;
  assign \nz.mem [1369] = \nz.mem_1369_sv2v_reg ;
  assign \nz.mem [1368] = \nz.mem_1368_sv2v_reg ;
  assign \nz.mem [1367] = \nz.mem_1367_sv2v_reg ;
  assign \nz.mem [1366] = \nz.mem_1366_sv2v_reg ;
  assign \nz.mem [1365] = \nz.mem_1365_sv2v_reg ;
  assign \nz.mem [1364] = \nz.mem_1364_sv2v_reg ;
  assign \nz.mem [1363] = \nz.mem_1363_sv2v_reg ;
  assign \nz.mem [1362] = \nz.mem_1362_sv2v_reg ;
  assign \nz.mem [1361] = \nz.mem_1361_sv2v_reg ;
  assign \nz.mem [1360] = \nz.mem_1360_sv2v_reg ;
  assign \nz.mem [1359] = \nz.mem_1359_sv2v_reg ;
  assign \nz.mem [1358] = \nz.mem_1358_sv2v_reg ;
  assign \nz.mem [1357] = \nz.mem_1357_sv2v_reg ;
  assign \nz.mem [1356] = \nz.mem_1356_sv2v_reg ;
  assign \nz.mem [1355] = \nz.mem_1355_sv2v_reg ;
  assign \nz.mem [1354] = \nz.mem_1354_sv2v_reg ;
  assign \nz.mem [1353] = \nz.mem_1353_sv2v_reg ;
  assign \nz.mem [1352] = \nz.mem_1352_sv2v_reg ;
  assign \nz.mem [1351] = \nz.mem_1351_sv2v_reg ;
  assign \nz.mem [1350] = \nz.mem_1350_sv2v_reg ;
  assign \nz.mem [1349] = \nz.mem_1349_sv2v_reg ;
  assign \nz.mem [1348] = \nz.mem_1348_sv2v_reg ;
  assign \nz.mem [1347] = \nz.mem_1347_sv2v_reg ;
  assign \nz.mem [1346] = \nz.mem_1346_sv2v_reg ;
  assign \nz.mem [1345] = \nz.mem_1345_sv2v_reg ;
  assign \nz.mem [1344] = \nz.mem_1344_sv2v_reg ;
  assign \nz.mem [1343] = \nz.mem_1343_sv2v_reg ;
  assign \nz.mem [1342] = \nz.mem_1342_sv2v_reg ;
  assign \nz.mem [1341] = \nz.mem_1341_sv2v_reg ;
  assign \nz.mem [1340] = \nz.mem_1340_sv2v_reg ;
  assign \nz.mem [1339] = \nz.mem_1339_sv2v_reg ;
  assign \nz.mem [1338] = \nz.mem_1338_sv2v_reg ;
  assign \nz.mem [1337] = \nz.mem_1337_sv2v_reg ;
  assign \nz.mem [1336] = \nz.mem_1336_sv2v_reg ;
  assign \nz.mem [1335] = \nz.mem_1335_sv2v_reg ;
  assign \nz.mem [1334] = \nz.mem_1334_sv2v_reg ;
  assign \nz.mem [1333] = \nz.mem_1333_sv2v_reg ;
  assign \nz.mem [1332] = \nz.mem_1332_sv2v_reg ;
  assign \nz.mem [1331] = \nz.mem_1331_sv2v_reg ;
  assign \nz.mem [1330] = \nz.mem_1330_sv2v_reg ;
  assign \nz.mem [1329] = \nz.mem_1329_sv2v_reg ;
  assign \nz.mem [1328] = \nz.mem_1328_sv2v_reg ;
  assign \nz.mem [1327] = \nz.mem_1327_sv2v_reg ;
  assign \nz.mem [1326] = \nz.mem_1326_sv2v_reg ;
  assign \nz.mem [1325] = \nz.mem_1325_sv2v_reg ;
  assign \nz.mem [1324] = \nz.mem_1324_sv2v_reg ;
  assign \nz.mem [1323] = \nz.mem_1323_sv2v_reg ;
  assign \nz.mem [1322] = \nz.mem_1322_sv2v_reg ;
  assign \nz.mem [1321] = \nz.mem_1321_sv2v_reg ;
  assign \nz.mem [1320] = \nz.mem_1320_sv2v_reg ;
  assign \nz.mem [1319] = \nz.mem_1319_sv2v_reg ;
  assign \nz.mem [1318] = \nz.mem_1318_sv2v_reg ;
  assign \nz.mem [1317] = \nz.mem_1317_sv2v_reg ;
  assign \nz.mem [1316] = \nz.mem_1316_sv2v_reg ;
  assign \nz.mem [1315] = \nz.mem_1315_sv2v_reg ;
  assign \nz.mem [1314] = \nz.mem_1314_sv2v_reg ;
  assign \nz.mem [1313] = \nz.mem_1313_sv2v_reg ;
  assign \nz.mem [1312] = \nz.mem_1312_sv2v_reg ;
  assign \nz.mem [1311] = \nz.mem_1311_sv2v_reg ;
  assign \nz.mem [1310] = \nz.mem_1310_sv2v_reg ;
  assign \nz.mem [1309] = \nz.mem_1309_sv2v_reg ;
  assign \nz.mem [1308] = \nz.mem_1308_sv2v_reg ;
  assign \nz.mem [1307] = \nz.mem_1307_sv2v_reg ;
  assign \nz.mem [1306] = \nz.mem_1306_sv2v_reg ;
  assign \nz.mem [1305] = \nz.mem_1305_sv2v_reg ;
  assign \nz.mem [1304] = \nz.mem_1304_sv2v_reg ;
  assign \nz.mem [1303] = \nz.mem_1303_sv2v_reg ;
  assign \nz.mem [1302] = \nz.mem_1302_sv2v_reg ;
  assign \nz.mem [1301] = \nz.mem_1301_sv2v_reg ;
  assign \nz.mem [1300] = \nz.mem_1300_sv2v_reg ;
  assign \nz.mem [1299] = \nz.mem_1299_sv2v_reg ;
  assign \nz.mem [1298] = \nz.mem_1298_sv2v_reg ;
  assign \nz.mem [1297] = \nz.mem_1297_sv2v_reg ;
  assign \nz.mem [1296] = \nz.mem_1296_sv2v_reg ;
  assign \nz.mem [1295] = \nz.mem_1295_sv2v_reg ;
  assign \nz.mem [1294] = \nz.mem_1294_sv2v_reg ;
  assign \nz.mem [1293] = \nz.mem_1293_sv2v_reg ;
  assign \nz.mem [1292] = \nz.mem_1292_sv2v_reg ;
  assign \nz.mem [1291] = \nz.mem_1291_sv2v_reg ;
  assign \nz.mem [1290] = \nz.mem_1290_sv2v_reg ;
  assign \nz.mem [1289] = \nz.mem_1289_sv2v_reg ;
  assign \nz.mem [1288] = \nz.mem_1288_sv2v_reg ;
  assign \nz.mem [1287] = \nz.mem_1287_sv2v_reg ;
  assign \nz.mem [1286] = \nz.mem_1286_sv2v_reg ;
  assign \nz.mem [1285] = \nz.mem_1285_sv2v_reg ;
  assign \nz.mem [1284] = \nz.mem_1284_sv2v_reg ;
  assign \nz.mem [1283] = \nz.mem_1283_sv2v_reg ;
  assign \nz.mem [1282] = \nz.mem_1282_sv2v_reg ;
  assign \nz.mem [1281] = \nz.mem_1281_sv2v_reg ;
  assign \nz.mem [1280] = \nz.mem_1280_sv2v_reg ;
  assign \nz.mem [1279] = \nz.mem_1279_sv2v_reg ;
  assign \nz.mem [1278] = \nz.mem_1278_sv2v_reg ;
  assign \nz.mem [1277] = \nz.mem_1277_sv2v_reg ;
  assign \nz.mem [1276] = \nz.mem_1276_sv2v_reg ;
  assign \nz.mem [1275] = \nz.mem_1275_sv2v_reg ;
  assign \nz.mem [1274] = \nz.mem_1274_sv2v_reg ;
  assign \nz.mem [1273] = \nz.mem_1273_sv2v_reg ;
  assign \nz.mem [1272] = \nz.mem_1272_sv2v_reg ;
  assign \nz.mem [1271] = \nz.mem_1271_sv2v_reg ;
  assign \nz.mem [1270] = \nz.mem_1270_sv2v_reg ;
  assign \nz.mem [1269] = \nz.mem_1269_sv2v_reg ;
  assign \nz.mem [1268] = \nz.mem_1268_sv2v_reg ;
  assign \nz.mem [1267] = \nz.mem_1267_sv2v_reg ;
  assign \nz.mem [1266] = \nz.mem_1266_sv2v_reg ;
  assign \nz.mem [1265] = \nz.mem_1265_sv2v_reg ;
  assign \nz.mem [1264] = \nz.mem_1264_sv2v_reg ;
  assign \nz.mem [1263] = \nz.mem_1263_sv2v_reg ;
  assign \nz.mem [1262] = \nz.mem_1262_sv2v_reg ;
  assign \nz.mem [1261] = \nz.mem_1261_sv2v_reg ;
  assign \nz.mem [1260] = \nz.mem_1260_sv2v_reg ;
  assign \nz.mem [1259] = \nz.mem_1259_sv2v_reg ;
  assign \nz.mem [1258] = \nz.mem_1258_sv2v_reg ;
  assign \nz.mem [1257] = \nz.mem_1257_sv2v_reg ;
  assign \nz.mem [1256] = \nz.mem_1256_sv2v_reg ;
  assign \nz.mem [1255] = \nz.mem_1255_sv2v_reg ;
  assign \nz.mem [1254] = \nz.mem_1254_sv2v_reg ;
  assign \nz.mem [1253] = \nz.mem_1253_sv2v_reg ;
  assign \nz.mem [1252] = \nz.mem_1252_sv2v_reg ;
  assign \nz.mem [1251] = \nz.mem_1251_sv2v_reg ;
  assign \nz.mem [1250] = \nz.mem_1250_sv2v_reg ;
  assign \nz.mem [1249] = \nz.mem_1249_sv2v_reg ;
  assign \nz.mem [1248] = \nz.mem_1248_sv2v_reg ;
  assign \nz.mem [1247] = \nz.mem_1247_sv2v_reg ;
  assign \nz.mem [1246] = \nz.mem_1246_sv2v_reg ;
  assign \nz.mem [1245] = \nz.mem_1245_sv2v_reg ;
  assign \nz.mem [1244] = \nz.mem_1244_sv2v_reg ;
  assign \nz.mem [1243] = \nz.mem_1243_sv2v_reg ;
  assign \nz.mem [1242] = \nz.mem_1242_sv2v_reg ;
  assign \nz.mem [1241] = \nz.mem_1241_sv2v_reg ;
  assign \nz.mem [1240] = \nz.mem_1240_sv2v_reg ;
  assign \nz.mem [1239] = \nz.mem_1239_sv2v_reg ;
  assign \nz.mem [1238] = \nz.mem_1238_sv2v_reg ;
  assign \nz.mem [1237] = \nz.mem_1237_sv2v_reg ;
  assign \nz.mem [1236] = \nz.mem_1236_sv2v_reg ;
  assign \nz.mem [1235] = \nz.mem_1235_sv2v_reg ;
  assign \nz.mem [1234] = \nz.mem_1234_sv2v_reg ;
  assign \nz.mem [1233] = \nz.mem_1233_sv2v_reg ;
  assign \nz.mem [1232] = \nz.mem_1232_sv2v_reg ;
  assign \nz.mem [1231] = \nz.mem_1231_sv2v_reg ;
  assign \nz.mem [1230] = \nz.mem_1230_sv2v_reg ;
  assign \nz.mem [1229] = \nz.mem_1229_sv2v_reg ;
  assign \nz.mem [1228] = \nz.mem_1228_sv2v_reg ;
  assign \nz.mem [1227] = \nz.mem_1227_sv2v_reg ;
  assign \nz.mem [1226] = \nz.mem_1226_sv2v_reg ;
  assign \nz.mem [1225] = \nz.mem_1225_sv2v_reg ;
  assign \nz.mem [1224] = \nz.mem_1224_sv2v_reg ;
  assign \nz.mem [1223] = \nz.mem_1223_sv2v_reg ;
  assign \nz.mem [1222] = \nz.mem_1222_sv2v_reg ;
  assign \nz.mem [1221] = \nz.mem_1221_sv2v_reg ;
  assign \nz.mem [1220] = \nz.mem_1220_sv2v_reg ;
  assign \nz.mem [1219] = \nz.mem_1219_sv2v_reg ;
  assign \nz.mem [1218] = \nz.mem_1218_sv2v_reg ;
  assign \nz.mem [1217] = \nz.mem_1217_sv2v_reg ;
  assign \nz.mem [1216] = \nz.mem_1216_sv2v_reg ;
  assign \nz.mem [1215] = \nz.mem_1215_sv2v_reg ;
  assign \nz.mem [1214] = \nz.mem_1214_sv2v_reg ;
  assign \nz.mem [1213] = \nz.mem_1213_sv2v_reg ;
  assign \nz.mem [1212] = \nz.mem_1212_sv2v_reg ;
  assign \nz.mem [1211] = \nz.mem_1211_sv2v_reg ;
  assign \nz.mem [1210] = \nz.mem_1210_sv2v_reg ;
  assign \nz.mem [1209] = \nz.mem_1209_sv2v_reg ;
  assign \nz.mem [1208] = \nz.mem_1208_sv2v_reg ;
  assign \nz.mem [1207] = \nz.mem_1207_sv2v_reg ;
  assign \nz.mem [1206] = \nz.mem_1206_sv2v_reg ;
  assign \nz.mem [1205] = \nz.mem_1205_sv2v_reg ;
  assign \nz.mem [1204] = \nz.mem_1204_sv2v_reg ;
  assign \nz.mem [1203] = \nz.mem_1203_sv2v_reg ;
  assign \nz.mem [1202] = \nz.mem_1202_sv2v_reg ;
  assign \nz.mem [1201] = \nz.mem_1201_sv2v_reg ;
  assign \nz.mem [1200] = \nz.mem_1200_sv2v_reg ;
  assign \nz.mem [1199] = \nz.mem_1199_sv2v_reg ;
  assign \nz.mem [1198] = \nz.mem_1198_sv2v_reg ;
  assign \nz.mem [1197] = \nz.mem_1197_sv2v_reg ;
  assign \nz.mem [1196] = \nz.mem_1196_sv2v_reg ;
  assign \nz.mem [1195] = \nz.mem_1195_sv2v_reg ;
  assign \nz.mem [1194] = \nz.mem_1194_sv2v_reg ;
  assign \nz.mem [1193] = \nz.mem_1193_sv2v_reg ;
  assign \nz.mem [1192] = \nz.mem_1192_sv2v_reg ;
  assign \nz.mem [1191] = \nz.mem_1191_sv2v_reg ;
  assign \nz.mem [1190] = \nz.mem_1190_sv2v_reg ;
  assign \nz.mem [1189] = \nz.mem_1189_sv2v_reg ;
  assign \nz.mem [1188] = \nz.mem_1188_sv2v_reg ;
  assign \nz.mem [1187] = \nz.mem_1187_sv2v_reg ;
  assign \nz.mem [1186] = \nz.mem_1186_sv2v_reg ;
  assign \nz.mem [1185] = \nz.mem_1185_sv2v_reg ;
  assign \nz.mem [1184] = \nz.mem_1184_sv2v_reg ;
  assign \nz.mem [1183] = \nz.mem_1183_sv2v_reg ;
  assign \nz.mem [1182] = \nz.mem_1182_sv2v_reg ;
  assign \nz.mem [1181] = \nz.mem_1181_sv2v_reg ;
  assign \nz.mem [1180] = \nz.mem_1180_sv2v_reg ;
  assign \nz.mem [1179] = \nz.mem_1179_sv2v_reg ;
  assign \nz.mem [1178] = \nz.mem_1178_sv2v_reg ;
  assign \nz.mem [1177] = \nz.mem_1177_sv2v_reg ;
  assign \nz.mem [1176] = \nz.mem_1176_sv2v_reg ;
  assign \nz.mem [1175] = \nz.mem_1175_sv2v_reg ;
  assign \nz.mem [1174] = \nz.mem_1174_sv2v_reg ;
  assign \nz.mem [1173] = \nz.mem_1173_sv2v_reg ;
  assign \nz.mem [1172] = \nz.mem_1172_sv2v_reg ;
  assign \nz.mem [1171] = \nz.mem_1171_sv2v_reg ;
  assign \nz.mem [1170] = \nz.mem_1170_sv2v_reg ;
  assign \nz.mem [1169] = \nz.mem_1169_sv2v_reg ;
  assign \nz.mem [1168] = \nz.mem_1168_sv2v_reg ;
  assign \nz.mem [1167] = \nz.mem_1167_sv2v_reg ;
  assign \nz.mem [1166] = \nz.mem_1166_sv2v_reg ;
  assign \nz.mem [1165] = \nz.mem_1165_sv2v_reg ;
  assign \nz.mem [1164] = \nz.mem_1164_sv2v_reg ;
  assign \nz.mem [1163] = \nz.mem_1163_sv2v_reg ;
  assign \nz.mem [1162] = \nz.mem_1162_sv2v_reg ;
  assign \nz.mem [1161] = \nz.mem_1161_sv2v_reg ;
  assign \nz.mem [1160] = \nz.mem_1160_sv2v_reg ;
  assign \nz.mem [1159] = \nz.mem_1159_sv2v_reg ;
  assign \nz.mem [1158] = \nz.mem_1158_sv2v_reg ;
  assign \nz.mem [1157] = \nz.mem_1157_sv2v_reg ;
  assign \nz.mem [1156] = \nz.mem_1156_sv2v_reg ;
  assign \nz.mem [1155] = \nz.mem_1155_sv2v_reg ;
  assign \nz.mem [1154] = \nz.mem_1154_sv2v_reg ;
  assign \nz.mem [1153] = \nz.mem_1153_sv2v_reg ;
  assign \nz.mem [1152] = \nz.mem_1152_sv2v_reg ;
  assign \nz.mem [1151] = \nz.mem_1151_sv2v_reg ;
  assign \nz.mem [1150] = \nz.mem_1150_sv2v_reg ;
  assign \nz.mem [1149] = \nz.mem_1149_sv2v_reg ;
  assign \nz.mem [1148] = \nz.mem_1148_sv2v_reg ;
  assign \nz.mem [1147] = \nz.mem_1147_sv2v_reg ;
  assign \nz.mem [1146] = \nz.mem_1146_sv2v_reg ;
  assign \nz.mem [1145] = \nz.mem_1145_sv2v_reg ;
  assign \nz.mem [1144] = \nz.mem_1144_sv2v_reg ;
  assign \nz.mem [1143] = \nz.mem_1143_sv2v_reg ;
  assign \nz.mem [1142] = \nz.mem_1142_sv2v_reg ;
  assign \nz.mem [1141] = \nz.mem_1141_sv2v_reg ;
  assign \nz.mem [1140] = \nz.mem_1140_sv2v_reg ;
  assign \nz.mem [1139] = \nz.mem_1139_sv2v_reg ;
  assign \nz.mem [1138] = \nz.mem_1138_sv2v_reg ;
  assign \nz.mem [1137] = \nz.mem_1137_sv2v_reg ;
  assign \nz.mem [1136] = \nz.mem_1136_sv2v_reg ;
  assign \nz.mem [1135] = \nz.mem_1135_sv2v_reg ;
  assign \nz.mem [1134] = \nz.mem_1134_sv2v_reg ;
  assign \nz.mem [1133] = \nz.mem_1133_sv2v_reg ;
  assign \nz.mem [1132] = \nz.mem_1132_sv2v_reg ;
  assign \nz.mem [1131] = \nz.mem_1131_sv2v_reg ;
  assign \nz.mem [1130] = \nz.mem_1130_sv2v_reg ;
  assign \nz.mem [1129] = \nz.mem_1129_sv2v_reg ;
  assign \nz.mem [1128] = \nz.mem_1128_sv2v_reg ;
  assign \nz.mem [1127] = \nz.mem_1127_sv2v_reg ;
  assign \nz.mem [1126] = \nz.mem_1126_sv2v_reg ;
  assign \nz.mem [1125] = \nz.mem_1125_sv2v_reg ;
  assign \nz.mem [1124] = \nz.mem_1124_sv2v_reg ;
  assign \nz.mem [1123] = \nz.mem_1123_sv2v_reg ;
  assign \nz.mem [1122] = \nz.mem_1122_sv2v_reg ;
  assign \nz.mem [1121] = \nz.mem_1121_sv2v_reg ;
  assign \nz.mem [1120] = \nz.mem_1120_sv2v_reg ;
  assign \nz.mem [1119] = \nz.mem_1119_sv2v_reg ;
  assign \nz.mem [1118] = \nz.mem_1118_sv2v_reg ;
  assign \nz.mem [1117] = \nz.mem_1117_sv2v_reg ;
  assign \nz.mem [1116] = \nz.mem_1116_sv2v_reg ;
  assign \nz.mem [1115] = \nz.mem_1115_sv2v_reg ;
  assign \nz.mem [1114] = \nz.mem_1114_sv2v_reg ;
  assign \nz.mem [1113] = \nz.mem_1113_sv2v_reg ;
  assign \nz.mem [1112] = \nz.mem_1112_sv2v_reg ;
  assign \nz.mem [1111] = \nz.mem_1111_sv2v_reg ;
  assign \nz.mem [1110] = \nz.mem_1110_sv2v_reg ;
  assign \nz.mem [1109] = \nz.mem_1109_sv2v_reg ;
  assign \nz.mem [1108] = \nz.mem_1108_sv2v_reg ;
  assign \nz.mem [1107] = \nz.mem_1107_sv2v_reg ;
  assign \nz.mem [1106] = \nz.mem_1106_sv2v_reg ;
  assign \nz.mem [1105] = \nz.mem_1105_sv2v_reg ;
  assign \nz.mem [1104] = \nz.mem_1104_sv2v_reg ;
  assign \nz.mem [1103] = \nz.mem_1103_sv2v_reg ;
  assign \nz.mem [1102] = \nz.mem_1102_sv2v_reg ;
  assign \nz.mem [1101] = \nz.mem_1101_sv2v_reg ;
  assign \nz.mem [1100] = \nz.mem_1100_sv2v_reg ;
  assign \nz.mem [1099] = \nz.mem_1099_sv2v_reg ;
  assign \nz.mem [1098] = \nz.mem_1098_sv2v_reg ;
  assign \nz.mem [1097] = \nz.mem_1097_sv2v_reg ;
  assign \nz.mem [1096] = \nz.mem_1096_sv2v_reg ;
  assign \nz.mem [1095] = \nz.mem_1095_sv2v_reg ;
  assign \nz.mem [1094] = \nz.mem_1094_sv2v_reg ;
  assign \nz.mem [1093] = \nz.mem_1093_sv2v_reg ;
  assign \nz.mem [1092] = \nz.mem_1092_sv2v_reg ;
  assign \nz.mem [1091] = \nz.mem_1091_sv2v_reg ;
  assign \nz.mem [1090] = \nz.mem_1090_sv2v_reg ;
  assign \nz.mem [1089] = \nz.mem_1089_sv2v_reg ;
  assign \nz.mem [1088] = \nz.mem_1088_sv2v_reg ;
  assign \nz.mem [1087] = \nz.mem_1087_sv2v_reg ;
  assign \nz.mem [1086] = \nz.mem_1086_sv2v_reg ;
  assign \nz.mem [1085] = \nz.mem_1085_sv2v_reg ;
  assign \nz.mem [1084] = \nz.mem_1084_sv2v_reg ;
  assign \nz.mem [1083] = \nz.mem_1083_sv2v_reg ;
  assign \nz.mem [1082] = \nz.mem_1082_sv2v_reg ;
  assign \nz.mem [1081] = \nz.mem_1081_sv2v_reg ;
  assign \nz.mem [1080] = \nz.mem_1080_sv2v_reg ;
  assign \nz.mem [1079] = \nz.mem_1079_sv2v_reg ;
  assign \nz.mem [1078] = \nz.mem_1078_sv2v_reg ;
  assign \nz.mem [1077] = \nz.mem_1077_sv2v_reg ;
  assign \nz.mem [1076] = \nz.mem_1076_sv2v_reg ;
  assign \nz.mem [1075] = \nz.mem_1075_sv2v_reg ;
  assign \nz.mem [1074] = \nz.mem_1074_sv2v_reg ;
  assign \nz.mem [1073] = \nz.mem_1073_sv2v_reg ;
  assign \nz.mem [1072] = \nz.mem_1072_sv2v_reg ;
  assign \nz.mem [1071] = \nz.mem_1071_sv2v_reg ;
  assign \nz.mem [1070] = \nz.mem_1070_sv2v_reg ;
  assign \nz.mem [1069] = \nz.mem_1069_sv2v_reg ;
  assign \nz.mem [1068] = \nz.mem_1068_sv2v_reg ;
  assign \nz.mem [1067] = \nz.mem_1067_sv2v_reg ;
  assign \nz.mem [1066] = \nz.mem_1066_sv2v_reg ;
  assign \nz.mem [1065] = \nz.mem_1065_sv2v_reg ;
  assign \nz.mem [1064] = \nz.mem_1064_sv2v_reg ;
  assign \nz.mem [1063] = \nz.mem_1063_sv2v_reg ;
  assign \nz.mem [1062] = \nz.mem_1062_sv2v_reg ;
  assign \nz.mem [1061] = \nz.mem_1061_sv2v_reg ;
  assign \nz.mem [1060] = \nz.mem_1060_sv2v_reg ;
  assign \nz.mem [1059] = \nz.mem_1059_sv2v_reg ;
  assign \nz.mem [1058] = \nz.mem_1058_sv2v_reg ;
  assign \nz.mem [1057] = \nz.mem_1057_sv2v_reg ;
  assign \nz.mem [1056] = \nz.mem_1056_sv2v_reg ;
  assign \nz.mem [1055] = \nz.mem_1055_sv2v_reg ;
  assign \nz.mem [1054] = \nz.mem_1054_sv2v_reg ;
  assign \nz.mem [1053] = \nz.mem_1053_sv2v_reg ;
  assign \nz.mem [1052] = \nz.mem_1052_sv2v_reg ;
  assign \nz.mem [1051] = \nz.mem_1051_sv2v_reg ;
  assign \nz.mem [1050] = \nz.mem_1050_sv2v_reg ;
  assign \nz.mem [1049] = \nz.mem_1049_sv2v_reg ;
  assign \nz.mem [1048] = \nz.mem_1048_sv2v_reg ;
  assign \nz.mem [1047] = \nz.mem_1047_sv2v_reg ;
  assign \nz.mem [1046] = \nz.mem_1046_sv2v_reg ;
  assign \nz.mem [1045] = \nz.mem_1045_sv2v_reg ;
  assign \nz.mem [1044] = \nz.mem_1044_sv2v_reg ;
  assign \nz.mem [1043] = \nz.mem_1043_sv2v_reg ;
  assign \nz.mem [1042] = \nz.mem_1042_sv2v_reg ;
  assign \nz.mem [1041] = \nz.mem_1041_sv2v_reg ;
  assign \nz.mem [1040] = \nz.mem_1040_sv2v_reg ;
  assign \nz.mem [1039] = \nz.mem_1039_sv2v_reg ;
  assign \nz.mem [1038] = \nz.mem_1038_sv2v_reg ;
  assign \nz.mem [1037] = \nz.mem_1037_sv2v_reg ;
  assign \nz.mem [1036] = \nz.mem_1036_sv2v_reg ;
  assign \nz.mem [1035] = \nz.mem_1035_sv2v_reg ;
  assign \nz.mem [1034] = \nz.mem_1034_sv2v_reg ;
  assign \nz.mem [1033] = \nz.mem_1033_sv2v_reg ;
  assign \nz.mem [1032] = \nz.mem_1032_sv2v_reg ;
  assign \nz.mem [1031] = \nz.mem_1031_sv2v_reg ;
  assign \nz.mem [1030] = \nz.mem_1030_sv2v_reg ;
  assign \nz.mem [1029] = \nz.mem_1029_sv2v_reg ;
  assign \nz.mem [1028] = \nz.mem_1028_sv2v_reg ;
  assign \nz.mem [1027] = \nz.mem_1027_sv2v_reg ;
  assign \nz.mem [1026] = \nz.mem_1026_sv2v_reg ;
  assign \nz.mem [1025] = \nz.mem_1025_sv2v_reg ;
  assign \nz.mem [1024] = \nz.mem_1024_sv2v_reg ;
  assign \nz.mem [1023] = \nz.mem_1023_sv2v_reg ;
  assign \nz.mem [1022] = \nz.mem_1022_sv2v_reg ;
  assign \nz.mem [1021] = \nz.mem_1021_sv2v_reg ;
  assign \nz.mem [1020] = \nz.mem_1020_sv2v_reg ;
  assign \nz.mem [1019] = \nz.mem_1019_sv2v_reg ;
  assign \nz.mem [1018] = \nz.mem_1018_sv2v_reg ;
  assign \nz.mem [1017] = \nz.mem_1017_sv2v_reg ;
  assign \nz.mem [1016] = \nz.mem_1016_sv2v_reg ;
  assign \nz.mem [1015] = \nz.mem_1015_sv2v_reg ;
  assign \nz.mem [1014] = \nz.mem_1014_sv2v_reg ;
  assign \nz.mem [1013] = \nz.mem_1013_sv2v_reg ;
  assign \nz.mem [1012] = \nz.mem_1012_sv2v_reg ;
  assign \nz.mem [1011] = \nz.mem_1011_sv2v_reg ;
  assign \nz.mem [1010] = \nz.mem_1010_sv2v_reg ;
  assign \nz.mem [1009] = \nz.mem_1009_sv2v_reg ;
  assign \nz.mem [1008] = \nz.mem_1008_sv2v_reg ;
  assign \nz.mem [1007] = \nz.mem_1007_sv2v_reg ;
  assign \nz.mem [1006] = \nz.mem_1006_sv2v_reg ;
  assign \nz.mem [1005] = \nz.mem_1005_sv2v_reg ;
  assign \nz.mem [1004] = \nz.mem_1004_sv2v_reg ;
  assign \nz.mem [1003] = \nz.mem_1003_sv2v_reg ;
  assign \nz.mem [1002] = \nz.mem_1002_sv2v_reg ;
  assign \nz.mem [1001] = \nz.mem_1001_sv2v_reg ;
  assign \nz.mem [1000] = \nz.mem_1000_sv2v_reg ;
  assign \nz.mem [999] = \nz.mem_999_sv2v_reg ;
  assign \nz.mem [998] = \nz.mem_998_sv2v_reg ;
  assign \nz.mem [997] = \nz.mem_997_sv2v_reg ;
  assign \nz.mem [996] = \nz.mem_996_sv2v_reg ;
  assign \nz.mem [995] = \nz.mem_995_sv2v_reg ;
  assign \nz.mem [994] = \nz.mem_994_sv2v_reg ;
  assign \nz.mem [993] = \nz.mem_993_sv2v_reg ;
  assign \nz.mem [992] = \nz.mem_992_sv2v_reg ;
  assign \nz.mem [991] = \nz.mem_991_sv2v_reg ;
  assign \nz.mem [990] = \nz.mem_990_sv2v_reg ;
  assign \nz.mem [989] = \nz.mem_989_sv2v_reg ;
  assign \nz.mem [988] = \nz.mem_988_sv2v_reg ;
  assign \nz.mem [987] = \nz.mem_987_sv2v_reg ;
  assign \nz.mem [986] = \nz.mem_986_sv2v_reg ;
  assign \nz.mem [985] = \nz.mem_985_sv2v_reg ;
  assign \nz.mem [984] = \nz.mem_984_sv2v_reg ;
  assign \nz.mem [983] = \nz.mem_983_sv2v_reg ;
  assign \nz.mem [982] = \nz.mem_982_sv2v_reg ;
  assign \nz.mem [981] = \nz.mem_981_sv2v_reg ;
  assign \nz.mem [980] = \nz.mem_980_sv2v_reg ;
  assign \nz.mem [979] = \nz.mem_979_sv2v_reg ;
  assign \nz.mem [978] = \nz.mem_978_sv2v_reg ;
  assign \nz.mem [977] = \nz.mem_977_sv2v_reg ;
  assign \nz.mem [976] = \nz.mem_976_sv2v_reg ;
  assign \nz.mem [975] = \nz.mem_975_sv2v_reg ;
  assign \nz.mem [974] = \nz.mem_974_sv2v_reg ;
  assign \nz.mem [973] = \nz.mem_973_sv2v_reg ;
  assign \nz.mem [972] = \nz.mem_972_sv2v_reg ;
  assign \nz.mem [971] = \nz.mem_971_sv2v_reg ;
  assign \nz.mem [970] = \nz.mem_970_sv2v_reg ;
  assign \nz.mem [969] = \nz.mem_969_sv2v_reg ;
  assign \nz.mem [968] = \nz.mem_968_sv2v_reg ;
  assign \nz.mem [967] = \nz.mem_967_sv2v_reg ;
  assign \nz.mem [966] = \nz.mem_966_sv2v_reg ;
  assign \nz.mem [965] = \nz.mem_965_sv2v_reg ;
  assign \nz.mem [964] = \nz.mem_964_sv2v_reg ;
  assign \nz.mem [963] = \nz.mem_963_sv2v_reg ;
  assign \nz.mem [962] = \nz.mem_962_sv2v_reg ;
  assign \nz.mem [961] = \nz.mem_961_sv2v_reg ;
  assign \nz.mem [960] = \nz.mem_960_sv2v_reg ;
  assign \nz.mem [959] = \nz.mem_959_sv2v_reg ;
  assign \nz.mem [958] = \nz.mem_958_sv2v_reg ;
  assign \nz.mem [957] = \nz.mem_957_sv2v_reg ;
  assign \nz.mem [956] = \nz.mem_956_sv2v_reg ;
  assign \nz.mem [955] = \nz.mem_955_sv2v_reg ;
  assign \nz.mem [954] = \nz.mem_954_sv2v_reg ;
  assign \nz.mem [953] = \nz.mem_953_sv2v_reg ;
  assign \nz.mem [952] = \nz.mem_952_sv2v_reg ;
  assign \nz.mem [951] = \nz.mem_951_sv2v_reg ;
  assign \nz.mem [950] = \nz.mem_950_sv2v_reg ;
  assign \nz.mem [949] = \nz.mem_949_sv2v_reg ;
  assign \nz.mem [948] = \nz.mem_948_sv2v_reg ;
  assign \nz.mem [947] = \nz.mem_947_sv2v_reg ;
  assign \nz.mem [946] = \nz.mem_946_sv2v_reg ;
  assign \nz.mem [945] = \nz.mem_945_sv2v_reg ;
  assign \nz.mem [944] = \nz.mem_944_sv2v_reg ;
  assign \nz.mem [943] = \nz.mem_943_sv2v_reg ;
  assign \nz.mem [942] = \nz.mem_942_sv2v_reg ;
  assign \nz.mem [941] = \nz.mem_941_sv2v_reg ;
  assign \nz.mem [940] = \nz.mem_940_sv2v_reg ;
  assign \nz.mem [939] = \nz.mem_939_sv2v_reg ;
  assign \nz.mem [938] = \nz.mem_938_sv2v_reg ;
  assign \nz.mem [937] = \nz.mem_937_sv2v_reg ;
  assign \nz.mem [936] = \nz.mem_936_sv2v_reg ;
  assign \nz.mem [935] = \nz.mem_935_sv2v_reg ;
  assign \nz.mem [934] = \nz.mem_934_sv2v_reg ;
  assign \nz.mem [933] = \nz.mem_933_sv2v_reg ;
  assign \nz.mem [932] = \nz.mem_932_sv2v_reg ;
  assign \nz.mem [931] = \nz.mem_931_sv2v_reg ;
  assign \nz.mem [930] = \nz.mem_930_sv2v_reg ;
  assign \nz.mem [929] = \nz.mem_929_sv2v_reg ;
  assign \nz.mem [928] = \nz.mem_928_sv2v_reg ;
  assign \nz.mem [927] = \nz.mem_927_sv2v_reg ;
  assign \nz.mem [926] = \nz.mem_926_sv2v_reg ;
  assign \nz.mem [925] = \nz.mem_925_sv2v_reg ;
  assign \nz.mem [924] = \nz.mem_924_sv2v_reg ;
  assign \nz.mem [923] = \nz.mem_923_sv2v_reg ;
  assign \nz.mem [922] = \nz.mem_922_sv2v_reg ;
  assign \nz.mem [921] = \nz.mem_921_sv2v_reg ;
  assign \nz.mem [920] = \nz.mem_920_sv2v_reg ;
  assign \nz.mem [919] = \nz.mem_919_sv2v_reg ;
  assign \nz.mem [918] = \nz.mem_918_sv2v_reg ;
  assign \nz.mem [917] = \nz.mem_917_sv2v_reg ;
  assign \nz.mem [916] = \nz.mem_916_sv2v_reg ;
  assign \nz.mem [915] = \nz.mem_915_sv2v_reg ;
  assign \nz.mem [914] = \nz.mem_914_sv2v_reg ;
  assign \nz.mem [913] = \nz.mem_913_sv2v_reg ;
  assign \nz.mem [912] = \nz.mem_912_sv2v_reg ;
  assign \nz.mem [911] = \nz.mem_911_sv2v_reg ;
  assign \nz.mem [910] = \nz.mem_910_sv2v_reg ;
  assign \nz.mem [909] = \nz.mem_909_sv2v_reg ;
  assign \nz.mem [908] = \nz.mem_908_sv2v_reg ;
  assign \nz.mem [907] = \nz.mem_907_sv2v_reg ;
  assign \nz.mem [906] = \nz.mem_906_sv2v_reg ;
  assign \nz.mem [905] = \nz.mem_905_sv2v_reg ;
  assign \nz.mem [904] = \nz.mem_904_sv2v_reg ;
  assign \nz.mem [903] = \nz.mem_903_sv2v_reg ;
  assign \nz.mem [902] = \nz.mem_902_sv2v_reg ;
  assign \nz.mem [901] = \nz.mem_901_sv2v_reg ;
  assign \nz.mem [900] = \nz.mem_900_sv2v_reg ;
  assign \nz.mem [899] = \nz.mem_899_sv2v_reg ;
  assign \nz.mem [898] = \nz.mem_898_sv2v_reg ;
  assign \nz.mem [897] = \nz.mem_897_sv2v_reg ;
  assign \nz.mem [896] = \nz.mem_896_sv2v_reg ;
  assign \nz.mem [895] = \nz.mem_895_sv2v_reg ;
  assign \nz.mem [894] = \nz.mem_894_sv2v_reg ;
  assign \nz.mem [893] = \nz.mem_893_sv2v_reg ;
  assign \nz.mem [892] = \nz.mem_892_sv2v_reg ;
  assign \nz.mem [891] = \nz.mem_891_sv2v_reg ;
  assign \nz.mem [890] = \nz.mem_890_sv2v_reg ;
  assign \nz.mem [889] = \nz.mem_889_sv2v_reg ;
  assign \nz.mem [888] = \nz.mem_888_sv2v_reg ;
  assign \nz.mem [887] = \nz.mem_887_sv2v_reg ;
  assign \nz.mem [886] = \nz.mem_886_sv2v_reg ;
  assign \nz.mem [885] = \nz.mem_885_sv2v_reg ;
  assign \nz.mem [884] = \nz.mem_884_sv2v_reg ;
  assign \nz.mem [883] = \nz.mem_883_sv2v_reg ;
  assign \nz.mem [882] = \nz.mem_882_sv2v_reg ;
  assign \nz.mem [881] = \nz.mem_881_sv2v_reg ;
  assign \nz.mem [880] = \nz.mem_880_sv2v_reg ;
  assign \nz.mem [879] = \nz.mem_879_sv2v_reg ;
  assign \nz.mem [878] = \nz.mem_878_sv2v_reg ;
  assign \nz.mem [877] = \nz.mem_877_sv2v_reg ;
  assign \nz.mem [876] = \nz.mem_876_sv2v_reg ;
  assign \nz.mem [875] = \nz.mem_875_sv2v_reg ;
  assign \nz.mem [874] = \nz.mem_874_sv2v_reg ;
  assign \nz.mem [873] = \nz.mem_873_sv2v_reg ;
  assign \nz.mem [872] = \nz.mem_872_sv2v_reg ;
  assign \nz.mem [871] = \nz.mem_871_sv2v_reg ;
  assign \nz.mem [870] = \nz.mem_870_sv2v_reg ;
  assign \nz.mem [869] = \nz.mem_869_sv2v_reg ;
  assign \nz.mem [868] = \nz.mem_868_sv2v_reg ;
  assign \nz.mem [867] = \nz.mem_867_sv2v_reg ;
  assign \nz.mem [866] = \nz.mem_866_sv2v_reg ;
  assign \nz.mem [865] = \nz.mem_865_sv2v_reg ;
  assign \nz.mem [864] = \nz.mem_864_sv2v_reg ;
  assign \nz.mem [863] = \nz.mem_863_sv2v_reg ;
  assign \nz.mem [862] = \nz.mem_862_sv2v_reg ;
  assign \nz.mem [861] = \nz.mem_861_sv2v_reg ;
  assign \nz.mem [860] = \nz.mem_860_sv2v_reg ;
  assign \nz.mem [859] = \nz.mem_859_sv2v_reg ;
  assign \nz.mem [858] = \nz.mem_858_sv2v_reg ;
  assign \nz.mem [857] = \nz.mem_857_sv2v_reg ;
  assign \nz.mem [856] = \nz.mem_856_sv2v_reg ;
  assign \nz.mem [855] = \nz.mem_855_sv2v_reg ;
  assign \nz.mem [854] = \nz.mem_854_sv2v_reg ;
  assign \nz.mem [853] = \nz.mem_853_sv2v_reg ;
  assign \nz.mem [852] = \nz.mem_852_sv2v_reg ;
  assign \nz.mem [851] = \nz.mem_851_sv2v_reg ;
  assign \nz.mem [850] = \nz.mem_850_sv2v_reg ;
  assign \nz.mem [849] = \nz.mem_849_sv2v_reg ;
  assign \nz.mem [848] = \nz.mem_848_sv2v_reg ;
  assign \nz.mem [847] = \nz.mem_847_sv2v_reg ;
  assign \nz.mem [846] = \nz.mem_846_sv2v_reg ;
  assign \nz.mem [845] = \nz.mem_845_sv2v_reg ;
  assign \nz.mem [844] = \nz.mem_844_sv2v_reg ;
  assign \nz.mem [843] = \nz.mem_843_sv2v_reg ;
  assign \nz.mem [842] = \nz.mem_842_sv2v_reg ;
  assign \nz.mem [841] = \nz.mem_841_sv2v_reg ;
  assign \nz.mem [840] = \nz.mem_840_sv2v_reg ;
  assign \nz.mem [839] = \nz.mem_839_sv2v_reg ;
  assign \nz.mem [838] = \nz.mem_838_sv2v_reg ;
  assign \nz.mem [837] = \nz.mem_837_sv2v_reg ;
  assign \nz.mem [836] = \nz.mem_836_sv2v_reg ;
  assign \nz.mem [835] = \nz.mem_835_sv2v_reg ;
  assign \nz.mem [834] = \nz.mem_834_sv2v_reg ;
  assign \nz.mem [833] = \nz.mem_833_sv2v_reg ;
  assign \nz.mem [832] = \nz.mem_832_sv2v_reg ;
  assign \nz.mem [831] = \nz.mem_831_sv2v_reg ;
  assign \nz.mem [830] = \nz.mem_830_sv2v_reg ;
  assign \nz.mem [829] = \nz.mem_829_sv2v_reg ;
  assign \nz.mem [828] = \nz.mem_828_sv2v_reg ;
  assign \nz.mem [827] = \nz.mem_827_sv2v_reg ;
  assign \nz.mem [826] = \nz.mem_826_sv2v_reg ;
  assign \nz.mem [825] = \nz.mem_825_sv2v_reg ;
  assign \nz.mem [824] = \nz.mem_824_sv2v_reg ;
  assign \nz.mem [823] = \nz.mem_823_sv2v_reg ;
  assign \nz.mem [822] = \nz.mem_822_sv2v_reg ;
  assign \nz.mem [821] = \nz.mem_821_sv2v_reg ;
  assign \nz.mem [820] = \nz.mem_820_sv2v_reg ;
  assign \nz.mem [819] = \nz.mem_819_sv2v_reg ;
  assign \nz.mem [818] = \nz.mem_818_sv2v_reg ;
  assign \nz.mem [817] = \nz.mem_817_sv2v_reg ;
  assign \nz.mem [816] = \nz.mem_816_sv2v_reg ;
  assign \nz.mem [815] = \nz.mem_815_sv2v_reg ;
  assign \nz.mem [814] = \nz.mem_814_sv2v_reg ;
  assign \nz.mem [813] = \nz.mem_813_sv2v_reg ;
  assign \nz.mem [812] = \nz.mem_812_sv2v_reg ;
  assign \nz.mem [811] = \nz.mem_811_sv2v_reg ;
  assign \nz.mem [810] = \nz.mem_810_sv2v_reg ;
  assign \nz.mem [809] = \nz.mem_809_sv2v_reg ;
  assign \nz.mem [808] = \nz.mem_808_sv2v_reg ;
  assign \nz.mem [807] = \nz.mem_807_sv2v_reg ;
  assign \nz.mem [806] = \nz.mem_806_sv2v_reg ;
  assign \nz.mem [805] = \nz.mem_805_sv2v_reg ;
  assign \nz.mem [804] = \nz.mem_804_sv2v_reg ;
  assign \nz.mem [803] = \nz.mem_803_sv2v_reg ;
  assign \nz.mem [802] = \nz.mem_802_sv2v_reg ;
  assign \nz.mem [801] = \nz.mem_801_sv2v_reg ;
  assign \nz.mem [800] = \nz.mem_800_sv2v_reg ;
  assign \nz.mem [799] = \nz.mem_799_sv2v_reg ;
  assign \nz.mem [798] = \nz.mem_798_sv2v_reg ;
  assign \nz.mem [797] = \nz.mem_797_sv2v_reg ;
  assign \nz.mem [796] = \nz.mem_796_sv2v_reg ;
  assign \nz.mem [795] = \nz.mem_795_sv2v_reg ;
  assign \nz.mem [794] = \nz.mem_794_sv2v_reg ;
  assign \nz.mem [793] = \nz.mem_793_sv2v_reg ;
  assign \nz.mem [792] = \nz.mem_792_sv2v_reg ;
  assign \nz.mem [791] = \nz.mem_791_sv2v_reg ;
  assign \nz.mem [790] = \nz.mem_790_sv2v_reg ;
  assign \nz.mem [789] = \nz.mem_789_sv2v_reg ;
  assign \nz.mem [788] = \nz.mem_788_sv2v_reg ;
  assign \nz.mem [787] = \nz.mem_787_sv2v_reg ;
  assign \nz.mem [786] = \nz.mem_786_sv2v_reg ;
  assign \nz.mem [785] = \nz.mem_785_sv2v_reg ;
  assign \nz.mem [784] = \nz.mem_784_sv2v_reg ;
  assign \nz.mem [783] = \nz.mem_783_sv2v_reg ;
  assign \nz.mem [782] = \nz.mem_782_sv2v_reg ;
  assign \nz.mem [781] = \nz.mem_781_sv2v_reg ;
  assign \nz.mem [780] = \nz.mem_780_sv2v_reg ;
  assign \nz.mem [779] = \nz.mem_779_sv2v_reg ;
  assign \nz.mem [778] = \nz.mem_778_sv2v_reg ;
  assign \nz.mem [777] = \nz.mem_777_sv2v_reg ;
  assign \nz.mem [776] = \nz.mem_776_sv2v_reg ;
  assign \nz.mem [775] = \nz.mem_775_sv2v_reg ;
  assign \nz.mem [774] = \nz.mem_774_sv2v_reg ;
  assign \nz.mem [773] = \nz.mem_773_sv2v_reg ;
  assign \nz.mem [772] = \nz.mem_772_sv2v_reg ;
  assign \nz.mem [771] = \nz.mem_771_sv2v_reg ;
  assign \nz.mem [770] = \nz.mem_770_sv2v_reg ;
  assign \nz.mem [769] = \nz.mem_769_sv2v_reg ;
  assign \nz.mem [768] = \nz.mem_768_sv2v_reg ;
  assign \nz.mem [767] = \nz.mem_767_sv2v_reg ;
  assign \nz.mem [766] = \nz.mem_766_sv2v_reg ;
  assign \nz.mem [765] = \nz.mem_765_sv2v_reg ;
  assign \nz.mem [764] = \nz.mem_764_sv2v_reg ;
  assign \nz.mem [763] = \nz.mem_763_sv2v_reg ;
  assign \nz.mem [762] = \nz.mem_762_sv2v_reg ;
  assign \nz.mem [761] = \nz.mem_761_sv2v_reg ;
  assign \nz.mem [760] = \nz.mem_760_sv2v_reg ;
  assign \nz.mem [759] = \nz.mem_759_sv2v_reg ;
  assign \nz.mem [758] = \nz.mem_758_sv2v_reg ;
  assign \nz.mem [757] = \nz.mem_757_sv2v_reg ;
  assign \nz.mem [756] = \nz.mem_756_sv2v_reg ;
  assign \nz.mem [755] = \nz.mem_755_sv2v_reg ;
  assign \nz.mem [754] = \nz.mem_754_sv2v_reg ;
  assign \nz.mem [753] = \nz.mem_753_sv2v_reg ;
  assign \nz.mem [752] = \nz.mem_752_sv2v_reg ;
  assign \nz.mem [751] = \nz.mem_751_sv2v_reg ;
  assign \nz.mem [750] = \nz.mem_750_sv2v_reg ;
  assign \nz.mem [749] = \nz.mem_749_sv2v_reg ;
  assign \nz.mem [748] = \nz.mem_748_sv2v_reg ;
  assign \nz.mem [747] = \nz.mem_747_sv2v_reg ;
  assign \nz.mem [746] = \nz.mem_746_sv2v_reg ;
  assign \nz.mem [745] = \nz.mem_745_sv2v_reg ;
  assign \nz.mem [744] = \nz.mem_744_sv2v_reg ;
  assign \nz.mem [743] = \nz.mem_743_sv2v_reg ;
  assign \nz.mem [742] = \nz.mem_742_sv2v_reg ;
  assign \nz.mem [741] = \nz.mem_741_sv2v_reg ;
  assign \nz.mem [740] = \nz.mem_740_sv2v_reg ;
  assign \nz.mem [739] = \nz.mem_739_sv2v_reg ;
  assign \nz.mem [738] = \nz.mem_738_sv2v_reg ;
  assign \nz.mem [737] = \nz.mem_737_sv2v_reg ;
  assign \nz.mem [736] = \nz.mem_736_sv2v_reg ;
  assign \nz.mem [735] = \nz.mem_735_sv2v_reg ;
  assign \nz.mem [734] = \nz.mem_734_sv2v_reg ;
  assign \nz.mem [733] = \nz.mem_733_sv2v_reg ;
  assign \nz.mem [732] = \nz.mem_732_sv2v_reg ;
  assign \nz.mem [731] = \nz.mem_731_sv2v_reg ;
  assign \nz.mem [730] = \nz.mem_730_sv2v_reg ;
  assign \nz.mem [729] = \nz.mem_729_sv2v_reg ;
  assign \nz.mem [728] = \nz.mem_728_sv2v_reg ;
  assign \nz.mem [727] = \nz.mem_727_sv2v_reg ;
  assign \nz.mem [726] = \nz.mem_726_sv2v_reg ;
  assign \nz.mem [725] = \nz.mem_725_sv2v_reg ;
  assign \nz.mem [724] = \nz.mem_724_sv2v_reg ;
  assign \nz.mem [723] = \nz.mem_723_sv2v_reg ;
  assign \nz.mem [722] = \nz.mem_722_sv2v_reg ;
  assign \nz.mem [721] = \nz.mem_721_sv2v_reg ;
  assign \nz.mem [720] = \nz.mem_720_sv2v_reg ;
  assign \nz.mem [719] = \nz.mem_719_sv2v_reg ;
  assign \nz.mem [718] = \nz.mem_718_sv2v_reg ;
  assign \nz.mem [717] = \nz.mem_717_sv2v_reg ;
  assign \nz.mem [716] = \nz.mem_716_sv2v_reg ;
  assign \nz.mem [715] = \nz.mem_715_sv2v_reg ;
  assign \nz.mem [714] = \nz.mem_714_sv2v_reg ;
  assign \nz.mem [713] = \nz.mem_713_sv2v_reg ;
  assign \nz.mem [712] = \nz.mem_712_sv2v_reg ;
  assign \nz.mem [711] = \nz.mem_711_sv2v_reg ;
  assign \nz.mem [710] = \nz.mem_710_sv2v_reg ;
  assign \nz.mem [709] = \nz.mem_709_sv2v_reg ;
  assign \nz.mem [708] = \nz.mem_708_sv2v_reg ;
  assign \nz.mem [707] = \nz.mem_707_sv2v_reg ;
  assign \nz.mem [706] = \nz.mem_706_sv2v_reg ;
  assign \nz.mem [705] = \nz.mem_705_sv2v_reg ;
  assign \nz.mem [704] = \nz.mem_704_sv2v_reg ;
  assign \nz.mem [703] = \nz.mem_703_sv2v_reg ;
  assign \nz.mem [702] = \nz.mem_702_sv2v_reg ;
  assign \nz.mem [701] = \nz.mem_701_sv2v_reg ;
  assign \nz.mem [700] = \nz.mem_700_sv2v_reg ;
  assign \nz.mem [699] = \nz.mem_699_sv2v_reg ;
  assign \nz.mem [698] = \nz.mem_698_sv2v_reg ;
  assign \nz.mem [697] = \nz.mem_697_sv2v_reg ;
  assign \nz.mem [696] = \nz.mem_696_sv2v_reg ;
  assign \nz.mem [695] = \nz.mem_695_sv2v_reg ;
  assign \nz.mem [694] = \nz.mem_694_sv2v_reg ;
  assign \nz.mem [693] = \nz.mem_693_sv2v_reg ;
  assign \nz.mem [692] = \nz.mem_692_sv2v_reg ;
  assign \nz.mem [691] = \nz.mem_691_sv2v_reg ;
  assign \nz.mem [690] = \nz.mem_690_sv2v_reg ;
  assign \nz.mem [689] = \nz.mem_689_sv2v_reg ;
  assign \nz.mem [688] = \nz.mem_688_sv2v_reg ;
  assign \nz.mem [687] = \nz.mem_687_sv2v_reg ;
  assign \nz.mem [686] = \nz.mem_686_sv2v_reg ;
  assign \nz.mem [685] = \nz.mem_685_sv2v_reg ;
  assign \nz.mem [684] = \nz.mem_684_sv2v_reg ;
  assign \nz.mem [683] = \nz.mem_683_sv2v_reg ;
  assign \nz.mem [682] = \nz.mem_682_sv2v_reg ;
  assign \nz.mem [681] = \nz.mem_681_sv2v_reg ;
  assign \nz.mem [680] = \nz.mem_680_sv2v_reg ;
  assign \nz.mem [679] = \nz.mem_679_sv2v_reg ;
  assign \nz.mem [678] = \nz.mem_678_sv2v_reg ;
  assign \nz.mem [677] = \nz.mem_677_sv2v_reg ;
  assign \nz.mem [676] = \nz.mem_676_sv2v_reg ;
  assign \nz.mem [675] = \nz.mem_675_sv2v_reg ;
  assign \nz.mem [674] = \nz.mem_674_sv2v_reg ;
  assign \nz.mem [673] = \nz.mem_673_sv2v_reg ;
  assign \nz.mem [672] = \nz.mem_672_sv2v_reg ;
  assign \nz.mem [671] = \nz.mem_671_sv2v_reg ;
  assign \nz.mem [670] = \nz.mem_670_sv2v_reg ;
  assign \nz.mem [669] = \nz.mem_669_sv2v_reg ;
  assign \nz.mem [668] = \nz.mem_668_sv2v_reg ;
  assign \nz.mem [667] = \nz.mem_667_sv2v_reg ;
  assign \nz.mem [666] = \nz.mem_666_sv2v_reg ;
  assign \nz.mem [665] = \nz.mem_665_sv2v_reg ;
  assign \nz.mem [664] = \nz.mem_664_sv2v_reg ;
  assign \nz.mem [663] = \nz.mem_663_sv2v_reg ;
  assign \nz.mem [662] = \nz.mem_662_sv2v_reg ;
  assign \nz.mem [661] = \nz.mem_661_sv2v_reg ;
  assign \nz.mem [660] = \nz.mem_660_sv2v_reg ;
  assign \nz.mem [659] = \nz.mem_659_sv2v_reg ;
  assign \nz.mem [658] = \nz.mem_658_sv2v_reg ;
  assign \nz.mem [657] = \nz.mem_657_sv2v_reg ;
  assign \nz.mem [656] = \nz.mem_656_sv2v_reg ;
  assign \nz.mem [655] = \nz.mem_655_sv2v_reg ;
  assign \nz.mem [654] = \nz.mem_654_sv2v_reg ;
  assign \nz.mem [653] = \nz.mem_653_sv2v_reg ;
  assign \nz.mem [652] = \nz.mem_652_sv2v_reg ;
  assign \nz.mem [651] = \nz.mem_651_sv2v_reg ;
  assign \nz.mem [650] = \nz.mem_650_sv2v_reg ;
  assign \nz.mem [649] = \nz.mem_649_sv2v_reg ;
  assign \nz.mem [648] = \nz.mem_648_sv2v_reg ;
  assign \nz.mem [647] = \nz.mem_647_sv2v_reg ;
  assign \nz.mem [646] = \nz.mem_646_sv2v_reg ;
  assign \nz.mem [645] = \nz.mem_645_sv2v_reg ;
  assign \nz.mem [644] = \nz.mem_644_sv2v_reg ;
  assign \nz.mem [643] = \nz.mem_643_sv2v_reg ;
  assign \nz.mem [642] = \nz.mem_642_sv2v_reg ;
  assign \nz.mem [641] = \nz.mem_641_sv2v_reg ;
  assign \nz.mem [640] = \nz.mem_640_sv2v_reg ;
  assign \nz.mem [639] = \nz.mem_639_sv2v_reg ;
  assign \nz.mem [638] = \nz.mem_638_sv2v_reg ;
  assign \nz.mem [637] = \nz.mem_637_sv2v_reg ;
  assign \nz.mem [636] = \nz.mem_636_sv2v_reg ;
  assign \nz.mem [635] = \nz.mem_635_sv2v_reg ;
  assign \nz.mem [634] = \nz.mem_634_sv2v_reg ;
  assign \nz.mem [633] = \nz.mem_633_sv2v_reg ;
  assign \nz.mem [632] = \nz.mem_632_sv2v_reg ;
  assign \nz.mem [631] = \nz.mem_631_sv2v_reg ;
  assign \nz.mem [630] = \nz.mem_630_sv2v_reg ;
  assign \nz.mem [629] = \nz.mem_629_sv2v_reg ;
  assign \nz.mem [628] = \nz.mem_628_sv2v_reg ;
  assign \nz.mem [627] = \nz.mem_627_sv2v_reg ;
  assign \nz.mem [626] = \nz.mem_626_sv2v_reg ;
  assign \nz.mem [625] = \nz.mem_625_sv2v_reg ;
  assign \nz.mem [624] = \nz.mem_624_sv2v_reg ;
  assign \nz.mem [623] = \nz.mem_623_sv2v_reg ;
  assign \nz.mem [622] = \nz.mem_622_sv2v_reg ;
  assign \nz.mem [621] = \nz.mem_621_sv2v_reg ;
  assign \nz.mem [620] = \nz.mem_620_sv2v_reg ;
  assign \nz.mem [619] = \nz.mem_619_sv2v_reg ;
  assign \nz.mem [618] = \nz.mem_618_sv2v_reg ;
  assign \nz.mem [617] = \nz.mem_617_sv2v_reg ;
  assign \nz.mem [616] = \nz.mem_616_sv2v_reg ;
  assign \nz.mem [615] = \nz.mem_615_sv2v_reg ;
  assign \nz.mem [614] = \nz.mem_614_sv2v_reg ;
  assign \nz.mem [613] = \nz.mem_613_sv2v_reg ;
  assign \nz.mem [612] = \nz.mem_612_sv2v_reg ;
  assign \nz.mem [611] = \nz.mem_611_sv2v_reg ;
  assign \nz.mem [610] = \nz.mem_610_sv2v_reg ;
  assign \nz.mem [609] = \nz.mem_609_sv2v_reg ;
  assign \nz.mem [608] = \nz.mem_608_sv2v_reg ;
  assign \nz.mem [607] = \nz.mem_607_sv2v_reg ;
  assign \nz.mem [606] = \nz.mem_606_sv2v_reg ;
  assign \nz.mem [605] = \nz.mem_605_sv2v_reg ;
  assign \nz.mem [604] = \nz.mem_604_sv2v_reg ;
  assign \nz.mem [603] = \nz.mem_603_sv2v_reg ;
  assign \nz.mem [602] = \nz.mem_602_sv2v_reg ;
  assign \nz.mem [601] = \nz.mem_601_sv2v_reg ;
  assign \nz.mem [600] = \nz.mem_600_sv2v_reg ;
  assign \nz.mem [599] = \nz.mem_599_sv2v_reg ;
  assign \nz.mem [598] = \nz.mem_598_sv2v_reg ;
  assign \nz.mem [597] = \nz.mem_597_sv2v_reg ;
  assign \nz.mem [596] = \nz.mem_596_sv2v_reg ;
  assign \nz.mem [595] = \nz.mem_595_sv2v_reg ;
  assign \nz.mem [594] = \nz.mem_594_sv2v_reg ;
  assign \nz.mem [593] = \nz.mem_593_sv2v_reg ;
  assign \nz.mem [592] = \nz.mem_592_sv2v_reg ;
  assign \nz.mem [591] = \nz.mem_591_sv2v_reg ;
  assign \nz.mem [590] = \nz.mem_590_sv2v_reg ;
  assign \nz.mem [589] = \nz.mem_589_sv2v_reg ;
  assign \nz.mem [588] = \nz.mem_588_sv2v_reg ;
  assign \nz.mem [587] = \nz.mem_587_sv2v_reg ;
  assign \nz.mem [586] = \nz.mem_586_sv2v_reg ;
  assign \nz.mem [585] = \nz.mem_585_sv2v_reg ;
  assign \nz.mem [584] = \nz.mem_584_sv2v_reg ;
  assign \nz.mem [583] = \nz.mem_583_sv2v_reg ;
  assign \nz.mem [582] = \nz.mem_582_sv2v_reg ;
  assign \nz.mem [581] = \nz.mem_581_sv2v_reg ;
  assign \nz.mem [580] = \nz.mem_580_sv2v_reg ;
  assign \nz.mem [579] = \nz.mem_579_sv2v_reg ;
  assign \nz.mem [578] = \nz.mem_578_sv2v_reg ;
  assign \nz.mem [577] = \nz.mem_577_sv2v_reg ;
  assign \nz.mem [576] = \nz.mem_576_sv2v_reg ;
  assign \nz.mem [575] = \nz.mem_575_sv2v_reg ;
  assign \nz.mem [574] = \nz.mem_574_sv2v_reg ;
  assign \nz.mem [573] = \nz.mem_573_sv2v_reg ;
  assign \nz.mem [572] = \nz.mem_572_sv2v_reg ;
  assign \nz.mem [571] = \nz.mem_571_sv2v_reg ;
  assign \nz.mem [570] = \nz.mem_570_sv2v_reg ;
  assign \nz.mem [569] = \nz.mem_569_sv2v_reg ;
  assign \nz.mem [568] = \nz.mem_568_sv2v_reg ;
  assign \nz.mem [567] = \nz.mem_567_sv2v_reg ;
  assign \nz.mem [566] = \nz.mem_566_sv2v_reg ;
  assign \nz.mem [565] = \nz.mem_565_sv2v_reg ;
  assign \nz.mem [564] = \nz.mem_564_sv2v_reg ;
  assign \nz.mem [563] = \nz.mem_563_sv2v_reg ;
  assign \nz.mem [562] = \nz.mem_562_sv2v_reg ;
  assign \nz.mem [561] = \nz.mem_561_sv2v_reg ;
  assign \nz.mem [560] = \nz.mem_560_sv2v_reg ;
  assign \nz.mem [559] = \nz.mem_559_sv2v_reg ;
  assign \nz.mem [558] = \nz.mem_558_sv2v_reg ;
  assign \nz.mem [557] = \nz.mem_557_sv2v_reg ;
  assign \nz.mem [556] = \nz.mem_556_sv2v_reg ;
  assign \nz.mem [555] = \nz.mem_555_sv2v_reg ;
  assign \nz.mem [554] = \nz.mem_554_sv2v_reg ;
  assign \nz.mem [553] = \nz.mem_553_sv2v_reg ;
  assign \nz.mem [552] = \nz.mem_552_sv2v_reg ;
  assign \nz.mem [551] = \nz.mem_551_sv2v_reg ;
  assign \nz.mem [550] = \nz.mem_550_sv2v_reg ;
  assign \nz.mem [549] = \nz.mem_549_sv2v_reg ;
  assign \nz.mem [548] = \nz.mem_548_sv2v_reg ;
  assign \nz.mem [547] = \nz.mem_547_sv2v_reg ;
  assign \nz.mem [546] = \nz.mem_546_sv2v_reg ;
  assign \nz.mem [545] = \nz.mem_545_sv2v_reg ;
  assign \nz.mem [544] = \nz.mem_544_sv2v_reg ;
  assign \nz.mem [543] = \nz.mem_543_sv2v_reg ;
  assign \nz.mem [542] = \nz.mem_542_sv2v_reg ;
  assign \nz.mem [541] = \nz.mem_541_sv2v_reg ;
  assign \nz.mem [540] = \nz.mem_540_sv2v_reg ;
  assign \nz.mem [539] = \nz.mem_539_sv2v_reg ;
  assign \nz.mem [538] = \nz.mem_538_sv2v_reg ;
  assign \nz.mem [537] = \nz.mem_537_sv2v_reg ;
  assign \nz.mem [536] = \nz.mem_536_sv2v_reg ;
  assign \nz.mem [535] = \nz.mem_535_sv2v_reg ;
  assign \nz.mem [534] = \nz.mem_534_sv2v_reg ;
  assign \nz.mem [533] = \nz.mem_533_sv2v_reg ;
  assign \nz.mem [532] = \nz.mem_532_sv2v_reg ;
  assign \nz.mem [531] = \nz.mem_531_sv2v_reg ;
  assign \nz.mem [530] = \nz.mem_530_sv2v_reg ;
  assign \nz.mem [529] = \nz.mem_529_sv2v_reg ;
  assign \nz.mem [528] = \nz.mem_528_sv2v_reg ;
  assign \nz.mem [527] = \nz.mem_527_sv2v_reg ;
  assign \nz.mem [526] = \nz.mem_526_sv2v_reg ;
  assign \nz.mem [525] = \nz.mem_525_sv2v_reg ;
  assign \nz.mem [524] = \nz.mem_524_sv2v_reg ;
  assign \nz.mem [523] = \nz.mem_523_sv2v_reg ;
  assign \nz.mem [522] = \nz.mem_522_sv2v_reg ;
  assign \nz.mem [521] = \nz.mem_521_sv2v_reg ;
  assign \nz.mem [520] = \nz.mem_520_sv2v_reg ;
  assign \nz.mem [519] = \nz.mem_519_sv2v_reg ;
  assign \nz.mem [518] = \nz.mem_518_sv2v_reg ;
  assign \nz.mem [517] = \nz.mem_517_sv2v_reg ;
  assign \nz.mem [516] = \nz.mem_516_sv2v_reg ;
  assign \nz.mem [515] = \nz.mem_515_sv2v_reg ;
  assign \nz.mem [514] = \nz.mem_514_sv2v_reg ;
  assign \nz.mem [513] = \nz.mem_513_sv2v_reg ;
  assign \nz.mem [512] = \nz.mem_512_sv2v_reg ;
  assign \nz.mem [511] = \nz.mem_511_sv2v_reg ;
  assign \nz.mem [510] = \nz.mem_510_sv2v_reg ;
  assign \nz.mem [509] = \nz.mem_509_sv2v_reg ;
  assign \nz.mem [508] = \nz.mem_508_sv2v_reg ;
  assign \nz.mem [507] = \nz.mem_507_sv2v_reg ;
  assign \nz.mem [506] = \nz.mem_506_sv2v_reg ;
  assign \nz.mem [505] = \nz.mem_505_sv2v_reg ;
  assign \nz.mem [504] = \nz.mem_504_sv2v_reg ;
  assign \nz.mem [503] = \nz.mem_503_sv2v_reg ;
  assign \nz.mem [502] = \nz.mem_502_sv2v_reg ;
  assign \nz.mem [501] = \nz.mem_501_sv2v_reg ;
  assign \nz.mem [500] = \nz.mem_500_sv2v_reg ;
  assign \nz.mem [499] = \nz.mem_499_sv2v_reg ;
  assign \nz.mem [498] = \nz.mem_498_sv2v_reg ;
  assign \nz.mem [497] = \nz.mem_497_sv2v_reg ;
  assign \nz.mem [496] = \nz.mem_496_sv2v_reg ;
  assign \nz.mem [495] = \nz.mem_495_sv2v_reg ;
  assign \nz.mem [494] = \nz.mem_494_sv2v_reg ;
  assign \nz.mem [493] = \nz.mem_493_sv2v_reg ;
  assign \nz.mem [492] = \nz.mem_492_sv2v_reg ;
  assign \nz.mem [491] = \nz.mem_491_sv2v_reg ;
  assign \nz.mem [490] = \nz.mem_490_sv2v_reg ;
  assign \nz.mem [489] = \nz.mem_489_sv2v_reg ;
  assign \nz.mem [488] = \nz.mem_488_sv2v_reg ;
  assign \nz.mem [487] = \nz.mem_487_sv2v_reg ;
  assign \nz.mem [486] = \nz.mem_486_sv2v_reg ;
  assign \nz.mem [485] = \nz.mem_485_sv2v_reg ;
  assign \nz.mem [484] = \nz.mem_484_sv2v_reg ;
  assign \nz.mem [483] = \nz.mem_483_sv2v_reg ;
  assign \nz.mem [482] = \nz.mem_482_sv2v_reg ;
  assign \nz.mem [481] = \nz.mem_481_sv2v_reg ;
  assign \nz.mem [480] = \nz.mem_480_sv2v_reg ;
  assign \nz.mem [479] = \nz.mem_479_sv2v_reg ;
  assign \nz.mem [478] = \nz.mem_478_sv2v_reg ;
  assign \nz.mem [477] = \nz.mem_477_sv2v_reg ;
  assign \nz.mem [476] = \nz.mem_476_sv2v_reg ;
  assign \nz.mem [475] = \nz.mem_475_sv2v_reg ;
  assign \nz.mem [474] = \nz.mem_474_sv2v_reg ;
  assign \nz.mem [473] = \nz.mem_473_sv2v_reg ;
  assign \nz.mem [472] = \nz.mem_472_sv2v_reg ;
  assign \nz.mem [471] = \nz.mem_471_sv2v_reg ;
  assign \nz.mem [470] = \nz.mem_470_sv2v_reg ;
  assign \nz.mem [469] = \nz.mem_469_sv2v_reg ;
  assign \nz.mem [468] = \nz.mem_468_sv2v_reg ;
  assign \nz.mem [467] = \nz.mem_467_sv2v_reg ;
  assign \nz.mem [466] = \nz.mem_466_sv2v_reg ;
  assign \nz.mem [465] = \nz.mem_465_sv2v_reg ;
  assign \nz.mem [464] = \nz.mem_464_sv2v_reg ;
  assign \nz.mem [463] = \nz.mem_463_sv2v_reg ;
  assign \nz.mem [462] = \nz.mem_462_sv2v_reg ;
  assign \nz.mem [461] = \nz.mem_461_sv2v_reg ;
  assign \nz.mem [460] = \nz.mem_460_sv2v_reg ;
  assign \nz.mem [459] = \nz.mem_459_sv2v_reg ;
  assign \nz.mem [458] = \nz.mem_458_sv2v_reg ;
  assign \nz.mem [457] = \nz.mem_457_sv2v_reg ;
  assign \nz.mem [456] = \nz.mem_456_sv2v_reg ;
  assign \nz.mem [455] = \nz.mem_455_sv2v_reg ;
  assign \nz.mem [454] = \nz.mem_454_sv2v_reg ;
  assign \nz.mem [453] = \nz.mem_453_sv2v_reg ;
  assign \nz.mem [452] = \nz.mem_452_sv2v_reg ;
  assign \nz.mem [451] = \nz.mem_451_sv2v_reg ;
  assign \nz.mem [450] = \nz.mem_450_sv2v_reg ;
  assign \nz.mem [449] = \nz.mem_449_sv2v_reg ;
  assign \nz.mem [448] = \nz.mem_448_sv2v_reg ;
  assign \nz.mem [447] = \nz.mem_447_sv2v_reg ;
  assign \nz.mem [446] = \nz.mem_446_sv2v_reg ;
  assign \nz.mem [445] = \nz.mem_445_sv2v_reg ;
  assign \nz.mem [444] = \nz.mem_444_sv2v_reg ;
  assign \nz.mem [443] = \nz.mem_443_sv2v_reg ;
  assign \nz.mem [442] = \nz.mem_442_sv2v_reg ;
  assign \nz.mem [441] = \nz.mem_441_sv2v_reg ;
  assign \nz.mem [440] = \nz.mem_440_sv2v_reg ;
  assign \nz.mem [439] = \nz.mem_439_sv2v_reg ;
  assign \nz.mem [438] = \nz.mem_438_sv2v_reg ;
  assign \nz.mem [437] = \nz.mem_437_sv2v_reg ;
  assign \nz.mem [436] = \nz.mem_436_sv2v_reg ;
  assign \nz.mem [435] = \nz.mem_435_sv2v_reg ;
  assign \nz.mem [434] = \nz.mem_434_sv2v_reg ;
  assign \nz.mem [433] = \nz.mem_433_sv2v_reg ;
  assign \nz.mem [432] = \nz.mem_432_sv2v_reg ;
  assign \nz.mem [431] = \nz.mem_431_sv2v_reg ;
  assign \nz.mem [430] = \nz.mem_430_sv2v_reg ;
  assign \nz.mem [429] = \nz.mem_429_sv2v_reg ;
  assign \nz.mem [428] = \nz.mem_428_sv2v_reg ;
  assign \nz.mem [427] = \nz.mem_427_sv2v_reg ;
  assign \nz.mem [426] = \nz.mem_426_sv2v_reg ;
  assign \nz.mem [425] = \nz.mem_425_sv2v_reg ;
  assign \nz.mem [424] = \nz.mem_424_sv2v_reg ;
  assign \nz.mem [423] = \nz.mem_423_sv2v_reg ;
  assign \nz.mem [422] = \nz.mem_422_sv2v_reg ;
  assign \nz.mem [421] = \nz.mem_421_sv2v_reg ;
  assign \nz.mem [420] = \nz.mem_420_sv2v_reg ;
  assign \nz.mem [419] = \nz.mem_419_sv2v_reg ;
  assign \nz.mem [418] = \nz.mem_418_sv2v_reg ;
  assign \nz.mem [417] = \nz.mem_417_sv2v_reg ;
  assign \nz.mem [416] = \nz.mem_416_sv2v_reg ;
  assign \nz.mem [415] = \nz.mem_415_sv2v_reg ;
  assign \nz.mem [414] = \nz.mem_414_sv2v_reg ;
  assign \nz.mem [413] = \nz.mem_413_sv2v_reg ;
  assign \nz.mem [412] = \nz.mem_412_sv2v_reg ;
  assign \nz.mem [411] = \nz.mem_411_sv2v_reg ;
  assign \nz.mem [410] = \nz.mem_410_sv2v_reg ;
  assign \nz.mem [409] = \nz.mem_409_sv2v_reg ;
  assign \nz.mem [408] = \nz.mem_408_sv2v_reg ;
  assign \nz.mem [407] = \nz.mem_407_sv2v_reg ;
  assign \nz.mem [406] = \nz.mem_406_sv2v_reg ;
  assign \nz.mem [405] = \nz.mem_405_sv2v_reg ;
  assign \nz.mem [404] = \nz.mem_404_sv2v_reg ;
  assign \nz.mem [403] = \nz.mem_403_sv2v_reg ;
  assign \nz.mem [402] = \nz.mem_402_sv2v_reg ;
  assign \nz.mem [401] = \nz.mem_401_sv2v_reg ;
  assign \nz.mem [400] = \nz.mem_400_sv2v_reg ;
  assign \nz.mem [399] = \nz.mem_399_sv2v_reg ;
  assign \nz.mem [398] = \nz.mem_398_sv2v_reg ;
  assign \nz.mem [397] = \nz.mem_397_sv2v_reg ;
  assign \nz.mem [396] = \nz.mem_396_sv2v_reg ;
  assign \nz.mem [395] = \nz.mem_395_sv2v_reg ;
  assign \nz.mem [394] = \nz.mem_394_sv2v_reg ;
  assign \nz.mem [393] = \nz.mem_393_sv2v_reg ;
  assign \nz.mem [392] = \nz.mem_392_sv2v_reg ;
  assign \nz.mem [391] = \nz.mem_391_sv2v_reg ;
  assign \nz.mem [390] = \nz.mem_390_sv2v_reg ;
  assign \nz.mem [389] = \nz.mem_389_sv2v_reg ;
  assign \nz.mem [388] = \nz.mem_388_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[173] = (N17)? \nz.mem [173] : 
                         (N19)? \nz.mem [347] : 
                         (N21)? \nz.mem [521] : 
                         (N23)? \nz.mem [695] : 
                         (N18)? \nz.mem [869] : 
                         (N20)? \nz.mem [1043] : 
                         (N22)? \nz.mem [1217] : 
                         (N24)? \nz.mem [1391] : 1'b0;
  assign r_data_o[172] = (N17)? \nz.mem [172] : 
                         (N19)? \nz.mem [346] : 
                         (N21)? \nz.mem [520] : 
                         (N23)? \nz.mem [694] : 
                         (N18)? \nz.mem [868] : 
                         (N20)? \nz.mem [1042] : 
                         (N22)? \nz.mem [1216] : 
                         (N24)? \nz.mem [1390] : 1'b0;
  assign r_data_o[171] = (N17)? \nz.mem [171] : 
                         (N19)? \nz.mem [345] : 
                         (N21)? \nz.mem [519] : 
                         (N23)? \nz.mem [693] : 
                         (N18)? \nz.mem [867] : 
                         (N20)? \nz.mem [1041] : 
                         (N22)? \nz.mem [1215] : 
                         (N24)? \nz.mem [1389] : 1'b0;
  assign r_data_o[170] = (N17)? \nz.mem [170] : 
                         (N19)? \nz.mem [344] : 
                         (N21)? \nz.mem [518] : 
                         (N23)? \nz.mem [692] : 
                         (N18)? \nz.mem [866] : 
                         (N20)? \nz.mem [1040] : 
                         (N22)? \nz.mem [1214] : 
                         (N24)? \nz.mem [1388] : 1'b0;
  assign r_data_o[169] = (N17)? \nz.mem [169] : 
                         (N19)? \nz.mem [343] : 
                         (N21)? \nz.mem [517] : 
                         (N23)? \nz.mem [691] : 
                         (N18)? \nz.mem [865] : 
                         (N20)? \nz.mem [1039] : 
                         (N22)? \nz.mem [1213] : 
                         (N24)? \nz.mem [1387] : 1'b0;
  assign r_data_o[168] = (N17)? \nz.mem [168] : 
                         (N19)? \nz.mem [342] : 
                         (N21)? \nz.mem [516] : 
                         (N23)? \nz.mem [690] : 
                         (N18)? \nz.mem [864] : 
                         (N20)? \nz.mem [1038] : 
                         (N22)? \nz.mem [1212] : 
                         (N24)? \nz.mem [1386] : 1'b0;
  assign r_data_o[167] = (N17)? \nz.mem [167] : 
                         (N19)? \nz.mem [341] : 
                         (N21)? \nz.mem [515] : 
                         (N23)? \nz.mem [689] : 
                         (N18)? \nz.mem [863] : 
                         (N20)? \nz.mem [1037] : 
                         (N22)? \nz.mem [1211] : 
                         (N24)? \nz.mem [1385] : 1'b0;
  assign r_data_o[166] = (N17)? \nz.mem [166] : 
                         (N19)? \nz.mem [340] : 
                         (N21)? \nz.mem [514] : 
                         (N23)? \nz.mem [688] : 
                         (N18)? \nz.mem [862] : 
                         (N20)? \nz.mem [1036] : 
                         (N22)? \nz.mem [1210] : 
                         (N24)? \nz.mem [1384] : 1'b0;
  assign r_data_o[165] = (N17)? \nz.mem [165] : 
                         (N19)? \nz.mem [339] : 
                         (N21)? \nz.mem [513] : 
                         (N23)? \nz.mem [687] : 
                         (N18)? \nz.mem [861] : 
                         (N20)? \nz.mem [1035] : 
                         (N22)? \nz.mem [1209] : 
                         (N24)? \nz.mem [1383] : 1'b0;
  assign r_data_o[164] = (N17)? \nz.mem [164] : 
                         (N19)? \nz.mem [338] : 
                         (N21)? \nz.mem [512] : 
                         (N23)? \nz.mem [686] : 
                         (N18)? \nz.mem [860] : 
                         (N20)? \nz.mem [1034] : 
                         (N22)? \nz.mem [1208] : 
                         (N24)? \nz.mem [1382] : 1'b0;
  assign r_data_o[163] = (N17)? \nz.mem [163] : 
                         (N19)? \nz.mem [337] : 
                         (N21)? \nz.mem [511] : 
                         (N23)? \nz.mem [685] : 
                         (N18)? \nz.mem [859] : 
                         (N20)? \nz.mem [1033] : 
                         (N22)? \nz.mem [1207] : 
                         (N24)? \nz.mem [1381] : 1'b0;
  assign r_data_o[162] = (N17)? \nz.mem [162] : 
                         (N19)? \nz.mem [336] : 
                         (N21)? \nz.mem [510] : 
                         (N23)? \nz.mem [684] : 
                         (N18)? \nz.mem [858] : 
                         (N20)? \nz.mem [1032] : 
                         (N22)? \nz.mem [1206] : 
                         (N24)? \nz.mem [1380] : 1'b0;
  assign r_data_o[161] = (N17)? \nz.mem [161] : 
                         (N19)? \nz.mem [335] : 
                         (N21)? \nz.mem [509] : 
                         (N23)? \nz.mem [683] : 
                         (N18)? \nz.mem [857] : 
                         (N20)? \nz.mem [1031] : 
                         (N22)? \nz.mem [1205] : 
                         (N24)? \nz.mem [1379] : 1'b0;
  assign r_data_o[160] = (N17)? \nz.mem [160] : 
                         (N19)? \nz.mem [334] : 
                         (N21)? \nz.mem [508] : 
                         (N23)? \nz.mem [682] : 
                         (N18)? \nz.mem [856] : 
                         (N20)? \nz.mem [1030] : 
                         (N22)? \nz.mem [1204] : 
                         (N24)? \nz.mem [1378] : 1'b0;
  assign r_data_o[159] = (N17)? \nz.mem [159] : 
                         (N19)? \nz.mem [333] : 
                         (N21)? \nz.mem [507] : 
                         (N23)? \nz.mem [681] : 
                         (N18)? \nz.mem [855] : 
                         (N20)? \nz.mem [1029] : 
                         (N22)? \nz.mem [1203] : 
                         (N24)? \nz.mem [1377] : 1'b0;
  assign r_data_o[158] = (N17)? \nz.mem [158] : 
                         (N19)? \nz.mem [332] : 
                         (N21)? \nz.mem [506] : 
                         (N23)? \nz.mem [680] : 
                         (N18)? \nz.mem [854] : 
                         (N20)? \nz.mem [1028] : 
                         (N22)? \nz.mem [1202] : 
                         (N24)? \nz.mem [1376] : 1'b0;
  assign r_data_o[157] = (N17)? \nz.mem [157] : 
                         (N19)? \nz.mem [331] : 
                         (N21)? \nz.mem [505] : 
                         (N23)? \nz.mem [679] : 
                         (N18)? \nz.mem [853] : 
                         (N20)? \nz.mem [1027] : 
                         (N22)? \nz.mem [1201] : 
                         (N24)? \nz.mem [1375] : 1'b0;
  assign r_data_o[156] = (N17)? \nz.mem [156] : 
                         (N19)? \nz.mem [330] : 
                         (N21)? \nz.mem [504] : 
                         (N23)? \nz.mem [678] : 
                         (N18)? \nz.mem [852] : 
                         (N20)? \nz.mem [1026] : 
                         (N22)? \nz.mem [1200] : 
                         (N24)? \nz.mem [1374] : 1'b0;
  assign r_data_o[155] = (N17)? \nz.mem [155] : 
                         (N19)? \nz.mem [329] : 
                         (N21)? \nz.mem [503] : 
                         (N23)? \nz.mem [677] : 
                         (N18)? \nz.mem [851] : 
                         (N20)? \nz.mem [1025] : 
                         (N22)? \nz.mem [1199] : 
                         (N24)? \nz.mem [1373] : 1'b0;
  assign r_data_o[154] = (N17)? \nz.mem [154] : 
                         (N19)? \nz.mem [328] : 
                         (N21)? \nz.mem [502] : 
                         (N23)? \nz.mem [676] : 
                         (N18)? \nz.mem [850] : 
                         (N20)? \nz.mem [1024] : 
                         (N22)? \nz.mem [1198] : 
                         (N24)? \nz.mem [1372] : 1'b0;
  assign r_data_o[153] = (N17)? \nz.mem [153] : 
                         (N19)? \nz.mem [327] : 
                         (N21)? \nz.mem [501] : 
                         (N23)? \nz.mem [675] : 
                         (N18)? \nz.mem [849] : 
                         (N20)? \nz.mem [1023] : 
                         (N22)? \nz.mem [1197] : 
                         (N24)? \nz.mem [1371] : 1'b0;
  assign r_data_o[152] = (N17)? \nz.mem [152] : 
                         (N19)? \nz.mem [326] : 
                         (N21)? \nz.mem [500] : 
                         (N23)? \nz.mem [674] : 
                         (N18)? \nz.mem [848] : 
                         (N20)? \nz.mem [1022] : 
                         (N22)? \nz.mem [1196] : 
                         (N24)? \nz.mem [1370] : 1'b0;
  assign r_data_o[151] = (N17)? \nz.mem [151] : 
                         (N19)? \nz.mem [325] : 
                         (N21)? \nz.mem [499] : 
                         (N23)? \nz.mem [673] : 
                         (N18)? \nz.mem [847] : 
                         (N20)? \nz.mem [1021] : 
                         (N22)? \nz.mem [1195] : 
                         (N24)? \nz.mem [1369] : 1'b0;
  assign r_data_o[150] = (N17)? \nz.mem [150] : 
                         (N19)? \nz.mem [324] : 
                         (N21)? \nz.mem [498] : 
                         (N23)? \nz.mem [672] : 
                         (N18)? \nz.mem [846] : 
                         (N20)? \nz.mem [1020] : 
                         (N22)? \nz.mem [1194] : 
                         (N24)? \nz.mem [1368] : 1'b0;
  assign r_data_o[149] = (N17)? \nz.mem [149] : 
                         (N19)? \nz.mem [323] : 
                         (N21)? \nz.mem [497] : 
                         (N23)? \nz.mem [671] : 
                         (N18)? \nz.mem [845] : 
                         (N20)? \nz.mem [1019] : 
                         (N22)? \nz.mem [1193] : 
                         (N24)? \nz.mem [1367] : 1'b0;
  assign r_data_o[148] = (N17)? \nz.mem [148] : 
                         (N19)? \nz.mem [322] : 
                         (N21)? \nz.mem [496] : 
                         (N23)? \nz.mem [670] : 
                         (N18)? \nz.mem [844] : 
                         (N20)? \nz.mem [1018] : 
                         (N22)? \nz.mem [1192] : 
                         (N24)? \nz.mem [1366] : 1'b0;
  assign r_data_o[147] = (N17)? \nz.mem [147] : 
                         (N19)? \nz.mem [321] : 
                         (N21)? \nz.mem [495] : 
                         (N23)? \nz.mem [669] : 
                         (N18)? \nz.mem [843] : 
                         (N20)? \nz.mem [1017] : 
                         (N22)? \nz.mem [1191] : 
                         (N24)? \nz.mem [1365] : 1'b0;
  assign r_data_o[146] = (N17)? \nz.mem [146] : 
                         (N19)? \nz.mem [320] : 
                         (N21)? \nz.mem [494] : 
                         (N23)? \nz.mem [668] : 
                         (N18)? \nz.mem [842] : 
                         (N20)? \nz.mem [1016] : 
                         (N22)? \nz.mem [1190] : 
                         (N24)? \nz.mem [1364] : 1'b0;
  assign r_data_o[145] = (N17)? \nz.mem [145] : 
                         (N19)? \nz.mem [319] : 
                         (N21)? \nz.mem [493] : 
                         (N23)? \nz.mem [667] : 
                         (N18)? \nz.mem [841] : 
                         (N20)? \nz.mem [1015] : 
                         (N22)? \nz.mem [1189] : 
                         (N24)? \nz.mem [1363] : 1'b0;
  assign r_data_o[144] = (N17)? \nz.mem [144] : 
                         (N19)? \nz.mem [318] : 
                         (N21)? \nz.mem [492] : 
                         (N23)? \nz.mem [666] : 
                         (N18)? \nz.mem [840] : 
                         (N20)? \nz.mem [1014] : 
                         (N22)? \nz.mem [1188] : 
                         (N24)? \nz.mem [1362] : 1'b0;
  assign r_data_o[143] = (N17)? \nz.mem [143] : 
                         (N19)? \nz.mem [317] : 
                         (N21)? \nz.mem [491] : 
                         (N23)? \nz.mem [665] : 
                         (N18)? \nz.mem [839] : 
                         (N20)? \nz.mem [1013] : 
                         (N22)? \nz.mem [1187] : 
                         (N24)? \nz.mem [1361] : 1'b0;
  assign r_data_o[142] = (N17)? \nz.mem [142] : 
                         (N19)? \nz.mem [316] : 
                         (N21)? \nz.mem [490] : 
                         (N23)? \nz.mem [664] : 
                         (N18)? \nz.mem [838] : 
                         (N20)? \nz.mem [1012] : 
                         (N22)? \nz.mem [1186] : 
                         (N24)? \nz.mem [1360] : 1'b0;
  assign r_data_o[141] = (N17)? \nz.mem [141] : 
                         (N19)? \nz.mem [315] : 
                         (N21)? \nz.mem [489] : 
                         (N23)? \nz.mem [663] : 
                         (N18)? \nz.mem [837] : 
                         (N20)? \nz.mem [1011] : 
                         (N22)? \nz.mem [1185] : 
                         (N24)? \nz.mem [1359] : 1'b0;
  assign r_data_o[140] = (N17)? \nz.mem [140] : 
                         (N19)? \nz.mem [314] : 
                         (N21)? \nz.mem [488] : 
                         (N23)? \nz.mem [662] : 
                         (N18)? \nz.mem [836] : 
                         (N20)? \nz.mem [1010] : 
                         (N22)? \nz.mem [1184] : 
                         (N24)? \nz.mem [1358] : 1'b0;
  assign r_data_o[139] = (N17)? \nz.mem [139] : 
                         (N19)? \nz.mem [313] : 
                         (N21)? \nz.mem [487] : 
                         (N23)? \nz.mem [661] : 
                         (N18)? \nz.mem [835] : 
                         (N20)? \nz.mem [1009] : 
                         (N22)? \nz.mem [1183] : 
                         (N24)? \nz.mem [1357] : 1'b0;
  assign r_data_o[138] = (N17)? \nz.mem [138] : 
                         (N19)? \nz.mem [312] : 
                         (N21)? \nz.mem [486] : 
                         (N23)? \nz.mem [660] : 
                         (N18)? \nz.mem [834] : 
                         (N20)? \nz.mem [1008] : 
                         (N22)? \nz.mem [1182] : 
                         (N24)? \nz.mem [1356] : 1'b0;
  assign r_data_o[137] = (N17)? \nz.mem [137] : 
                         (N19)? \nz.mem [311] : 
                         (N21)? \nz.mem [485] : 
                         (N23)? \nz.mem [659] : 
                         (N18)? \nz.mem [833] : 
                         (N20)? \nz.mem [1007] : 
                         (N22)? \nz.mem [1181] : 
                         (N24)? \nz.mem [1355] : 1'b0;
  assign r_data_o[136] = (N17)? \nz.mem [136] : 
                         (N19)? \nz.mem [310] : 
                         (N21)? \nz.mem [484] : 
                         (N23)? \nz.mem [658] : 
                         (N18)? \nz.mem [832] : 
                         (N20)? \nz.mem [1006] : 
                         (N22)? \nz.mem [1180] : 
                         (N24)? \nz.mem [1354] : 1'b0;
  assign r_data_o[135] = (N17)? \nz.mem [135] : 
                         (N19)? \nz.mem [309] : 
                         (N21)? \nz.mem [483] : 
                         (N23)? \nz.mem [657] : 
                         (N18)? \nz.mem [831] : 
                         (N20)? \nz.mem [1005] : 
                         (N22)? \nz.mem [1179] : 
                         (N24)? \nz.mem [1353] : 1'b0;
  assign r_data_o[134] = (N17)? \nz.mem [134] : 
                         (N19)? \nz.mem [308] : 
                         (N21)? \nz.mem [482] : 
                         (N23)? \nz.mem [656] : 
                         (N18)? \nz.mem [830] : 
                         (N20)? \nz.mem [1004] : 
                         (N22)? \nz.mem [1178] : 
                         (N24)? \nz.mem [1352] : 1'b0;
  assign r_data_o[133] = (N17)? \nz.mem [133] : 
                         (N19)? \nz.mem [307] : 
                         (N21)? \nz.mem [481] : 
                         (N23)? \nz.mem [655] : 
                         (N18)? \nz.mem [829] : 
                         (N20)? \nz.mem [1003] : 
                         (N22)? \nz.mem [1177] : 
                         (N24)? \nz.mem [1351] : 1'b0;
  assign r_data_o[132] = (N17)? \nz.mem [132] : 
                         (N19)? \nz.mem [306] : 
                         (N21)? \nz.mem [480] : 
                         (N23)? \nz.mem [654] : 
                         (N18)? \nz.mem [828] : 
                         (N20)? \nz.mem [1002] : 
                         (N22)? \nz.mem [1176] : 
                         (N24)? \nz.mem [1350] : 1'b0;
  assign r_data_o[131] = (N17)? \nz.mem [131] : 
                         (N19)? \nz.mem [305] : 
                         (N21)? \nz.mem [479] : 
                         (N23)? \nz.mem [653] : 
                         (N18)? \nz.mem [827] : 
                         (N20)? \nz.mem [1001] : 
                         (N22)? \nz.mem [1175] : 
                         (N24)? \nz.mem [1349] : 1'b0;
  assign r_data_o[130] = (N17)? \nz.mem [130] : 
                         (N19)? \nz.mem [304] : 
                         (N21)? \nz.mem [478] : 
                         (N23)? \nz.mem [652] : 
                         (N18)? \nz.mem [826] : 
                         (N20)? \nz.mem [1000] : 
                         (N22)? \nz.mem [1174] : 
                         (N24)? \nz.mem [1348] : 1'b0;
  assign r_data_o[129] = (N17)? \nz.mem [129] : 
                         (N19)? \nz.mem [303] : 
                         (N21)? \nz.mem [477] : 
                         (N23)? \nz.mem [651] : 
                         (N18)? \nz.mem [825] : 
                         (N20)? \nz.mem [999] : 
                         (N22)? \nz.mem [1173] : 
                         (N24)? \nz.mem [1347] : 1'b0;
  assign r_data_o[128] = (N17)? \nz.mem [128] : 
                         (N19)? \nz.mem [302] : 
                         (N21)? \nz.mem [476] : 
                         (N23)? \nz.mem [650] : 
                         (N18)? \nz.mem [824] : 
                         (N20)? \nz.mem [998] : 
                         (N22)? \nz.mem [1172] : 
                         (N24)? \nz.mem [1346] : 1'b0;
  assign r_data_o[127] = (N17)? \nz.mem [127] : 
                         (N19)? \nz.mem [301] : 
                         (N21)? \nz.mem [475] : 
                         (N23)? \nz.mem [649] : 
                         (N18)? \nz.mem [823] : 
                         (N20)? \nz.mem [997] : 
                         (N22)? \nz.mem [1171] : 
                         (N24)? \nz.mem [1345] : 1'b0;
  assign r_data_o[126] = (N17)? \nz.mem [126] : 
                         (N19)? \nz.mem [300] : 
                         (N21)? \nz.mem [474] : 
                         (N23)? \nz.mem [648] : 
                         (N18)? \nz.mem [822] : 
                         (N20)? \nz.mem [996] : 
                         (N22)? \nz.mem [1170] : 
                         (N24)? \nz.mem [1344] : 1'b0;
  assign r_data_o[125] = (N17)? \nz.mem [125] : 
                         (N19)? \nz.mem [299] : 
                         (N21)? \nz.mem [473] : 
                         (N23)? \nz.mem [647] : 
                         (N18)? \nz.mem [821] : 
                         (N20)? \nz.mem [995] : 
                         (N22)? \nz.mem [1169] : 
                         (N24)? \nz.mem [1343] : 1'b0;
  assign r_data_o[124] = (N17)? \nz.mem [124] : 
                         (N19)? \nz.mem [298] : 
                         (N21)? \nz.mem [472] : 
                         (N23)? \nz.mem [646] : 
                         (N18)? \nz.mem [820] : 
                         (N20)? \nz.mem [994] : 
                         (N22)? \nz.mem [1168] : 
                         (N24)? \nz.mem [1342] : 1'b0;
  assign r_data_o[123] = (N17)? \nz.mem [123] : 
                         (N19)? \nz.mem [297] : 
                         (N21)? \nz.mem [471] : 
                         (N23)? \nz.mem [645] : 
                         (N18)? \nz.mem [819] : 
                         (N20)? \nz.mem [993] : 
                         (N22)? \nz.mem [1167] : 
                         (N24)? \nz.mem [1341] : 1'b0;
  assign r_data_o[122] = (N17)? \nz.mem [122] : 
                         (N19)? \nz.mem [296] : 
                         (N21)? \nz.mem [470] : 
                         (N23)? \nz.mem [644] : 
                         (N18)? \nz.mem [818] : 
                         (N20)? \nz.mem [992] : 
                         (N22)? \nz.mem [1166] : 
                         (N24)? \nz.mem [1340] : 1'b0;
  assign r_data_o[121] = (N17)? \nz.mem [121] : 
                         (N19)? \nz.mem [295] : 
                         (N21)? \nz.mem [469] : 
                         (N23)? \nz.mem [643] : 
                         (N18)? \nz.mem [817] : 
                         (N20)? \nz.mem [991] : 
                         (N22)? \nz.mem [1165] : 
                         (N24)? \nz.mem [1339] : 1'b0;
  assign r_data_o[120] = (N17)? \nz.mem [120] : 
                         (N19)? \nz.mem [294] : 
                         (N21)? \nz.mem [468] : 
                         (N23)? \nz.mem [642] : 
                         (N18)? \nz.mem [816] : 
                         (N20)? \nz.mem [990] : 
                         (N22)? \nz.mem [1164] : 
                         (N24)? \nz.mem [1338] : 1'b0;
  assign r_data_o[119] = (N17)? \nz.mem [119] : 
                         (N19)? \nz.mem [293] : 
                         (N21)? \nz.mem [467] : 
                         (N23)? \nz.mem [641] : 
                         (N18)? \nz.mem [815] : 
                         (N20)? \nz.mem [989] : 
                         (N22)? \nz.mem [1163] : 
                         (N24)? \nz.mem [1337] : 1'b0;
  assign r_data_o[118] = (N17)? \nz.mem [118] : 
                         (N19)? \nz.mem [292] : 
                         (N21)? \nz.mem [466] : 
                         (N23)? \nz.mem [640] : 
                         (N18)? \nz.mem [814] : 
                         (N20)? \nz.mem [988] : 
                         (N22)? \nz.mem [1162] : 
                         (N24)? \nz.mem [1336] : 1'b0;
  assign r_data_o[117] = (N17)? \nz.mem [117] : 
                         (N19)? \nz.mem [291] : 
                         (N21)? \nz.mem [465] : 
                         (N23)? \nz.mem [639] : 
                         (N18)? \nz.mem [813] : 
                         (N20)? \nz.mem [987] : 
                         (N22)? \nz.mem [1161] : 
                         (N24)? \nz.mem [1335] : 1'b0;
  assign r_data_o[116] = (N17)? \nz.mem [116] : 
                         (N19)? \nz.mem [290] : 
                         (N21)? \nz.mem [464] : 
                         (N23)? \nz.mem [638] : 
                         (N18)? \nz.mem [812] : 
                         (N20)? \nz.mem [986] : 
                         (N22)? \nz.mem [1160] : 
                         (N24)? \nz.mem [1334] : 1'b0;
  assign r_data_o[115] = (N17)? \nz.mem [115] : 
                         (N19)? \nz.mem [289] : 
                         (N21)? \nz.mem [463] : 
                         (N23)? \nz.mem [637] : 
                         (N18)? \nz.mem [811] : 
                         (N20)? \nz.mem [985] : 
                         (N22)? \nz.mem [1159] : 
                         (N24)? \nz.mem [1333] : 1'b0;
  assign r_data_o[114] = (N17)? \nz.mem [114] : 
                         (N19)? \nz.mem [288] : 
                         (N21)? \nz.mem [462] : 
                         (N23)? \nz.mem [636] : 
                         (N18)? \nz.mem [810] : 
                         (N20)? \nz.mem [984] : 
                         (N22)? \nz.mem [1158] : 
                         (N24)? \nz.mem [1332] : 1'b0;
  assign r_data_o[113] = (N17)? \nz.mem [113] : 
                         (N19)? \nz.mem [287] : 
                         (N21)? \nz.mem [461] : 
                         (N23)? \nz.mem [635] : 
                         (N18)? \nz.mem [809] : 
                         (N20)? \nz.mem [983] : 
                         (N22)? \nz.mem [1157] : 
                         (N24)? \nz.mem [1331] : 1'b0;
  assign r_data_o[112] = (N17)? \nz.mem [112] : 
                         (N19)? \nz.mem [286] : 
                         (N21)? \nz.mem [460] : 
                         (N23)? \nz.mem [634] : 
                         (N18)? \nz.mem [808] : 
                         (N20)? \nz.mem [982] : 
                         (N22)? \nz.mem [1156] : 
                         (N24)? \nz.mem [1330] : 1'b0;
  assign r_data_o[111] = (N17)? \nz.mem [111] : 
                         (N19)? \nz.mem [285] : 
                         (N21)? \nz.mem [459] : 
                         (N23)? \nz.mem [633] : 
                         (N18)? \nz.mem [807] : 
                         (N20)? \nz.mem [981] : 
                         (N22)? \nz.mem [1155] : 
                         (N24)? \nz.mem [1329] : 1'b0;
  assign r_data_o[110] = (N17)? \nz.mem [110] : 
                         (N19)? \nz.mem [284] : 
                         (N21)? \nz.mem [458] : 
                         (N23)? \nz.mem [632] : 
                         (N18)? \nz.mem [806] : 
                         (N20)? \nz.mem [980] : 
                         (N22)? \nz.mem [1154] : 
                         (N24)? \nz.mem [1328] : 1'b0;
  assign r_data_o[109] = (N17)? \nz.mem [109] : 
                         (N19)? \nz.mem [283] : 
                         (N21)? \nz.mem [457] : 
                         (N23)? \nz.mem [631] : 
                         (N18)? \nz.mem [805] : 
                         (N20)? \nz.mem [979] : 
                         (N22)? \nz.mem [1153] : 
                         (N24)? \nz.mem [1327] : 1'b0;
  assign r_data_o[108] = (N17)? \nz.mem [108] : 
                         (N19)? \nz.mem [282] : 
                         (N21)? \nz.mem [456] : 
                         (N23)? \nz.mem [630] : 
                         (N18)? \nz.mem [804] : 
                         (N20)? \nz.mem [978] : 
                         (N22)? \nz.mem [1152] : 
                         (N24)? \nz.mem [1326] : 1'b0;
  assign r_data_o[107] = (N17)? \nz.mem [107] : 
                         (N19)? \nz.mem [281] : 
                         (N21)? \nz.mem [455] : 
                         (N23)? \nz.mem [629] : 
                         (N18)? \nz.mem [803] : 
                         (N20)? \nz.mem [977] : 
                         (N22)? \nz.mem [1151] : 
                         (N24)? \nz.mem [1325] : 1'b0;
  assign r_data_o[106] = (N17)? \nz.mem [106] : 
                         (N19)? \nz.mem [280] : 
                         (N21)? \nz.mem [454] : 
                         (N23)? \nz.mem [628] : 
                         (N18)? \nz.mem [802] : 
                         (N20)? \nz.mem [976] : 
                         (N22)? \nz.mem [1150] : 
                         (N24)? \nz.mem [1324] : 1'b0;
  assign r_data_o[105] = (N17)? \nz.mem [105] : 
                         (N19)? \nz.mem [279] : 
                         (N21)? \nz.mem [453] : 
                         (N23)? \nz.mem [627] : 
                         (N18)? \nz.mem [801] : 
                         (N20)? \nz.mem [975] : 
                         (N22)? \nz.mem [1149] : 
                         (N24)? \nz.mem [1323] : 1'b0;
  assign r_data_o[104] = (N17)? \nz.mem [104] : 
                         (N19)? \nz.mem [278] : 
                         (N21)? \nz.mem [452] : 
                         (N23)? \nz.mem [626] : 
                         (N18)? \nz.mem [800] : 
                         (N20)? \nz.mem [974] : 
                         (N22)? \nz.mem [1148] : 
                         (N24)? \nz.mem [1322] : 1'b0;
  assign r_data_o[103] = (N17)? \nz.mem [103] : 
                         (N19)? \nz.mem [277] : 
                         (N21)? \nz.mem [451] : 
                         (N23)? \nz.mem [625] : 
                         (N18)? \nz.mem [799] : 
                         (N20)? \nz.mem [973] : 
                         (N22)? \nz.mem [1147] : 
                         (N24)? \nz.mem [1321] : 1'b0;
  assign r_data_o[102] = (N17)? \nz.mem [102] : 
                         (N19)? \nz.mem [276] : 
                         (N21)? \nz.mem [450] : 
                         (N23)? \nz.mem [624] : 
                         (N18)? \nz.mem [798] : 
                         (N20)? \nz.mem [972] : 
                         (N22)? \nz.mem [1146] : 
                         (N24)? \nz.mem [1320] : 1'b0;
  assign r_data_o[101] = (N17)? \nz.mem [101] : 
                         (N19)? \nz.mem [275] : 
                         (N21)? \nz.mem [449] : 
                         (N23)? \nz.mem [623] : 
                         (N18)? \nz.mem [797] : 
                         (N20)? \nz.mem [971] : 
                         (N22)? \nz.mem [1145] : 
                         (N24)? \nz.mem [1319] : 1'b0;
  assign r_data_o[100] = (N17)? \nz.mem [100] : 
                         (N19)? \nz.mem [274] : 
                         (N21)? \nz.mem [448] : 
                         (N23)? \nz.mem [622] : 
                         (N18)? \nz.mem [796] : 
                         (N20)? \nz.mem [970] : 
                         (N22)? \nz.mem [1144] : 
                         (N24)? \nz.mem [1318] : 1'b0;
  assign r_data_o[99] = (N17)? \nz.mem [99] : 
                        (N19)? \nz.mem [273] : 
                        (N21)? \nz.mem [447] : 
                        (N23)? \nz.mem [621] : 
                        (N18)? \nz.mem [795] : 
                        (N20)? \nz.mem [969] : 
                        (N22)? \nz.mem [1143] : 
                        (N24)? \nz.mem [1317] : 1'b0;
  assign r_data_o[98] = (N17)? \nz.mem [98] : 
                        (N19)? \nz.mem [272] : 
                        (N21)? \nz.mem [446] : 
                        (N23)? \nz.mem [620] : 
                        (N18)? \nz.mem [794] : 
                        (N20)? \nz.mem [968] : 
                        (N22)? \nz.mem [1142] : 
                        (N24)? \nz.mem [1316] : 1'b0;
  assign r_data_o[97] = (N17)? \nz.mem [97] : 
                        (N19)? \nz.mem [271] : 
                        (N21)? \nz.mem [445] : 
                        (N23)? \nz.mem [619] : 
                        (N18)? \nz.mem [793] : 
                        (N20)? \nz.mem [967] : 
                        (N22)? \nz.mem [1141] : 
                        (N24)? \nz.mem [1315] : 1'b0;
  assign r_data_o[96] = (N17)? \nz.mem [96] : 
                        (N19)? \nz.mem [270] : 
                        (N21)? \nz.mem [444] : 
                        (N23)? \nz.mem [618] : 
                        (N18)? \nz.mem [792] : 
                        (N20)? \nz.mem [966] : 
                        (N22)? \nz.mem [1140] : 
                        (N24)? \nz.mem [1314] : 1'b0;
  assign r_data_o[95] = (N17)? \nz.mem [95] : 
                        (N19)? \nz.mem [269] : 
                        (N21)? \nz.mem [443] : 
                        (N23)? \nz.mem [617] : 
                        (N18)? \nz.mem [791] : 
                        (N20)? \nz.mem [965] : 
                        (N22)? \nz.mem [1139] : 
                        (N24)? \nz.mem [1313] : 1'b0;
  assign r_data_o[94] = (N17)? \nz.mem [94] : 
                        (N19)? \nz.mem [268] : 
                        (N21)? \nz.mem [442] : 
                        (N23)? \nz.mem [616] : 
                        (N18)? \nz.mem [790] : 
                        (N20)? \nz.mem [964] : 
                        (N22)? \nz.mem [1138] : 
                        (N24)? \nz.mem [1312] : 1'b0;
  assign r_data_o[93] = (N17)? \nz.mem [93] : 
                        (N19)? \nz.mem [267] : 
                        (N21)? \nz.mem [441] : 
                        (N23)? \nz.mem [615] : 
                        (N18)? \nz.mem [789] : 
                        (N20)? \nz.mem [963] : 
                        (N22)? \nz.mem [1137] : 
                        (N24)? \nz.mem [1311] : 1'b0;
  assign r_data_o[92] = (N17)? \nz.mem [92] : 
                        (N19)? \nz.mem [266] : 
                        (N21)? \nz.mem [440] : 
                        (N23)? \nz.mem [614] : 
                        (N18)? \nz.mem [788] : 
                        (N20)? \nz.mem [962] : 
                        (N22)? \nz.mem [1136] : 
                        (N24)? \nz.mem [1310] : 1'b0;
  assign r_data_o[91] = (N17)? \nz.mem [91] : 
                        (N19)? \nz.mem [265] : 
                        (N21)? \nz.mem [439] : 
                        (N23)? \nz.mem [613] : 
                        (N18)? \nz.mem [787] : 
                        (N20)? \nz.mem [961] : 
                        (N22)? \nz.mem [1135] : 
                        (N24)? \nz.mem [1309] : 1'b0;
  assign r_data_o[90] = (N17)? \nz.mem [90] : 
                        (N19)? \nz.mem [264] : 
                        (N21)? \nz.mem [438] : 
                        (N23)? \nz.mem [612] : 
                        (N18)? \nz.mem [786] : 
                        (N20)? \nz.mem [960] : 
                        (N22)? \nz.mem [1134] : 
                        (N24)? \nz.mem [1308] : 1'b0;
  assign r_data_o[89] = (N17)? \nz.mem [89] : 
                        (N19)? \nz.mem [263] : 
                        (N21)? \nz.mem [437] : 
                        (N23)? \nz.mem [611] : 
                        (N18)? \nz.mem [785] : 
                        (N20)? \nz.mem [959] : 
                        (N22)? \nz.mem [1133] : 
                        (N24)? \nz.mem [1307] : 1'b0;
  assign r_data_o[88] = (N17)? \nz.mem [88] : 
                        (N19)? \nz.mem [262] : 
                        (N21)? \nz.mem [436] : 
                        (N23)? \nz.mem [610] : 
                        (N18)? \nz.mem [784] : 
                        (N20)? \nz.mem [958] : 
                        (N22)? \nz.mem [1132] : 
                        (N24)? \nz.mem [1306] : 1'b0;
  assign r_data_o[87] = (N17)? \nz.mem [87] : 
                        (N19)? \nz.mem [261] : 
                        (N21)? \nz.mem [435] : 
                        (N23)? \nz.mem [609] : 
                        (N18)? \nz.mem [783] : 
                        (N20)? \nz.mem [957] : 
                        (N22)? \nz.mem [1131] : 
                        (N24)? \nz.mem [1305] : 1'b0;
  assign r_data_o[86] = (N17)? \nz.mem [86] : 
                        (N19)? \nz.mem [260] : 
                        (N21)? \nz.mem [434] : 
                        (N23)? \nz.mem [608] : 
                        (N18)? \nz.mem [782] : 
                        (N20)? \nz.mem [956] : 
                        (N22)? \nz.mem [1130] : 
                        (N24)? \nz.mem [1304] : 1'b0;
  assign r_data_o[85] = (N17)? \nz.mem [85] : 
                        (N19)? \nz.mem [259] : 
                        (N21)? \nz.mem [433] : 
                        (N23)? \nz.mem [607] : 
                        (N18)? \nz.mem [781] : 
                        (N20)? \nz.mem [955] : 
                        (N22)? \nz.mem [1129] : 
                        (N24)? \nz.mem [1303] : 1'b0;
  assign r_data_o[84] = (N17)? \nz.mem [84] : 
                        (N19)? \nz.mem [258] : 
                        (N21)? \nz.mem [432] : 
                        (N23)? \nz.mem [606] : 
                        (N18)? \nz.mem [780] : 
                        (N20)? \nz.mem [954] : 
                        (N22)? \nz.mem [1128] : 
                        (N24)? \nz.mem [1302] : 1'b0;
  assign r_data_o[83] = (N17)? \nz.mem [83] : 
                        (N19)? \nz.mem [257] : 
                        (N21)? \nz.mem [431] : 
                        (N23)? \nz.mem [605] : 
                        (N18)? \nz.mem [779] : 
                        (N20)? \nz.mem [953] : 
                        (N22)? \nz.mem [1127] : 
                        (N24)? \nz.mem [1301] : 1'b0;
  assign r_data_o[82] = (N17)? \nz.mem [82] : 
                        (N19)? \nz.mem [256] : 
                        (N21)? \nz.mem [430] : 
                        (N23)? \nz.mem [604] : 
                        (N18)? \nz.mem [778] : 
                        (N20)? \nz.mem [952] : 
                        (N22)? \nz.mem [1126] : 
                        (N24)? \nz.mem [1300] : 1'b0;
  assign r_data_o[81] = (N17)? \nz.mem [81] : 
                        (N19)? \nz.mem [255] : 
                        (N21)? \nz.mem [429] : 
                        (N23)? \nz.mem [603] : 
                        (N18)? \nz.mem [777] : 
                        (N20)? \nz.mem [951] : 
                        (N22)? \nz.mem [1125] : 
                        (N24)? \nz.mem [1299] : 1'b0;
  assign r_data_o[80] = (N17)? \nz.mem [80] : 
                        (N19)? \nz.mem [254] : 
                        (N21)? \nz.mem [428] : 
                        (N23)? \nz.mem [602] : 
                        (N18)? \nz.mem [776] : 
                        (N20)? \nz.mem [950] : 
                        (N22)? \nz.mem [1124] : 
                        (N24)? \nz.mem [1298] : 1'b0;
  assign r_data_o[79] = (N17)? \nz.mem [79] : 
                        (N19)? \nz.mem [253] : 
                        (N21)? \nz.mem [427] : 
                        (N23)? \nz.mem [601] : 
                        (N18)? \nz.mem [775] : 
                        (N20)? \nz.mem [949] : 
                        (N22)? \nz.mem [1123] : 
                        (N24)? \nz.mem [1297] : 1'b0;
  assign r_data_o[78] = (N17)? \nz.mem [78] : 
                        (N19)? \nz.mem [252] : 
                        (N21)? \nz.mem [426] : 
                        (N23)? \nz.mem [600] : 
                        (N18)? \nz.mem [774] : 
                        (N20)? \nz.mem [948] : 
                        (N22)? \nz.mem [1122] : 
                        (N24)? \nz.mem [1296] : 1'b0;
  assign r_data_o[77] = (N17)? \nz.mem [77] : 
                        (N19)? \nz.mem [251] : 
                        (N21)? \nz.mem [425] : 
                        (N23)? \nz.mem [599] : 
                        (N18)? \nz.mem [773] : 
                        (N20)? \nz.mem [947] : 
                        (N22)? \nz.mem [1121] : 
                        (N24)? \nz.mem [1295] : 1'b0;
  assign r_data_o[76] = (N17)? \nz.mem [76] : 
                        (N19)? \nz.mem [250] : 
                        (N21)? \nz.mem [424] : 
                        (N23)? \nz.mem [598] : 
                        (N18)? \nz.mem [772] : 
                        (N20)? \nz.mem [946] : 
                        (N22)? \nz.mem [1120] : 
                        (N24)? \nz.mem [1294] : 1'b0;
  assign r_data_o[75] = (N17)? \nz.mem [75] : 
                        (N19)? \nz.mem [249] : 
                        (N21)? \nz.mem [423] : 
                        (N23)? \nz.mem [597] : 
                        (N18)? \nz.mem [771] : 
                        (N20)? \nz.mem [945] : 
                        (N22)? \nz.mem [1119] : 
                        (N24)? \nz.mem [1293] : 1'b0;
  assign r_data_o[74] = (N17)? \nz.mem [74] : 
                        (N19)? \nz.mem [248] : 
                        (N21)? \nz.mem [422] : 
                        (N23)? \nz.mem [596] : 
                        (N18)? \nz.mem [770] : 
                        (N20)? \nz.mem [944] : 
                        (N22)? \nz.mem [1118] : 
                        (N24)? \nz.mem [1292] : 1'b0;
  assign r_data_o[73] = (N17)? \nz.mem [73] : 
                        (N19)? \nz.mem [247] : 
                        (N21)? \nz.mem [421] : 
                        (N23)? \nz.mem [595] : 
                        (N18)? \nz.mem [769] : 
                        (N20)? \nz.mem [943] : 
                        (N22)? \nz.mem [1117] : 
                        (N24)? \nz.mem [1291] : 1'b0;
  assign r_data_o[72] = (N17)? \nz.mem [72] : 
                        (N19)? \nz.mem [246] : 
                        (N21)? \nz.mem [420] : 
                        (N23)? \nz.mem [594] : 
                        (N18)? \nz.mem [768] : 
                        (N20)? \nz.mem [942] : 
                        (N22)? \nz.mem [1116] : 
                        (N24)? \nz.mem [1290] : 1'b0;
  assign r_data_o[71] = (N17)? \nz.mem [71] : 
                        (N19)? \nz.mem [245] : 
                        (N21)? \nz.mem [419] : 
                        (N23)? \nz.mem [593] : 
                        (N18)? \nz.mem [767] : 
                        (N20)? \nz.mem [941] : 
                        (N22)? \nz.mem [1115] : 
                        (N24)? \nz.mem [1289] : 1'b0;
  assign r_data_o[70] = (N17)? \nz.mem [70] : 
                        (N19)? \nz.mem [244] : 
                        (N21)? \nz.mem [418] : 
                        (N23)? \nz.mem [592] : 
                        (N18)? \nz.mem [766] : 
                        (N20)? \nz.mem [940] : 
                        (N22)? \nz.mem [1114] : 
                        (N24)? \nz.mem [1288] : 1'b0;
  assign r_data_o[69] = (N17)? \nz.mem [69] : 
                        (N19)? \nz.mem [243] : 
                        (N21)? \nz.mem [417] : 
                        (N23)? \nz.mem [591] : 
                        (N18)? \nz.mem [765] : 
                        (N20)? \nz.mem [939] : 
                        (N22)? \nz.mem [1113] : 
                        (N24)? \nz.mem [1287] : 1'b0;
  assign r_data_o[68] = (N17)? \nz.mem [68] : 
                        (N19)? \nz.mem [242] : 
                        (N21)? \nz.mem [416] : 
                        (N23)? \nz.mem [590] : 
                        (N18)? \nz.mem [764] : 
                        (N20)? \nz.mem [938] : 
                        (N22)? \nz.mem [1112] : 
                        (N24)? \nz.mem [1286] : 1'b0;
  assign r_data_o[67] = (N17)? \nz.mem [67] : 
                        (N19)? \nz.mem [241] : 
                        (N21)? \nz.mem [415] : 
                        (N23)? \nz.mem [589] : 
                        (N18)? \nz.mem [763] : 
                        (N20)? \nz.mem [937] : 
                        (N22)? \nz.mem [1111] : 
                        (N24)? \nz.mem [1285] : 1'b0;
  assign r_data_o[66] = (N17)? \nz.mem [66] : 
                        (N19)? \nz.mem [240] : 
                        (N21)? \nz.mem [414] : 
                        (N23)? \nz.mem [588] : 
                        (N18)? \nz.mem [762] : 
                        (N20)? \nz.mem [936] : 
                        (N22)? \nz.mem [1110] : 
                        (N24)? \nz.mem [1284] : 1'b0;
  assign r_data_o[65] = (N17)? \nz.mem [65] : 
                        (N19)? \nz.mem [239] : 
                        (N21)? \nz.mem [413] : 
                        (N23)? \nz.mem [587] : 
                        (N18)? \nz.mem [761] : 
                        (N20)? \nz.mem [935] : 
                        (N22)? \nz.mem [1109] : 
                        (N24)? \nz.mem [1283] : 1'b0;
  assign r_data_o[64] = (N17)? \nz.mem [64] : 
                        (N19)? \nz.mem [238] : 
                        (N21)? \nz.mem [412] : 
                        (N23)? \nz.mem [586] : 
                        (N18)? \nz.mem [760] : 
                        (N20)? \nz.mem [934] : 
                        (N22)? \nz.mem [1108] : 
                        (N24)? \nz.mem [1282] : 1'b0;
  assign r_data_o[63] = (N17)? \nz.mem [63] : 
                        (N19)? \nz.mem [237] : 
                        (N21)? \nz.mem [411] : 
                        (N23)? \nz.mem [585] : 
                        (N18)? \nz.mem [759] : 
                        (N20)? \nz.mem [933] : 
                        (N22)? \nz.mem [1107] : 
                        (N24)? \nz.mem [1281] : 1'b0;
  assign r_data_o[62] = (N17)? \nz.mem [62] : 
                        (N19)? \nz.mem [236] : 
                        (N21)? \nz.mem [410] : 
                        (N23)? \nz.mem [584] : 
                        (N18)? \nz.mem [758] : 
                        (N20)? \nz.mem [932] : 
                        (N22)? \nz.mem [1106] : 
                        (N24)? \nz.mem [1280] : 1'b0;
  assign r_data_o[61] = (N17)? \nz.mem [61] : 
                        (N19)? \nz.mem [235] : 
                        (N21)? \nz.mem [409] : 
                        (N23)? \nz.mem [583] : 
                        (N18)? \nz.mem [757] : 
                        (N20)? \nz.mem [931] : 
                        (N22)? \nz.mem [1105] : 
                        (N24)? \nz.mem [1279] : 1'b0;
  assign r_data_o[60] = (N17)? \nz.mem [60] : 
                        (N19)? \nz.mem [234] : 
                        (N21)? \nz.mem [408] : 
                        (N23)? \nz.mem [582] : 
                        (N18)? \nz.mem [756] : 
                        (N20)? \nz.mem [930] : 
                        (N22)? \nz.mem [1104] : 
                        (N24)? \nz.mem [1278] : 1'b0;
  assign r_data_o[59] = (N17)? \nz.mem [59] : 
                        (N19)? \nz.mem [233] : 
                        (N21)? \nz.mem [407] : 
                        (N23)? \nz.mem [581] : 
                        (N18)? \nz.mem [755] : 
                        (N20)? \nz.mem [929] : 
                        (N22)? \nz.mem [1103] : 
                        (N24)? \nz.mem [1277] : 1'b0;
  assign r_data_o[58] = (N17)? \nz.mem [58] : 
                        (N19)? \nz.mem [232] : 
                        (N21)? \nz.mem [406] : 
                        (N23)? \nz.mem [580] : 
                        (N18)? \nz.mem [754] : 
                        (N20)? \nz.mem [928] : 
                        (N22)? \nz.mem [1102] : 
                        (N24)? \nz.mem [1276] : 1'b0;
  assign r_data_o[57] = (N17)? \nz.mem [57] : 
                        (N19)? \nz.mem [231] : 
                        (N21)? \nz.mem [405] : 
                        (N23)? \nz.mem [579] : 
                        (N18)? \nz.mem [753] : 
                        (N20)? \nz.mem [927] : 
                        (N22)? \nz.mem [1101] : 
                        (N24)? \nz.mem [1275] : 1'b0;
  assign r_data_o[56] = (N17)? \nz.mem [56] : 
                        (N19)? \nz.mem [230] : 
                        (N21)? \nz.mem [404] : 
                        (N23)? \nz.mem [578] : 
                        (N18)? \nz.mem [752] : 
                        (N20)? \nz.mem [926] : 
                        (N22)? \nz.mem [1100] : 
                        (N24)? \nz.mem [1274] : 1'b0;
  assign r_data_o[55] = (N17)? \nz.mem [55] : 
                        (N19)? \nz.mem [229] : 
                        (N21)? \nz.mem [403] : 
                        (N23)? \nz.mem [577] : 
                        (N18)? \nz.mem [751] : 
                        (N20)? \nz.mem [925] : 
                        (N22)? \nz.mem [1099] : 
                        (N24)? \nz.mem [1273] : 1'b0;
  assign r_data_o[54] = (N17)? \nz.mem [54] : 
                        (N19)? \nz.mem [228] : 
                        (N21)? \nz.mem [402] : 
                        (N23)? \nz.mem [576] : 
                        (N18)? \nz.mem [750] : 
                        (N20)? \nz.mem [924] : 
                        (N22)? \nz.mem [1098] : 
                        (N24)? \nz.mem [1272] : 1'b0;
  assign r_data_o[53] = (N17)? \nz.mem [53] : 
                        (N19)? \nz.mem [227] : 
                        (N21)? \nz.mem [401] : 
                        (N23)? \nz.mem [575] : 
                        (N18)? \nz.mem [749] : 
                        (N20)? \nz.mem [923] : 
                        (N22)? \nz.mem [1097] : 
                        (N24)? \nz.mem [1271] : 1'b0;
  assign r_data_o[52] = (N17)? \nz.mem [52] : 
                        (N19)? \nz.mem [226] : 
                        (N21)? \nz.mem [400] : 
                        (N23)? \nz.mem [574] : 
                        (N18)? \nz.mem [748] : 
                        (N20)? \nz.mem [922] : 
                        (N22)? \nz.mem [1096] : 
                        (N24)? \nz.mem [1270] : 1'b0;
  assign r_data_o[51] = (N17)? \nz.mem [51] : 
                        (N19)? \nz.mem [225] : 
                        (N21)? \nz.mem [399] : 
                        (N23)? \nz.mem [573] : 
                        (N18)? \nz.mem [747] : 
                        (N20)? \nz.mem [921] : 
                        (N22)? \nz.mem [1095] : 
                        (N24)? \nz.mem [1269] : 1'b0;
  assign r_data_o[50] = (N17)? \nz.mem [50] : 
                        (N19)? \nz.mem [224] : 
                        (N21)? \nz.mem [398] : 
                        (N23)? \nz.mem [572] : 
                        (N18)? \nz.mem [746] : 
                        (N20)? \nz.mem [920] : 
                        (N22)? \nz.mem [1094] : 
                        (N24)? \nz.mem [1268] : 1'b0;
  assign r_data_o[49] = (N17)? \nz.mem [49] : 
                        (N19)? \nz.mem [223] : 
                        (N21)? \nz.mem [397] : 
                        (N23)? \nz.mem [571] : 
                        (N18)? \nz.mem [745] : 
                        (N20)? \nz.mem [919] : 
                        (N22)? \nz.mem [1093] : 
                        (N24)? \nz.mem [1267] : 1'b0;
  assign r_data_o[48] = (N17)? \nz.mem [48] : 
                        (N19)? \nz.mem [222] : 
                        (N21)? \nz.mem [396] : 
                        (N23)? \nz.mem [570] : 
                        (N18)? \nz.mem [744] : 
                        (N20)? \nz.mem [918] : 
                        (N22)? \nz.mem [1092] : 
                        (N24)? \nz.mem [1266] : 1'b0;
  assign r_data_o[47] = (N17)? \nz.mem [47] : 
                        (N19)? \nz.mem [221] : 
                        (N21)? \nz.mem [395] : 
                        (N23)? \nz.mem [569] : 
                        (N18)? \nz.mem [743] : 
                        (N20)? \nz.mem [917] : 
                        (N22)? \nz.mem [1091] : 
                        (N24)? \nz.mem [1265] : 1'b0;
  assign r_data_o[46] = (N17)? \nz.mem [46] : 
                        (N19)? \nz.mem [220] : 
                        (N21)? \nz.mem [394] : 
                        (N23)? \nz.mem [568] : 
                        (N18)? \nz.mem [742] : 
                        (N20)? \nz.mem [916] : 
                        (N22)? \nz.mem [1090] : 
                        (N24)? \nz.mem [1264] : 1'b0;
  assign r_data_o[45] = (N17)? \nz.mem [45] : 
                        (N19)? \nz.mem [219] : 
                        (N21)? \nz.mem [393] : 
                        (N23)? \nz.mem [567] : 
                        (N18)? \nz.mem [741] : 
                        (N20)? \nz.mem [915] : 
                        (N22)? \nz.mem [1089] : 
                        (N24)? \nz.mem [1263] : 1'b0;
  assign r_data_o[44] = (N17)? \nz.mem [44] : 
                        (N19)? \nz.mem [218] : 
                        (N21)? \nz.mem [392] : 
                        (N23)? \nz.mem [566] : 
                        (N18)? \nz.mem [740] : 
                        (N20)? \nz.mem [914] : 
                        (N22)? \nz.mem [1088] : 
                        (N24)? \nz.mem [1262] : 1'b0;
  assign r_data_o[43] = (N17)? \nz.mem [43] : 
                        (N19)? \nz.mem [217] : 
                        (N21)? \nz.mem [391] : 
                        (N23)? \nz.mem [565] : 
                        (N18)? \nz.mem [739] : 
                        (N20)? \nz.mem [913] : 
                        (N22)? \nz.mem [1087] : 
                        (N24)? \nz.mem [1261] : 1'b0;
  assign r_data_o[42] = (N17)? \nz.mem [42] : 
                        (N19)? \nz.mem [216] : 
                        (N21)? \nz.mem [390] : 
                        (N23)? \nz.mem [564] : 
                        (N18)? \nz.mem [738] : 
                        (N20)? \nz.mem [912] : 
                        (N22)? \nz.mem [1086] : 
                        (N24)? \nz.mem [1260] : 1'b0;
  assign r_data_o[41] = (N17)? \nz.mem [41] : 
                        (N19)? \nz.mem [215] : 
                        (N21)? \nz.mem [389] : 
                        (N23)? \nz.mem [563] : 
                        (N18)? \nz.mem [737] : 
                        (N20)? \nz.mem [911] : 
                        (N22)? \nz.mem [1085] : 
                        (N24)? \nz.mem [1259] : 1'b0;
  assign r_data_o[40] = (N17)? \nz.mem [40] : 
                        (N19)? \nz.mem [214] : 
                        (N21)? \nz.mem [388] : 
                        (N23)? \nz.mem [562] : 
                        (N18)? \nz.mem [736] : 
                        (N20)? \nz.mem [910] : 
                        (N22)? \nz.mem [1084] : 
                        (N24)? \nz.mem [1258] : 1'b0;
  assign r_data_o[39] = (N17)? \nz.mem [39] : 
                        (N19)? \nz.mem [213] : 
                        (N21)? \nz.mem [387] : 
                        (N23)? \nz.mem [561] : 
                        (N18)? \nz.mem [735] : 
                        (N20)? \nz.mem [909] : 
                        (N22)? \nz.mem [1083] : 
                        (N24)? \nz.mem [1257] : 1'b0;
  assign r_data_o[38] = (N17)? \nz.mem [38] : 
                        (N19)? \nz.mem [212] : 
                        (N21)? \nz.mem [386] : 
                        (N23)? \nz.mem [560] : 
                        (N18)? \nz.mem [734] : 
                        (N20)? \nz.mem [908] : 
                        (N22)? \nz.mem [1082] : 
                        (N24)? \nz.mem [1256] : 1'b0;
  assign r_data_o[37] = (N17)? \nz.mem [37] : 
                        (N19)? \nz.mem [211] : 
                        (N21)? \nz.mem [385] : 
                        (N23)? \nz.mem [559] : 
                        (N18)? \nz.mem [733] : 
                        (N20)? \nz.mem [907] : 
                        (N22)? \nz.mem [1081] : 
                        (N24)? \nz.mem [1255] : 1'b0;
  assign r_data_o[36] = (N17)? \nz.mem [36] : 
                        (N19)? \nz.mem [210] : 
                        (N21)? \nz.mem [384] : 
                        (N23)? \nz.mem [558] : 
                        (N18)? \nz.mem [732] : 
                        (N20)? \nz.mem [906] : 
                        (N22)? \nz.mem [1080] : 
                        (N24)? \nz.mem [1254] : 1'b0;
  assign r_data_o[35] = (N17)? \nz.mem [35] : 
                        (N19)? \nz.mem [209] : 
                        (N21)? \nz.mem [383] : 
                        (N23)? \nz.mem [557] : 
                        (N18)? \nz.mem [731] : 
                        (N20)? \nz.mem [905] : 
                        (N22)? \nz.mem [1079] : 
                        (N24)? \nz.mem [1253] : 1'b0;
  assign r_data_o[34] = (N17)? \nz.mem [34] : 
                        (N19)? \nz.mem [208] : 
                        (N21)? \nz.mem [382] : 
                        (N23)? \nz.mem [556] : 
                        (N18)? \nz.mem [730] : 
                        (N20)? \nz.mem [904] : 
                        (N22)? \nz.mem [1078] : 
                        (N24)? \nz.mem [1252] : 1'b0;
  assign r_data_o[33] = (N17)? \nz.mem [33] : 
                        (N19)? \nz.mem [207] : 
                        (N21)? \nz.mem [381] : 
                        (N23)? \nz.mem [555] : 
                        (N18)? \nz.mem [729] : 
                        (N20)? \nz.mem [903] : 
                        (N22)? \nz.mem [1077] : 
                        (N24)? \nz.mem [1251] : 1'b0;
  assign r_data_o[32] = (N17)? \nz.mem [32] : 
                        (N19)? \nz.mem [206] : 
                        (N21)? \nz.mem [380] : 
                        (N23)? \nz.mem [554] : 
                        (N18)? \nz.mem [728] : 
                        (N20)? \nz.mem [902] : 
                        (N22)? \nz.mem [1076] : 
                        (N24)? \nz.mem [1250] : 1'b0;
  assign r_data_o[31] = (N17)? \nz.mem [31] : 
                        (N19)? \nz.mem [205] : 
                        (N21)? \nz.mem [379] : 
                        (N23)? \nz.mem [553] : 
                        (N18)? \nz.mem [727] : 
                        (N20)? \nz.mem [901] : 
                        (N22)? \nz.mem [1075] : 
                        (N24)? \nz.mem [1249] : 1'b0;
  assign r_data_o[30] = (N17)? \nz.mem [30] : 
                        (N19)? \nz.mem [204] : 
                        (N21)? \nz.mem [378] : 
                        (N23)? \nz.mem [552] : 
                        (N18)? \nz.mem [726] : 
                        (N20)? \nz.mem [900] : 
                        (N22)? \nz.mem [1074] : 
                        (N24)? \nz.mem [1248] : 1'b0;
  assign r_data_o[29] = (N17)? \nz.mem [29] : 
                        (N19)? \nz.mem [203] : 
                        (N21)? \nz.mem [377] : 
                        (N23)? \nz.mem [551] : 
                        (N18)? \nz.mem [725] : 
                        (N20)? \nz.mem [899] : 
                        (N22)? \nz.mem [1073] : 
                        (N24)? \nz.mem [1247] : 1'b0;
  assign r_data_o[28] = (N17)? \nz.mem [28] : 
                        (N19)? \nz.mem [202] : 
                        (N21)? \nz.mem [376] : 
                        (N23)? \nz.mem [550] : 
                        (N18)? \nz.mem [724] : 
                        (N20)? \nz.mem [898] : 
                        (N22)? \nz.mem [1072] : 
                        (N24)? \nz.mem [1246] : 1'b0;
  assign r_data_o[27] = (N17)? \nz.mem [27] : 
                        (N19)? \nz.mem [201] : 
                        (N21)? \nz.mem [375] : 
                        (N23)? \nz.mem [549] : 
                        (N18)? \nz.mem [723] : 
                        (N20)? \nz.mem [897] : 
                        (N22)? \nz.mem [1071] : 
                        (N24)? \nz.mem [1245] : 1'b0;
  assign r_data_o[26] = (N17)? \nz.mem [26] : 
                        (N19)? \nz.mem [200] : 
                        (N21)? \nz.mem [374] : 
                        (N23)? \nz.mem [548] : 
                        (N18)? \nz.mem [722] : 
                        (N20)? \nz.mem [896] : 
                        (N22)? \nz.mem [1070] : 
                        (N24)? \nz.mem [1244] : 1'b0;
  assign r_data_o[25] = (N17)? \nz.mem [25] : 
                        (N19)? \nz.mem [199] : 
                        (N21)? \nz.mem [373] : 
                        (N23)? \nz.mem [547] : 
                        (N18)? \nz.mem [721] : 
                        (N20)? \nz.mem [895] : 
                        (N22)? \nz.mem [1069] : 
                        (N24)? \nz.mem [1243] : 1'b0;
  assign r_data_o[24] = (N17)? \nz.mem [24] : 
                        (N19)? \nz.mem [198] : 
                        (N21)? \nz.mem [372] : 
                        (N23)? \nz.mem [546] : 
                        (N18)? \nz.mem [720] : 
                        (N20)? \nz.mem [894] : 
                        (N22)? \nz.mem [1068] : 
                        (N24)? \nz.mem [1242] : 1'b0;
  assign r_data_o[23] = (N17)? \nz.mem [23] : 
                        (N19)? \nz.mem [197] : 
                        (N21)? \nz.mem [371] : 
                        (N23)? \nz.mem [545] : 
                        (N18)? \nz.mem [719] : 
                        (N20)? \nz.mem [893] : 
                        (N22)? \nz.mem [1067] : 
                        (N24)? \nz.mem [1241] : 1'b0;
  assign r_data_o[22] = (N17)? \nz.mem [22] : 
                        (N19)? \nz.mem [196] : 
                        (N21)? \nz.mem [370] : 
                        (N23)? \nz.mem [544] : 
                        (N18)? \nz.mem [718] : 
                        (N20)? \nz.mem [892] : 
                        (N22)? \nz.mem [1066] : 
                        (N24)? \nz.mem [1240] : 1'b0;
  assign r_data_o[21] = (N17)? \nz.mem [21] : 
                        (N19)? \nz.mem [195] : 
                        (N21)? \nz.mem [369] : 
                        (N23)? \nz.mem [543] : 
                        (N18)? \nz.mem [717] : 
                        (N20)? \nz.mem [891] : 
                        (N22)? \nz.mem [1065] : 
                        (N24)? \nz.mem [1239] : 1'b0;
  assign r_data_o[20] = (N17)? \nz.mem [20] : 
                        (N19)? \nz.mem [194] : 
                        (N21)? \nz.mem [368] : 
                        (N23)? \nz.mem [542] : 
                        (N18)? \nz.mem [716] : 
                        (N20)? \nz.mem [890] : 
                        (N22)? \nz.mem [1064] : 
                        (N24)? \nz.mem [1238] : 1'b0;
  assign r_data_o[19] = (N17)? \nz.mem [19] : 
                        (N19)? \nz.mem [193] : 
                        (N21)? \nz.mem [367] : 
                        (N23)? \nz.mem [541] : 
                        (N18)? \nz.mem [715] : 
                        (N20)? \nz.mem [889] : 
                        (N22)? \nz.mem [1063] : 
                        (N24)? \nz.mem [1237] : 1'b0;
  assign r_data_o[18] = (N17)? \nz.mem [18] : 
                        (N19)? \nz.mem [192] : 
                        (N21)? \nz.mem [366] : 
                        (N23)? \nz.mem [540] : 
                        (N18)? \nz.mem [714] : 
                        (N20)? \nz.mem [888] : 
                        (N22)? \nz.mem [1062] : 
                        (N24)? \nz.mem [1236] : 1'b0;
  assign r_data_o[17] = (N17)? \nz.mem [17] : 
                        (N19)? \nz.mem [191] : 
                        (N21)? \nz.mem [365] : 
                        (N23)? \nz.mem [539] : 
                        (N18)? \nz.mem [713] : 
                        (N20)? \nz.mem [887] : 
                        (N22)? \nz.mem [1061] : 
                        (N24)? \nz.mem [1235] : 1'b0;
  assign r_data_o[16] = (N17)? \nz.mem [16] : 
                        (N19)? \nz.mem [190] : 
                        (N21)? \nz.mem [364] : 
                        (N23)? \nz.mem [538] : 
                        (N18)? \nz.mem [712] : 
                        (N20)? \nz.mem [886] : 
                        (N22)? \nz.mem [1060] : 
                        (N24)? \nz.mem [1234] : 1'b0;
  assign r_data_o[15] = (N17)? \nz.mem [15] : 
                        (N19)? \nz.mem [189] : 
                        (N21)? \nz.mem [363] : 
                        (N23)? \nz.mem [537] : 
                        (N18)? \nz.mem [711] : 
                        (N20)? \nz.mem [885] : 
                        (N22)? \nz.mem [1059] : 
                        (N24)? \nz.mem [1233] : 1'b0;
  assign r_data_o[14] = (N17)? \nz.mem [14] : 
                        (N19)? \nz.mem [188] : 
                        (N21)? \nz.mem [362] : 
                        (N23)? \nz.mem [536] : 
                        (N18)? \nz.mem [710] : 
                        (N20)? \nz.mem [884] : 
                        (N22)? \nz.mem [1058] : 
                        (N24)? \nz.mem [1232] : 1'b0;
  assign r_data_o[13] = (N17)? \nz.mem [13] : 
                        (N19)? \nz.mem [187] : 
                        (N21)? \nz.mem [361] : 
                        (N23)? \nz.mem [535] : 
                        (N18)? \nz.mem [709] : 
                        (N20)? \nz.mem [883] : 
                        (N22)? \nz.mem [1057] : 
                        (N24)? \nz.mem [1231] : 1'b0;
  assign r_data_o[12] = (N17)? \nz.mem [12] : 
                        (N19)? \nz.mem [186] : 
                        (N21)? \nz.mem [360] : 
                        (N23)? \nz.mem [534] : 
                        (N18)? \nz.mem [708] : 
                        (N20)? \nz.mem [882] : 
                        (N22)? \nz.mem [1056] : 
                        (N24)? \nz.mem [1230] : 1'b0;
  assign r_data_o[11] = (N17)? \nz.mem [11] : 
                        (N19)? \nz.mem [185] : 
                        (N21)? \nz.mem [359] : 
                        (N23)? \nz.mem [533] : 
                        (N18)? \nz.mem [707] : 
                        (N20)? \nz.mem [881] : 
                        (N22)? \nz.mem [1055] : 
                        (N24)? \nz.mem [1229] : 1'b0;
  assign r_data_o[10] = (N17)? \nz.mem [10] : 
                        (N19)? \nz.mem [184] : 
                        (N21)? \nz.mem [358] : 
                        (N23)? \nz.mem [532] : 
                        (N18)? \nz.mem [706] : 
                        (N20)? \nz.mem [880] : 
                        (N22)? \nz.mem [1054] : 
                        (N24)? \nz.mem [1228] : 1'b0;
  assign r_data_o[9] = (N17)? \nz.mem [9] : 
                       (N19)? \nz.mem [183] : 
                       (N21)? \nz.mem [357] : 
                       (N23)? \nz.mem [531] : 
                       (N18)? \nz.mem [705] : 
                       (N20)? \nz.mem [879] : 
                       (N22)? \nz.mem [1053] : 
                       (N24)? \nz.mem [1227] : 1'b0;
  assign r_data_o[8] = (N17)? \nz.mem [8] : 
                       (N19)? \nz.mem [182] : 
                       (N21)? \nz.mem [356] : 
                       (N23)? \nz.mem [530] : 
                       (N18)? \nz.mem [704] : 
                       (N20)? \nz.mem [878] : 
                       (N22)? \nz.mem [1052] : 
                       (N24)? \nz.mem [1226] : 1'b0;
  assign r_data_o[7] = (N17)? \nz.mem [7] : 
                       (N19)? \nz.mem [181] : 
                       (N21)? \nz.mem [355] : 
                       (N23)? \nz.mem [529] : 
                       (N18)? \nz.mem [703] : 
                       (N20)? \nz.mem [877] : 
                       (N22)? \nz.mem [1051] : 
                       (N24)? \nz.mem [1225] : 1'b0;
  assign r_data_o[6] = (N17)? \nz.mem [6] : 
                       (N19)? \nz.mem [180] : 
                       (N21)? \nz.mem [354] : 
                       (N23)? \nz.mem [528] : 
                       (N18)? \nz.mem [702] : 
                       (N20)? \nz.mem [876] : 
                       (N22)? \nz.mem [1050] : 
                       (N24)? \nz.mem [1224] : 1'b0;
  assign r_data_o[5] = (N17)? \nz.mem [5] : 
                       (N19)? \nz.mem [179] : 
                       (N21)? \nz.mem [353] : 
                       (N23)? \nz.mem [527] : 
                       (N18)? \nz.mem [701] : 
                       (N20)? \nz.mem [875] : 
                       (N22)? \nz.mem [1049] : 
                       (N24)? \nz.mem [1223] : 1'b0;
  assign r_data_o[4] = (N17)? \nz.mem [4] : 
                       (N19)? \nz.mem [178] : 
                       (N21)? \nz.mem [352] : 
                       (N23)? \nz.mem [526] : 
                       (N18)? \nz.mem [700] : 
                       (N20)? \nz.mem [874] : 
                       (N22)? \nz.mem [1048] : 
                       (N24)? \nz.mem [1222] : 1'b0;
  assign r_data_o[3] = (N17)? \nz.mem [3] : 
                       (N19)? \nz.mem [177] : 
                       (N21)? \nz.mem [351] : 
                       (N23)? \nz.mem [525] : 
                       (N18)? \nz.mem [699] : 
                       (N20)? \nz.mem [873] : 
                       (N22)? \nz.mem [1047] : 
                       (N24)? \nz.mem [1221] : 1'b0;
  assign r_data_o[2] = (N17)? \nz.mem [2] : 
                       (N19)? \nz.mem [176] : 
                       (N21)? \nz.mem [350] : 
                       (N23)? \nz.mem [524] : 
                       (N18)? \nz.mem [698] : 
                       (N20)? \nz.mem [872] : 
                       (N22)? \nz.mem [1046] : 
                       (N24)? \nz.mem [1220] : 1'b0;
  assign r_data_o[1] = (N17)? \nz.mem [1] : 
                       (N19)? \nz.mem [175] : 
                       (N21)? \nz.mem [349] : 
                       (N23)? \nz.mem [523] : 
                       (N18)? \nz.mem [697] : 
                       (N20)? \nz.mem [871] : 
                       (N22)? \nz.mem [1045] : 
                       (N24)? \nz.mem [1219] : 1'b0;
  assign r_data_o[0] = (N17)? \nz.mem [0] : 
                       (N19)? \nz.mem [174] : 
                       (N21)? \nz.mem [348] : 
                       (N23)? \nz.mem [522] : 
                       (N18)? \nz.mem [696] : 
                       (N20)? \nz.mem [870] : 
                       (N22)? \nz.mem [1044] : 
                       (N24)? \nz.mem [1218] : 1'b0;
  assign N50 = w_addr_i[0] & w_addr_i[1];
  assign N33 = N50 & w_addr_i[2];
  assign N51 = N0 & w_addr_i[1];
  assign N0 = ~w_addr_i[0];
  assign N32 = N51 & w_addr_i[2];
  assign N52 = w_addr_i[0] & N1;
  assign N1 = ~w_addr_i[1];
  assign N31 = N52 & w_addr_i[2];
  assign N53 = N2 & N3;
  assign N2 = ~w_addr_i[0];
  assign N3 = ~w_addr_i[1];
  assign N30 = N53 & w_addr_i[2];
  assign N29 = N50 & N4;
  assign N4 = ~w_addr_i[2];
  assign N28 = N51 & N5;
  assign N5 = ~w_addr_i[2];
  assign N27 = N52 & N6;
  assign N6 = ~w_addr_i[2];
  assign N26 = N53 & N7;
  assign N7 = ~w_addr_i[2];
  assign { N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34 } = (N8)? { N33, N33, N32, N32, N31, N31, N30, N30, N29, N29, N28, N28, N27, N27, N26, N26 } : 
                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N25;
  assign N10 = ~r_addr_i[0];
  assign N11 = ~r_addr_i[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r_addr_i[1];
  assign N14 = r_addr_i[0] & N11;
  assign N15 = r_addr_i[0] & r_addr_i[1];
  assign N16 = ~r_addr_i[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r_addr_i[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r_addr_i[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r_addr_i[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r_addr_i[2];
  assign N25 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N48) begin
      \nz.mem_1391_sv2v_reg  <= w_data_i[173];
      \nz.mem_1390_sv2v_reg  <= w_data_i[172];
      \nz.mem_1389_sv2v_reg  <= w_data_i[171];
      \nz.mem_1388_sv2v_reg  <= w_data_i[170];
      \nz.mem_1387_sv2v_reg  <= w_data_i[169];
      \nz.mem_1386_sv2v_reg  <= w_data_i[168];
      \nz.mem_1385_sv2v_reg  <= w_data_i[167];
      \nz.mem_1384_sv2v_reg  <= w_data_i[166];
      \nz.mem_1383_sv2v_reg  <= w_data_i[165];
      \nz.mem_1382_sv2v_reg  <= w_data_i[164];
      \nz.mem_1381_sv2v_reg  <= w_data_i[163];
      \nz.mem_1380_sv2v_reg  <= w_data_i[162];
      \nz.mem_1379_sv2v_reg  <= w_data_i[161];
      \nz.mem_1378_sv2v_reg  <= w_data_i[160];
      \nz.mem_1377_sv2v_reg  <= w_data_i[159];
      \nz.mem_1376_sv2v_reg  <= w_data_i[158];
      \nz.mem_1375_sv2v_reg  <= w_data_i[157];
      \nz.mem_1374_sv2v_reg  <= w_data_i[156];
      \nz.mem_1373_sv2v_reg  <= w_data_i[155];
      \nz.mem_1372_sv2v_reg  <= w_data_i[154];
      \nz.mem_1371_sv2v_reg  <= w_data_i[153];
      \nz.mem_1370_sv2v_reg  <= w_data_i[152];
      \nz.mem_1369_sv2v_reg  <= w_data_i[151];
      \nz.mem_1368_sv2v_reg  <= w_data_i[150];
      \nz.mem_1367_sv2v_reg  <= w_data_i[149];
      \nz.mem_1366_sv2v_reg  <= w_data_i[148];
      \nz.mem_1365_sv2v_reg  <= w_data_i[147];
      \nz.mem_1364_sv2v_reg  <= w_data_i[146];
      \nz.mem_1363_sv2v_reg  <= w_data_i[145];
      \nz.mem_1362_sv2v_reg  <= w_data_i[144];
      \nz.mem_1361_sv2v_reg  <= w_data_i[143];
      \nz.mem_1360_sv2v_reg  <= w_data_i[142];
      \nz.mem_1359_sv2v_reg  <= w_data_i[141];
      \nz.mem_1358_sv2v_reg  <= w_data_i[140];
      \nz.mem_1357_sv2v_reg  <= w_data_i[139];
      \nz.mem_1356_sv2v_reg  <= w_data_i[138];
      \nz.mem_1355_sv2v_reg  <= w_data_i[137];
      \nz.mem_1354_sv2v_reg  <= w_data_i[136];
      \nz.mem_1353_sv2v_reg  <= w_data_i[135];
      \nz.mem_1352_sv2v_reg  <= w_data_i[134];
      \nz.mem_1351_sv2v_reg  <= w_data_i[133];
      \nz.mem_1350_sv2v_reg  <= w_data_i[132];
      \nz.mem_1349_sv2v_reg  <= w_data_i[131];
      \nz.mem_1348_sv2v_reg  <= w_data_i[130];
      \nz.mem_1347_sv2v_reg  <= w_data_i[129];
      \nz.mem_1346_sv2v_reg  <= w_data_i[128];
      \nz.mem_1345_sv2v_reg  <= w_data_i[127];
      \nz.mem_1344_sv2v_reg  <= w_data_i[126];
      \nz.mem_1343_sv2v_reg  <= w_data_i[125];
      \nz.mem_1342_sv2v_reg  <= w_data_i[124];
      \nz.mem_1341_sv2v_reg  <= w_data_i[123];
      \nz.mem_1340_sv2v_reg  <= w_data_i[122];
      \nz.mem_1339_sv2v_reg  <= w_data_i[121];
      \nz.mem_1338_sv2v_reg  <= w_data_i[120];
      \nz.mem_1337_sv2v_reg  <= w_data_i[119];
      \nz.mem_1336_sv2v_reg  <= w_data_i[118];
      \nz.mem_1335_sv2v_reg  <= w_data_i[117];
      \nz.mem_1334_sv2v_reg  <= w_data_i[116];
      \nz.mem_1333_sv2v_reg  <= w_data_i[115];
      \nz.mem_1332_sv2v_reg  <= w_data_i[114];
      \nz.mem_1331_sv2v_reg  <= w_data_i[113];
      \nz.mem_1330_sv2v_reg  <= w_data_i[112];
      \nz.mem_1329_sv2v_reg  <= w_data_i[111];
      \nz.mem_1328_sv2v_reg  <= w_data_i[110];
      \nz.mem_1327_sv2v_reg  <= w_data_i[109];
      \nz.mem_1326_sv2v_reg  <= w_data_i[108];
      \nz.mem_1325_sv2v_reg  <= w_data_i[107];
      \nz.mem_1324_sv2v_reg  <= w_data_i[106];
      \nz.mem_1323_sv2v_reg  <= w_data_i[105];
      \nz.mem_1322_sv2v_reg  <= w_data_i[104];
      \nz.mem_1321_sv2v_reg  <= w_data_i[103];
      \nz.mem_1320_sv2v_reg  <= w_data_i[102];
      \nz.mem_1319_sv2v_reg  <= w_data_i[101];
      \nz.mem_1318_sv2v_reg  <= w_data_i[100];
      \nz.mem_1317_sv2v_reg  <= w_data_i[99];
      \nz.mem_1316_sv2v_reg  <= w_data_i[98];
      \nz.mem_1315_sv2v_reg  <= w_data_i[97];
      \nz.mem_1314_sv2v_reg  <= w_data_i[96];
      \nz.mem_1313_sv2v_reg  <= w_data_i[95];
      \nz.mem_1312_sv2v_reg  <= w_data_i[94];
      \nz.mem_1311_sv2v_reg  <= w_data_i[93];
      \nz.mem_1310_sv2v_reg  <= w_data_i[92];
      \nz.mem_1309_sv2v_reg  <= w_data_i[91];
      \nz.mem_1308_sv2v_reg  <= w_data_i[90];
      \nz.mem_1307_sv2v_reg  <= w_data_i[89];
      \nz.mem_1306_sv2v_reg  <= w_data_i[88];
      \nz.mem_1305_sv2v_reg  <= w_data_i[87];
      \nz.mem_1304_sv2v_reg  <= w_data_i[86];
      \nz.mem_1303_sv2v_reg  <= w_data_i[85];
      \nz.mem_1302_sv2v_reg  <= w_data_i[84];
      \nz.mem_1301_sv2v_reg  <= w_data_i[83];
      \nz.mem_1300_sv2v_reg  <= w_data_i[82];
      \nz.mem_1299_sv2v_reg  <= w_data_i[81];
      \nz.mem_1298_sv2v_reg  <= w_data_i[80];
      \nz.mem_1297_sv2v_reg  <= w_data_i[79];
      \nz.mem_1296_sv2v_reg  <= w_data_i[78];
      \nz.mem_1295_sv2v_reg  <= w_data_i[77];
      \nz.mem_1294_sv2v_reg  <= w_data_i[76];
      \nz.mem_1293_sv2v_reg  <= w_data_i[75];
      \nz.mem_1218_sv2v_reg  <= w_data_i[0];
    end 
    if(N49) begin
      \nz.mem_1292_sv2v_reg  <= w_data_i[74];
      \nz.mem_1291_sv2v_reg  <= w_data_i[73];
      \nz.mem_1290_sv2v_reg  <= w_data_i[72];
      \nz.mem_1289_sv2v_reg  <= w_data_i[71];
      \nz.mem_1288_sv2v_reg  <= w_data_i[70];
      \nz.mem_1287_sv2v_reg  <= w_data_i[69];
      \nz.mem_1286_sv2v_reg  <= w_data_i[68];
      \nz.mem_1285_sv2v_reg  <= w_data_i[67];
      \nz.mem_1284_sv2v_reg  <= w_data_i[66];
      \nz.mem_1283_sv2v_reg  <= w_data_i[65];
      \nz.mem_1282_sv2v_reg  <= w_data_i[64];
      \nz.mem_1281_sv2v_reg  <= w_data_i[63];
      \nz.mem_1280_sv2v_reg  <= w_data_i[62];
      \nz.mem_1279_sv2v_reg  <= w_data_i[61];
      \nz.mem_1278_sv2v_reg  <= w_data_i[60];
      \nz.mem_1277_sv2v_reg  <= w_data_i[59];
      \nz.mem_1276_sv2v_reg  <= w_data_i[58];
      \nz.mem_1275_sv2v_reg  <= w_data_i[57];
      \nz.mem_1274_sv2v_reg  <= w_data_i[56];
      \nz.mem_1273_sv2v_reg  <= w_data_i[55];
      \nz.mem_1272_sv2v_reg  <= w_data_i[54];
      \nz.mem_1271_sv2v_reg  <= w_data_i[53];
      \nz.mem_1270_sv2v_reg  <= w_data_i[52];
      \nz.mem_1269_sv2v_reg  <= w_data_i[51];
      \nz.mem_1268_sv2v_reg  <= w_data_i[50];
      \nz.mem_1267_sv2v_reg  <= w_data_i[49];
      \nz.mem_1266_sv2v_reg  <= w_data_i[48];
      \nz.mem_1265_sv2v_reg  <= w_data_i[47];
      \nz.mem_1264_sv2v_reg  <= w_data_i[46];
      \nz.mem_1263_sv2v_reg  <= w_data_i[45];
      \nz.mem_1262_sv2v_reg  <= w_data_i[44];
      \nz.mem_1261_sv2v_reg  <= w_data_i[43];
      \nz.mem_1260_sv2v_reg  <= w_data_i[42];
      \nz.mem_1259_sv2v_reg  <= w_data_i[41];
      \nz.mem_1258_sv2v_reg  <= w_data_i[40];
      \nz.mem_1257_sv2v_reg  <= w_data_i[39];
      \nz.mem_1256_sv2v_reg  <= w_data_i[38];
      \nz.mem_1255_sv2v_reg  <= w_data_i[37];
      \nz.mem_1254_sv2v_reg  <= w_data_i[36];
      \nz.mem_1253_sv2v_reg  <= w_data_i[35];
      \nz.mem_1252_sv2v_reg  <= w_data_i[34];
      \nz.mem_1251_sv2v_reg  <= w_data_i[33];
      \nz.mem_1250_sv2v_reg  <= w_data_i[32];
      \nz.mem_1249_sv2v_reg  <= w_data_i[31];
      \nz.mem_1248_sv2v_reg  <= w_data_i[30];
      \nz.mem_1247_sv2v_reg  <= w_data_i[29];
      \nz.mem_1246_sv2v_reg  <= w_data_i[28];
      \nz.mem_1245_sv2v_reg  <= w_data_i[27];
      \nz.mem_1244_sv2v_reg  <= w_data_i[26];
      \nz.mem_1243_sv2v_reg  <= w_data_i[25];
      \nz.mem_1242_sv2v_reg  <= w_data_i[24];
      \nz.mem_1241_sv2v_reg  <= w_data_i[23];
      \nz.mem_1240_sv2v_reg  <= w_data_i[22];
      \nz.mem_1239_sv2v_reg  <= w_data_i[21];
      \nz.mem_1238_sv2v_reg  <= w_data_i[20];
      \nz.mem_1237_sv2v_reg  <= w_data_i[19];
      \nz.mem_1236_sv2v_reg  <= w_data_i[18];
      \nz.mem_1235_sv2v_reg  <= w_data_i[17];
      \nz.mem_1234_sv2v_reg  <= w_data_i[16];
      \nz.mem_1233_sv2v_reg  <= w_data_i[15];
      \nz.mem_1232_sv2v_reg  <= w_data_i[14];
      \nz.mem_1231_sv2v_reg  <= w_data_i[13];
      \nz.mem_1230_sv2v_reg  <= w_data_i[12];
      \nz.mem_1229_sv2v_reg  <= w_data_i[11];
      \nz.mem_1228_sv2v_reg  <= w_data_i[10];
      \nz.mem_1227_sv2v_reg  <= w_data_i[9];
      \nz.mem_1226_sv2v_reg  <= w_data_i[8];
      \nz.mem_1225_sv2v_reg  <= w_data_i[7];
      \nz.mem_1224_sv2v_reg  <= w_data_i[6];
      \nz.mem_1223_sv2v_reg  <= w_data_i[5];
      \nz.mem_1222_sv2v_reg  <= w_data_i[4];
      \nz.mem_1221_sv2v_reg  <= w_data_i[3];
      \nz.mem_1220_sv2v_reg  <= w_data_i[2];
      \nz.mem_1219_sv2v_reg  <= w_data_i[1];
    end 
    if(N46) begin
      \nz.mem_1217_sv2v_reg  <= w_data_i[173];
      \nz.mem_1216_sv2v_reg  <= w_data_i[172];
      \nz.mem_1215_sv2v_reg  <= w_data_i[171];
      \nz.mem_1214_sv2v_reg  <= w_data_i[170];
      \nz.mem_1213_sv2v_reg  <= w_data_i[169];
      \nz.mem_1212_sv2v_reg  <= w_data_i[168];
      \nz.mem_1211_sv2v_reg  <= w_data_i[167];
      \nz.mem_1210_sv2v_reg  <= w_data_i[166];
      \nz.mem_1209_sv2v_reg  <= w_data_i[165];
      \nz.mem_1208_sv2v_reg  <= w_data_i[164];
      \nz.mem_1207_sv2v_reg  <= w_data_i[163];
      \nz.mem_1206_sv2v_reg  <= w_data_i[162];
      \nz.mem_1205_sv2v_reg  <= w_data_i[161];
      \nz.mem_1204_sv2v_reg  <= w_data_i[160];
      \nz.mem_1203_sv2v_reg  <= w_data_i[159];
      \nz.mem_1202_sv2v_reg  <= w_data_i[158];
      \nz.mem_1201_sv2v_reg  <= w_data_i[157];
      \nz.mem_1200_sv2v_reg  <= w_data_i[156];
      \nz.mem_1199_sv2v_reg  <= w_data_i[155];
      \nz.mem_1198_sv2v_reg  <= w_data_i[154];
      \nz.mem_1197_sv2v_reg  <= w_data_i[153];
      \nz.mem_1196_sv2v_reg  <= w_data_i[152];
      \nz.mem_1195_sv2v_reg  <= w_data_i[151];
      \nz.mem_1194_sv2v_reg  <= w_data_i[150];
      \nz.mem_1193_sv2v_reg  <= w_data_i[149];
      \nz.mem_1192_sv2v_reg  <= w_data_i[148];
      \nz.mem_1191_sv2v_reg  <= w_data_i[147];
      \nz.mem_1190_sv2v_reg  <= w_data_i[146];
      \nz.mem_1189_sv2v_reg  <= w_data_i[145];
      \nz.mem_1188_sv2v_reg  <= w_data_i[144];
      \nz.mem_1187_sv2v_reg  <= w_data_i[143];
      \nz.mem_1186_sv2v_reg  <= w_data_i[142];
      \nz.mem_1185_sv2v_reg  <= w_data_i[141];
      \nz.mem_1184_sv2v_reg  <= w_data_i[140];
      \nz.mem_1183_sv2v_reg  <= w_data_i[139];
      \nz.mem_1182_sv2v_reg  <= w_data_i[138];
      \nz.mem_1181_sv2v_reg  <= w_data_i[137];
      \nz.mem_1180_sv2v_reg  <= w_data_i[136];
      \nz.mem_1179_sv2v_reg  <= w_data_i[135];
      \nz.mem_1178_sv2v_reg  <= w_data_i[134];
      \nz.mem_1177_sv2v_reg  <= w_data_i[133];
      \nz.mem_1176_sv2v_reg  <= w_data_i[132];
      \nz.mem_1175_sv2v_reg  <= w_data_i[131];
      \nz.mem_1174_sv2v_reg  <= w_data_i[130];
      \nz.mem_1173_sv2v_reg  <= w_data_i[129];
      \nz.mem_1172_sv2v_reg  <= w_data_i[128];
      \nz.mem_1171_sv2v_reg  <= w_data_i[127];
      \nz.mem_1170_sv2v_reg  <= w_data_i[126];
      \nz.mem_1169_sv2v_reg  <= w_data_i[125];
      \nz.mem_1168_sv2v_reg  <= w_data_i[124];
      \nz.mem_1167_sv2v_reg  <= w_data_i[123];
      \nz.mem_1166_sv2v_reg  <= w_data_i[122];
      \nz.mem_1165_sv2v_reg  <= w_data_i[121];
      \nz.mem_1164_sv2v_reg  <= w_data_i[120];
      \nz.mem_1163_sv2v_reg  <= w_data_i[119];
      \nz.mem_1162_sv2v_reg  <= w_data_i[118];
      \nz.mem_1161_sv2v_reg  <= w_data_i[117];
      \nz.mem_1160_sv2v_reg  <= w_data_i[116];
      \nz.mem_1159_sv2v_reg  <= w_data_i[115];
      \nz.mem_1158_sv2v_reg  <= w_data_i[114];
      \nz.mem_1157_sv2v_reg  <= w_data_i[113];
      \nz.mem_1156_sv2v_reg  <= w_data_i[112];
      \nz.mem_1155_sv2v_reg  <= w_data_i[111];
      \nz.mem_1154_sv2v_reg  <= w_data_i[110];
      \nz.mem_1153_sv2v_reg  <= w_data_i[109];
      \nz.mem_1152_sv2v_reg  <= w_data_i[108];
      \nz.mem_1151_sv2v_reg  <= w_data_i[107];
      \nz.mem_1150_sv2v_reg  <= w_data_i[106];
      \nz.mem_1149_sv2v_reg  <= w_data_i[105];
      \nz.mem_1148_sv2v_reg  <= w_data_i[104];
      \nz.mem_1147_sv2v_reg  <= w_data_i[103];
      \nz.mem_1146_sv2v_reg  <= w_data_i[102];
      \nz.mem_1145_sv2v_reg  <= w_data_i[101];
      \nz.mem_1144_sv2v_reg  <= w_data_i[100];
      \nz.mem_1143_sv2v_reg  <= w_data_i[99];
      \nz.mem_1142_sv2v_reg  <= w_data_i[98];
      \nz.mem_1141_sv2v_reg  <= w_data_i[97];
      \nz.mem_1140_sv2v_reg  <= w_data_i[96];
      \nz.mem_1139_sv2v_reg  <= w_data_i[95];
      \nz.mem_1138_sv2v_reg  <= w_data_i[94];
      \nz.mem_1137_sv2v_reg  <= w_data_i[93];
      \nz.mem_1136_sv2v_reg  <= w_data_i[92];
      \nz.mem_1135_sv2v_reg  <= w_data_i[91];
      \nz.mem_1134_sv2v_reg  <= w_data_i[90];
      \nz.mem_1133_sv2v_reg  <= w_data_i[89];
      \nz.mem_1132_sv2v_reg  <= w_data_i[88];
      \nz.mem_1131_sv2v_reg  <= w_data_i[87];
      \nz.mem_1130_sv2v_reg  <= w_data_i[86];
      \nz.mem_1129_sv2v_reg  <= w_data_i[85];
      \nz.mem_1128_sv2v_reg  <= w_data_i[84];
      \nz.mem_1127_sv2v_reg  <= w_data_i[83];
      \nz.mem_1126_sv2v_reg  <= w_data_i[82];
      \nz.mem_1125_sv2v_reg  <= w_data_i[81];
      \nz.mem_1124_sv2v_reg  <= w_data_i[80];
      \nz.mem_1123_sv2v_reg  <= w_data_i[79];
      \nz.mem_1122_sv2v_reg  <= w_data_i[78];
      \nz.mem_1121_sv2v_reg  <= w_data_i[77];
      \nz.mem_1120_sv2v_reg  <= w_data_i[76];
      \nz.mem_1119_sv2v_reg  <= w_data_i[75];
      \nz.mem_1044_sv2v_reg  <= w_data_i[0];
    end 
    if(N47) begin
      \nz.mem_1118_sv2v_reg  <= w_data_i[74];
      \nz.mem_1117_sv2v_reg  <= w_data_i[73];
      \nz.mem_1116_sv2v_reg  <= w_data_i[72];
      \nz.mem_1115_sv2v_reg  <= w_data_i[71];
      \nz.mem_1114_sv2v_reg  <= w_data_i[70];
      \nz.mem_1113_sv2v_reg  <= w_data_i[69];
      \nz.mem_1112_sv2v_reg  <= w_data_i[68];
      \nz.mem_1111_sv2v_reg  <= w_data_i[67];
      \nz.mem_1110_sv2v_reg  <= w_data_i[66];
      \nz.mem_1109_sv2v_reg  <= w_data_i[65];
      \nz.mem_1108_sv2v_reg  <= w_data_i[64];
      \nz.mem_1107_sv2v_reg  <= w_data_i[63];
      \nz.mem_1106_sv2v_reg  <= w_data_i[62];
      \nz.mem_1105_sv2v_reg  <= w_data_i[61];
      \nz.mem_1104_sv2v_reg  <= w_data_i[60];
      \nz.mem_1103_sv2v_reg  <= w_data_i[59];
      \nz.mem_1102_sv2v_reg  <= w_data_i[58];
      \nz.mem_1101_sv2v_reg  <= w_data_i[57];
      \nz.mem_1100_sv2v_reg  <= w_data_i[56];
      \nz.mem_1099_sv2v_reg  <= w_data_i[55];
      \nz.mem_1098_sv2v_reg  <= w_data_i[54];
      \nz.mem_1097_sv2v_reg  <= w_data_i[53];
      \nz.mem_1096_sv2v_reg  <= w_data_i[52];
      \nz.mem_1095_sv2v_reg  <= w_data_i[51];
      \nz.mem_1094_sv2v_reg  <= w_data_i[50];
      \nz.mem_1093_sv2v_reg  <= w_data_i[49];
      \nz.mem_1092_sv2v_reg  <= w_data_i[48];
      \nz.mem_1091_sv2v_reg  <= w_data_i[47];
      \nz.mem_1090_sv2v_reg  <= w_data_i[46];
      \nz.mem_1089_sv2v_reg  <= w_data_i[45];
      \nz.mem_1088_sv2v_reg  <= w_data_i[44];
      \nz.mem_1087_sv2v_reg  <= w_data_i[43];
      \nz.mem_1086_sv2v_reg  <= w_data_i[42];
      \nz.mem_1085_sv2v_reg  <= w_data_i[41];
      \nz.mem_1084_sv2v_reg  <= w_data_i[40];
      \nz.mem_1083_sv2v_reg  <= w_data_i[39];
      \nz.mem_1082_sv2v_reg  <= w_data_i[38];
      \nz.mem_1081_sv2v_reg  <= w_data_i[37];
      \nz.mem_1080_sv2v_reg  <= w_data_i[36];
      \nz.mem_1079_sv2v_reg  <= w_data_i[35];
      \nz.mem_1078_sv2v_reg  <= w_data_i[34];
      \nz.mem_1077_sv2v_reg  <= w_data_i[33];
      \nz.mem_1076_sv2v_reg  <= w_data_i[32];
      \nz.mem_1075_sv2v_reg  <= w_data_i[31];
      \nz.mem_1074_sv2v_reg  <= w_data_i[30];
      \nz.mem_1073_sv2v_reg  <= w_data_i[29];
      \nz.mem_1072_sv2v_reg  <= w_data_i[28];
      \nz.mem_1071_sv2v_reg  <= w_data_i[27];
      \nz.mem_1070_sv2v_reg  <= w_data_i[26];
      \nz.mem_1069_sv2v_reg  <= w_data_i[25];
      \nz.mem_1068_sv2v_reg  <= w_data_i[24];
      \nz.mem_1067_sv2v_reg  <= w_data_i[23];
      \nz.mem_1066_sv2v_reg  <= w_data_i[22];
      \nz.mem_1065_sv2v_reg  <= w_data_i[21];
      \nz.mem_1064_sv2v_reg  <= w_data_i[20];
      \nz.mem_1063_sv2v_reg  <= w_data_i[19];
      \nz.mem_1062_sv2v_reg  <= w_data_i[18];
      \nz.mem_1061_sv2v_reg  <= w_data_i[17];
      \nz.mem_1060_sv2v_reg  <= w_data_i[16];
      \nz.mem_1059_sv2v_reg  <= w_data_i[15];
      \nz.mem_1058_sv2v_reg  <= w_data_i[14];
      \nz.mem_1057_sv2v_reg  <= w_data_i[13];
      \nz.mem_1056_sv2v_reg  <= w_data_i[12];
      \nz.mem_1055_sv2v_reg  <= w_data_i[11];
      \nz.mem_1054_sv2v_reg  <= w_data_i[10];
      \nz.mem_1053_sv2v_reg  <= w_data_i[9];
      \nz.mem_1052_sv2v_reg  <= w_data_i[8];
      \nz.mem_1051_sv2v_reg  <= w_data_i[7];
      \nz.mem_1050_sv2v_reg  <= w_data_i[6];
      \nz.mem_1049_sv2v_reg  <= w_data_i[5];
      \nz.mem_1048_sv2v_reg  <= w_data_i[4];
      \nz.mem_1047_sv2v_reg  <= w_data_i[3];
      \nz.mem_1046_sv2v_reg  <= w_data_i[2];
      \nz.mem_1045_sv2v_reg  <= w_data_i[1];
    end 
    if(N44) begin
      \nz.mem_1043_sv2v_reg  <= w_data_i[173];
      \nz.mem_1042_sv2v_reg  <= w_data_i[172];
      \nz.mem_1041_sv2v_reg  <= w_data_i[171];
      \nz.mem_1040_sv2v_reg  <= w_data_i[170];
      \nz.mem_1039_sv2v_reg  <= w_data_i[169];
      \nz.mem_1038_sv2v_reg  <= w_data_i[168];
      \nz.mem_1037_sv2v_reg  <= w_data_i[167];
      \nz.mem_1036_sv2v_reg  <= w_data_i[166];
      \nz.mem_1035_sv2v_reg  <= w_data_i[165];
      \nz.mem_1034_sv2v_reg  <= w_data_i[164];
      \nz.mem_1033_sv2v_reg  <= w_data_i[163];
      \nz.mem_1032_sv2v_reg  <= w_data_i[162];
      \nz.mem_1031_sv2v_reg  <= w_data_i[161];
      \nz.mem_1030_sv2v_reg  <= w_data_i[160];
      \nz.mem_1029_sv2v_reg  <= w_data_i[159];
      \nz.mem_1028_sv2v_reg  <= w_data_i[158];
      \nz.mem_1027_sv2v_reg  <= w_data_i[157];
      \nz.mem_1026_sv2v_reg  <= w_data_i[156];
      \nz.mem_1025_sv2v_reg  <= w_data_i[155];
      \nz.mem_1024_sv2v_reg  <= w_data_i[154];
      \nz.mem_1023_sv2v_reg  <= w_data_i[153];
      \nz.mem_1022_sv2v_reg  <= w_data_i[152];
      \nz.mem_1021_sv2v_reg  <= w_data_i[151];
      \nz.mem_1020_sv2v_reg  <= w_data_i[150];
      \nz.mem_1019_sv2v_reg  <= w_data_i[149];
      \nz.mem_1018_sv2v_reg  <= w_data_i[148];
      \nz.mem_1017_sv2v_reg  <= w_data_i[147];
      \nz.mem_1016_sv2v_reg  <= w_data_i[146];
      \nz.mem_1015_sv2v_reg  <= w_data_i[145];
      \nz.mem_1014_sv2v_reg  <= w_data_i[144];
      \nz.mem_1013_sv2v_reg  <= w_data_i[143];
      \nz.mem_1012_sv2v_reg  <= w_data_i[142];
      \nz.mem_1011_sv2v_reg  <= w_data_i[141];
      \nz.mem_1010_sv2v_reg  <= w_data_i[140];
      \nz.mem_1009_sv2v_reg  <= w_data_i[139];
      \nz.mem_1008_sv2v_reg  <= w_data_i[138];
      \nz.mem_1007_sv2v_reg  <= w_data_i[137];
      \nz.mem_1006_sv2v_reg  <= w_data_i[136];
      \nz.mem_1005_sv2v_reg  <= w_data_i[135];
      \nz.mem_1004_sv2v_reg  <= w_data_i[134];
      \nz.mem_1003_sv2v_reg  <= w_data_i[133];
      \nz.mem_1002_sv2v_reg  <= w_data_i[132];
      \nz.mem_1001_sv2v_reg  <= w_data_i[131];
      \nz.mem_1000_sv2v_reg  <= w_data_i[130];
      \nz.mem_999_sv2v_reg  <= w_data_i[129];
      \nz.mem_998_sv2v_reg  <= w_data_i[128];
      \nz.mem_997_sv2v_reg  <= w_data_i[127];
      \nz.mem_996_sv2v_reg  <= w_data_i[126];
      \nz.mem_995_sv2v_reg  <= w_data_i[125];
      \nz.mem_994_sv2v_reg  <= w_data_i[124];
      \nz.mem_993_sv2v_reg  <= w_data_i[123];
      \nz.mem_992_sv2v_reg  <= w_data_i[122];
      \nz.mem_991_sv2v_reg  <= w_data_i[121];
      \nz.mem_990_sv2v_reg  <= w_data_i[120];
      \nz.mem_989_sv2v_reg  <= w_data_i[119];
      \nz.mem_988_sv2v_reg  <= w_data_i[118];
      \nz.mem_987_sv2v_reg  <= w_data_i[117];
      \nz.mem_986_sv2v_reg  <= w_data_i[116];
      \nz.mem_985_sv2v_reg  <= w_data_i[115];
      \nz.mem_984_sv2v_reg  <= w_data_i[114];
      \nz.mem_983_sv2v_reg  <= w_data_i[113];
      \nz.mem_982_sv2v_reg  <= w_data_i[112];
      \nz.mem_981_sv2v_reg  <= w_data_i[111];
      \nz.mem_980_sv2v_reg  <= w_data_i[110];
      \nz.mem_979_sv2v_reg  <= w_data_i[109];
      \nz.mem_978_sv2v_reg  <= w_data_i[108];
      \nz.mem_977_sv2v_reg  <= w_data_i[107];
      \nz.mem_976_sv2v_reg  <= w_data_i[106];
      \nz.mem_975_sv2v_reg  <= w_data_i[105];
      \nz.mem_974_sv2v_reg  <= w_data_i[104];
      \nz.mem_973_sv2v_reg  <= w_data_i[103];
      \nz.mem_972_sv2v_reg  <= w_data_i[102];
      \nz.mem_971_sv2v_reg  <= w_data_i[101];
      \nz.mem_970_sv2v_reg  <= w_data_i[100];
      \nz.mem_969_sv2v_reg  <= w_data_i[99];
      \nz.mem_968_sv2v_reg  <= w_data_i[98];
      \nz.mem_967_sv2v_reg  <= w_data_i[97];
      \nz.mem_966_sv2v_reg  <= w_data_i[96];
      \nz.mem_965_sv2v_reg  <= w_data_i[95];
      \nz.mem_964_sv2v_reg  <= w_data_i[94];
      \nz.mem_963_sv2v_reg  <= w_data_i[93];
      \nz.mem_962_sv2v_reg  <= w_data_i[92];
      \nz.mem_961_sv2v_reg  <= w_data_i[91];
      \nz.mem_960_sv2v_reg  <= w_data_i[90];
      \nz.mem_959_sv2v_reg  <= w_data_i[89];
      \nz.mem_958_sv2v_reg  <= w_data_i[88];
      \nz.mem_957_sv2v_reg  <= w_data_i[87];
      \nz.mem_956_sv2v_reg  <= w_data_i[86];
      \nz.mem_955_sv2v_reg  <= w_data_i[85];
      \nz.mem_954_sv2v_reg  <= w_data_i[84];
      \nz.mem_953_sv2v_reg  <= w_data_i[83];
      \nz.mem_952_sv2v_reg  <= w_data_i[82];
      \nz.mem_951_sv2v_reg  <= w_data_i[81];
      \nz.mem_950_sv2v_reg  <= w_data_i[80];
      \nz.mem_949_sv2v_reg  <= w_data_i[79];
      \nz.mem_948_sv2v_reg  <= w_data_i[78];
      \nz.mem_947_sv2v_reg  <= w_data_i[77];
      \nz.mem_946_sv2v_reg  <= w_data_i[76];
      \nz.mem_945_sv2v_reg  <= w_data_i[75];
      \nz.mem_870_sv2v_reg  <= w_data_i[0];
    end 
    if(N45) begin
      \nz.mem_944_sv2v_reg  <= w_data_i[74];
      \nz.mem_943_sv2v_reg  <= w_data_i[73];
      \nz.mem_942_sv2v_reg  <= w_data_i[72];
      \nz.mem_941_sv2v_reg  <= w_data_i[71];
      \nz.mem_940_sv2v_reg  <= w_data_i[70];
      \nz.mem_939_sv2v_reg  <= w_data_i[69];
      \nz.mem_938_sv2v_reg  <= w_data_i[68];
      \nz.mem_937_sv2v_reg  <= w_data_i[67];
      \nz.mem_936_sv2v_reg  <= w_data_i[66];
      \nz.mem_935_sv2v_reg  <= w_data_i[65];
      \nz.mem_934_sv2v_reg  <= w_data_i[64];
      \nz.mem_933_sv2v_reg  <= w_data_i[63];
      \nz.mem_932_sv2v_reg  <= w_data_i[62];
      \nz.mem_931_sv2v_reg  <= w_data_i[61];
      \nz.mem_930_sv2v_reg  <= w_data_i[60];
      \nz.mem_929_sv2v_reg  <= w_data_i[59];
      \nz.mem_928_sv2v_reg  <= w_data_i[58];
      \nz.mem_927_sv2v_reg  <= w_data_i[57];
      \nz.mem_926_sv2v_reg  <= w_data_i[56];
      \nz.mem_925_sv2v_reg  <= w_data_i[55];
      \nz.mem_924_sv2v_reg  <= w_data_i[54];
      \nz.mem_923_sv2v_reg  <= w_data_i[53];
      \nz.mem_922_sv2v_reg  <= w_data_i[52];
      \nz.mem_921_sv2v_reg  <= w_data_i[51];
      \nz.mem_920_sv2v_reg  <= w_data_i[50];
      \nz.mem_919_sv2v_reg  <= w_data_i[49];
      \nz.mem_918_sv2v_reg  <= w_data_i[48];
      \nz.mem_917_sv2v_reg  <= w_data_i[47];
      \nz.mem_916_sv2v_reg  <= w_data_i[46];
      \nz.mem_915_sv2v_reg  <= w_data_i[45];
      \nz.mem_914_sv2v_reg  <= w_data_i[44];
      \nz.mem_913_sv2v_reg  <= w_data_i[43];
      \nz.mem_912_sv2v_reg  <= w_data_i[42];
      \nz.mem_911_sv2v_reg  <= w_data_i[41];
      \nz.mem_910_sv2v_reg  <= w_data_i[40];
      \nz.mem_909_sv2v_reg  <= w_data_i[39];
      \nz.mem_908_sv2v_reg  <= w_data_i[38];
      \nz.mem_907_sv2v_reg  <= w_data_i[37];
      \nz.mem_906_sv2v_reg  <= w_data_i[36];
      \nz.mem_905_sv2v_reg  <= w_data_i[35];
      \nz.mem_904_sv2v_reg  <= w_data_i[34];
      \nz.mem_903_sv2v_reg  <= w_data_i[33];
      \nz.mem_902_sv2v_reg  <= w_data_i[32];
      \nz.mem_901_sv2v_reg  <= w_data_i[31];
      \nz.mem_900_sv2v_reg  <= w_data_i[30];
      \nz.mem_899_sv2v_reg  <= w_data_i[29];
      \nz.mem_898_sv2v_reg  <= w_data_i[28];
      \nz.mem_897_sv2v_reg  <= w_data_i[27];
      \nz.mem_896_sv2v_reg  <= w_data_i[26];
      \nz.mem_895_sv2v_reg  <= w_data_i[25];
      \nz.mem_894_sv2v_reg  <= w_data_i[24];
      \nz.mem_893_sv2v_reg  <= w_data_i[23];
      \nz.mem_892_sv2v_reg  <= w_data_i[22];
      \nz.mem_891_sv2v_reg  <= w_data_i[21];
      \nz.mem_890_sv2v_reg  <= w_data_i[20];
      \nz.mem_889_sv2v_reg  <= w_data_i[19];
      \nz.mem_888_sv2v_reg  <= w_data_i[18];
      \nz.mem_887_sv2v_reg  <= w_data_i[17];
      \nz.mem_886_sv2v_reg  <= w_data_i[16];
      \nz.mem_885_sv2v_reg  <= w_data_i[15];
      \nz.mem_884_sv2v_reg  <= w_data_i[14];
      \nz.mem_883_sv2v_reg  <= w_data_i[13];
      \nz.mem_882_sv2v_reg  <= w_data_i[12];
      \nz.mem_881_sv2v_reg  <= w_data_i[11];
      \nz.mem_880_sv2v_reg  <= w_data_i[10];
      \nz.mem_879_sv2v_reg  <= w_data_i[9];
      \nz.mem_878_sv2v_reg  <= w_data_i[8];
      \nz.mem_877_sv2v_reg  <= w_data_i[7];
      \nz.mem_876_sv2v_reg  <= w_data_i[6];
      \nz.mem_875_sv2v_reg  <= w_data_i[5];
      \nz.mem_874_sv2v_reg  <= w_data_i[4];
      \nz.mem_873_sv2v_reg  <= w_data_i[3];
      \nz.mem_872_sv2v_reg  <= w_data_i[2];
      \nz.mem_871_sv2v_reg  <= w_data_i[1];
    end 
    if(N42) begin
      \nz.mem_869_sv2v_reg  <= w_data_i[173];
      \nz.mem_868_sv2v_reg  <= w_data_i[172];
      \nz.mem_867_sv2v_reg  <= w_data_i[171];
      \nz.mem_866_sv2v_reg  <= w_data_i[170];
      \nz.mem_865_sv2v_reg  <= w_data_i[169];
      \nz.mem_864_sv2v_reg  <= w_data_i[168];
      \nz.mem_863_sv2v_reg  <= w_data_i[167];
      \nz.mem_862_sv2v_reg  <= w_data_i[166];
      \nz.mem_861_sv2v_reg  <= w_data_i[165];
      \nz.mem_860_sv2v_reg  <= w_data_i[164];
      \nz.mem_859_sv2v_reg  <= w_data_i[163];
      \nz.mem_858_sv2v_reg  <= w_data_i[162];
      \nz.mem_857_sv2v_reg  <= w_data_i[161];
      \nz.mem_856_sv2v_reg  <= w_data_i[160];
      \nz.mem_855_sv2v_reg  <= w_data_i[159];
      \nz.mem_854_sv2v_reg  <= w_data_i[158];
      \nz.mem_853_sv2v_reg  <= w_data_i[157];
      \nz.mem_852_sv2v_reg  <= w_data_i[156];
      \nz.mem_851_sv2v_reg  <= w_data_i[155];
      \nz.mem_850_sv2v_reg  <= w_data_i[154];
      \nz.mem_849_sv2v_reg  <= w_data_i[153];
      \nz.mem_848_sv2v_reg  <= w_data_i[152];
      \nz.mem_847_sv2v_reg  <= w_data_i[151];
      \nz.mem_846_sv2v_reg  <= w_data_i[150];
      \nz.mem_845_sv2v_reg  <= w_data_i[149];
      \nz.mem_844_sv2v_reg  <= w_data_i[148];
      \nz.mem_843_sv2v_reg  <= w_data_i[147];
      \nz.mem_842_sv2v_reg  <= w_data_i[146];
      \nz.mem_841_sv2v_reg  <= w_data_i[145];
      \nz.mem_840_sv2v_reg  <= w_data_i[144];
      \nz.mem_839_sv2v_reg  <= w_data_i[143];
      \nz.mem_838_sv2v_reg  <= w_data_i[142];
      \nz.mem_837_sv2v_reg  <= w_data_i[141];
      \nz.mem_836_sv2v_reg  <= w_data_i[140];
      \nz.mem_835_sv2v_reg  <= w_data_i[139];
      \nz.mem_834_sv2v_reg  <= w_data_i[138];
      \nz.mem_833_sv2v_reg  <= w_data_i[137];
      \nz.mem_832_sv2v_reg  <= w_data_i[136];
      \nz.mem_831_sv2v_reg  <= w_data_i[135];
      \nz.mem_830_sv2v_reg  <= w_data_i[134];
      \nz.mem_829_sv2v_reg  <= w_data_i[133];
      \nz.mem_828_sv2v_reg  <= w_data_i[132];
      \nz.mem_827_sv2v_reg  <= w_data_i[131];
      \nz.mem_826_sv2v_reg  <= w_data_i[130];
      \nz.mem_825_sv2v_reg  <= w_data_i[129];
      \nz.mem_824_sv2v_reg  <= w_data_i[128];
      \nz.mem_823_sv2v_reg  <= w_data_i[127];
      \nz.mem_822_sv2v_reg  <= w_data_i[126];
      \nz.mem_821_sv2v_reg  <= w_data_i[125];
      \nz.mem_820_sv2v_reg  <= w_data_i[124];
      \nz.mem_819_sv2v_reg  <= w_data_i[123];
      \nz.mem_818_sv2v_reg  <= w_data_i[122];
      \nz.mem_817_sv2v_reg  <= w_data_i[121];
      \nz.mem_816_sv2v_reg  <= w_data_i[120];
      \nz.mem_815_sv2v_reg  <= w_data_i[119];
      \nz.mem_814_sv2v_reg  <= w_data_i[118];
      \nz.mem_813_sv2v_reg  <= w_data_i[117];
      \nz.mem_812_sv2v_reg  <= w_data_i[116];
      \nz.mem_811_sv2v_reg  <= w_data_i[115];
      \nz.mem_810_sv2v_reg  <= w_data_i[114];
      \nz.mem_809_sv2v_reg  <= w_data_i[113];
      \nz.mem_808_sv2v_reg  <= w_data_i[112];
      \nz.mem_807_sv2v_reg  <= w_data_i[111];
      \nz.mem_806_sv2v_reg  <= w_data_i[110];
      \nz.mem_805_sv2v_reg  <= w_data_i[109];
      \nz.mem_804_sv2v_reg  <= w_data_i[108];
      \nz.mem_803_sv2v_reg  <= w_data_i[107];
      \nz.mem_802_sv2v_reg  <= w_data_i[106];
      \nz.mem_801_sv2v_reg  <= w_data_i[105];
      \nz.mem_800_sv2v_reg  <= w_data_i[104];
      \nz.mem_799_sv2v_reg  <= w_data_i[103];
      \nz.mem_798_sv2v_reg  <= w_data_i[102];
      \nz.mem_797_sv2v_reg  <= w_data_i[101];
      \nz.mem_796_sv2v_reg  <= w_data_i[100];
      \nz.mem_795_sv2v_reg  <= w_data_i[99];
      \nz.mem_794_sv2v_reg  <= w_data_i[98];
      \nz.mem_793_sv2v_reg  <= w_data_i[97];
      \nz.mem_792_sv2v_reg  <= w_data_i[96];
      \nz.mem_791_sv2v_reg  <= w_data_i[95];
      \nz.mem_790_sv2v_reg  <= w_data_i[94];
      \nz.mem_789_sv2v_reg  <= w_data_i[93];
      \nz.mem_788_sv2v_reg  <= w_data_i[92];
      \nz.mem_787_sv2v_reg  <= w_data_i[91];
      \nz.mem_786_sv2v_reg  <= w_data_i[90];
      \nz.mem_785_sv2v_reg  <= w_data_i[89];
      \nz.mem_784_sv2v_reg  <= w_data_i[88];
      \nz.mem_783_sv2v_reg  <= w_data_i[87];
      \nz.mem_782_sv2v_reg  <= w_data_i[86];
      \nz.mem_781_sv2v_reg  <= w_data_i[85];
      \nz.mem_780_sv2v_reg  <= w_data_i[84];
      \nz.mem_779_sv2v_reg  <= w_data_i[83];
      \nz.mem_778_sv2v_reg  <= w_data_i[82];
      \nz.mem_777_sv2v_reg  <= w_data_i[81];
      \nz.mem_776_sv2v_reg  <= w_data_i[80];
      \nz.mem_775_sv2v_reg  <= w_data_i[79];
      \nz.mem_774_sv2v_reg  <= w_data_i[78];
      \nz.mem_773_sv2v_reg  <= w_data_i[77];
      \nz.mem_772_sv2v_reg  <= w_data_i[76];
      \nz.mem_771_sv2v_reg  <= w_data_i[75];
      \nz.mem_696_sv2v_reg  <= w_data_i[0];
    end 
    if(N43) begin
      \nz.mem_770_sv2v_reg  <= w_data_i[74];
      \nz.mem_769_sv2v_reg  <= w_data_i[73];
      \nz.mem_768_sv2v_reg  <= w_data_i[72];
      \nz.mem_767_sv2v_reg  <= w_data_i[71];
      \nz.mem_766_sv2v_reg  <= w_data_i[70];
      \nz.mem_765_sv2v_reg  <= w_data_i[69];
      \nz.mem_764_sv2v_reg  <= w_data_i[68];
      \nz.mem_763_sv2v_reg  <= w_data_i[67];
      \nz.mem_762_sv2v_reg  <= w_data_i[66];
      \nz.mem_761_sv2v_reg  <= w_data_i[65];
      \nz.mem_760_sv2v_reg  <= w_data_i[64];
      \nz.mem_759_sv2v_reg  <= w_data_i[63];
      \nz.mem_758_sv2v_reg  <= w_data_i[62];
      \nz.mem_757_sv2v_reg  <= w_data_i[61];
      \nz.mem_756_sv2v_reg  <= w_data_i[60];
      \nz.mem_755_sv2v_reg  <= w_data_i[59];
      \nz.mem_754_sv2v_reg  <= w_data_i[58];
      \nz.mem_753_sv2v_reg  <= w_data_i[57];
      \nz.mem_752_sv2v_reg  <= w_data_i[56];
      \nz.mem_751_sv2v_reg  <= w_data_i[55];
      \nz.mem_750_sv2v_reg  <= w_data_i[54];
      \nz.mem_749_sv2v_reg  <= w_data_i[53];
      \nz.mem_748_sv2v_reg  <= w_data_i[52];
      \nz.mem_747_sv2v_reg  <= w_data_i[51];
      \nz.mem_746_sv2v_reg  <= w_data_i[50];
      \nz.mem_745_sv2v_reg  <= w_data_i[49];
      \nz.mem_744_sv2v_reg  <= w_data_i[48];
      \nz.mem_743_sv2v_reg  <= w_data_i[47];
      \nz.mem_742_sv2v_reg  <= w_data_i[46];
      \nz.mem_741_sv2v_reg  <= w_data_i[45];
      \nz.mem_740_sv2v_reg  <= w_data_i[44];
      \nz.mem_739_sv2v_reg  <= w_data_i[43];
      \nz.mem_738_sv2v_reg  <= w_data_i[42];
      \nz.mem_737_sv2v_reg  <= w_data_i[41];
      \nz.mem_736_sv2v_reg  <= w_data_i[40];
      \nz.mem_735_sv2v_reg  <= w_data_i[39];
      \nz.mem_734_sv2v_reg  <= w_data_i[38];
      \nz.mem_733_sv2v_reg  <= w_data_i[37];
      \nz.mem_732_sv2v_reg  <= w_data_i[36];
      \nz.mem_731_sv2v_reg  <= w_data_i[35];
      \nz.mem_730_sv2v_reg  <= w_data_i[34];
      \nz.mem_729_sv2v_reg  <= w_data_i[33];
      \nz.mem_728_sv2v_reg  <= w_data_i[32];
      \nz.mem_727_sv2v_reg  <= w_data_i[31];
      \nz.mem_726_sv2v_reg  <= w_data_i[30];
      \nz.mem_725_sv2v_reg  <= w_data_i[29];
      \nz.mem_724_sv2v_reg  <= w_data_i[28];
      \nz.mem_723_sv2v_reg  <= w_data_i[27];
      \nz.mem_722_sv2v_reg  <= w_data_i[26];
      \nz.mem_721_sv2v_reg  <= w_data_i[25];
      \nz.mem_720_sv2v_reg  <= w_data_i[24];
      \nz.mem_719_sv2v_reg  <= w_data_i[23];
      \nz.mem_718_sv2v_reg  <= w_data_i[22];
      \nz.mem_717_sv2v_reg  <= w_data_i[21];
      \nz.mem_716_sv2v_reg  <= w_data_i[20];
      \nz.mem_715_sv2v_reg  <= w_data_i[19];
      \nz.mem_714_sv2v_reg  <= w_data_i[18];
      \nz.mem_713_sv2v_reg  <= w_data_i[17];
      \nz.mem_712_sv2v_reg  <= w_data_i[16];
      \nz.mem_711_sv2v_reg  <= w_data_i[15];
      \nz.mem_710_sv2v_reg  <= w_data_i[14];
      \nz.mem_709_sv2v_reg  <= w_data_i[13];
      \nz.mem_708_sv2v_reg  <= w_data_i[12];
      \nz.mem_707_sv2v_reg  <= w_data_i[11];
      \nz.mem_706_sv2v_reg  <= w_data_i[10];
      \nz.mem_705_sv2v_reg  <= w_data_i[9];
      \nz.mem_704_sv2v_reg  <= w_data_i[8];
      \nz.mem_703_sv2v_reg  <= w_data_i[7];
      \nz.mem_702_sv2v_reg  <= w_data_i[6];
      \nz.mem_701_sv2v_reg  <= w_data_i[5];
      \nz.mem_700_sv2v_reg  <= w_data_i[4];
      \nz.mem_699_sv2v_reg  <= w_data_i[3];
      \nz.mem_698_sv2v_reg  <= w_data_i[2];
      \nz.mem_697_sv2v_reg  <= w_data_i[1];
    end 
    if(N40) begin
      \nz.mem_695_sv2v_reg  <= w_data_i[173];
      \nz.mem_694_sv2v_reg  <= w_data_i[172];
      \nz.mem_693_sv2v_reg  <= w_data_i[171];
      \nz.mem_692_sv2v_reg  <= w_data_i[170];
      \nz.mem_691_sv2v_reg  <= w_data_i[169];
      \nz.mem_690_sv2v_reg  <= w_data_i[168];
      \nz.mem_689_sv2v_reg  <= w_data_i[167];
      \nz.mem_688_sv2v_reg  <= w_data_i[166];
      \nz.mem_687_sv2v_reg  <= w_data_i[165];
      \nz.mem_686_sv2v_reg  <= w_data_i[164];
      \nz.mem_685_sv2v_reg  <= w_data_i[163];
      \nz.mem_684_sv2v_reg  <= w_data_i[162];
      \nz.mem_683_sv2v_reg  <= w_data_i[161];
      \nz.mem_682_sv2v_reg  <= w_data_i[160];
      \nz.mem_681_sv2v_reg  <= w_data_i[159];
      \nz.mem_680_sv2v_reg  <= w_data_i[158];
      \nz.mem_679_sv2v_reg  <= w_data_i[157];
      \nz.mem_678_sv2v_reg  <= w_data_i[156];
      \nz.mem_677_sv2v_reg  <= w_data_i[155];
      \nz.mem_676_sv2v_reg  <= w_data_i[154];
      \nz.mem_675_sv2v_reg  <= w_data_i[153];
      \nz.mem_674_sv2v_reg  <= w_data_i[152];
      \nz.mem_673_sv2v_reg  <= w_data_i[151];
      \nz.mem_672_sv2v_reg  <= w_data_i[150];
      \nz.mem_671_sv2v_reg  <= w_data_i[149];
      \nz.mem_670_sv2v_reg  <= w_data_i[148];
      \nz.mem_669_sv2v_reg  <= w_data_i[147];
      \nz.mem_668_sv2v_reg  <= w_data_i[146];
      \nz.mem_667_sv2v_reg  <= w_data_i[145];
      \nz.mem_666_sv2v_reg  <= w_data_i[144];
      \nz.mem_665_sv2v_reg  <= w_data_i[143];
      \nz.mem_664_sv2v_reg  <= w_data_i[142];
      \nz.mem_663_sv2v_reg  <= w_data_i[141];
      \nz.mem_662_sv2v_reg  <= w_data_i[140];
      \nz.mem_661_sv2v_reg  <= w_data_i[139];
      \nz.mem_660_sv2v_reg  <= w_data_i[138];
      \nz.mem_659_sv2v_reg  <= w_data_i[137];
      \nz.mem_658_sv2v_reg  <= w_data_i[136];
      \nz.mem_657_sv2v_reg  <= w_data_i[135];
      \nz.mem_656_sv2v_reg  <= w_data_i[134];
      \nz.mem_655_sv2v_reg  <= w_data_i[133];
      \nz.mem_654_sv2v_reg  <= w_data_i[132];
      \nz.mem_653_sv2v_reg  <= w_data_i[131];
      \nz.mem_652_sv2v_reg  <= w_data_i[130];
      \nz.mem_651_sv2v_reg  <= w_data_i[129];
      \nz.mem_650_sv2v_reg  <= w_data_i[128];
      \nz.mem_649_sv2v_reg  <= w_data_i[127];
      \nz.mem_648_sv2v_reg  <= w_data_i[126];
      \nz.mem_647_sv2v_reg  <= w_data_i[125];
      \nz.mem_646_sv2v_reg  <= w_data_i[124];
      \nz.mem_645_sv2v_reg  <= w_data_i[123];
      \nz.mem_644_sv2v_reg  <= w_data_i[122];
      \nz.mem_643_sv2v_reg  <= w_data_i[121];
      \nz.mem_642_sv2v_reg  <= w_data_i[120];
      \nz.mem_641_sv2v_reg  <= w_data_i[119];
      \nz.mem_640_sv2v_reg  <= w_data_i[118];
      \nz.mem_639_sv2v_reg  <= w_data_i[117];
      \nz.mem_638_sv2v_reg  <= w_data_i[116];
      \nz.mem_637_sv2v_reg  <= w_data_i[115];
      \nz.mem_636_sv2v_reg  <= w_data_i[114];
      \nz.mem_635_sv2v_reg  <= w_data_i[113];
      \nz.mem_634_sv2v_reg  <= w_data_i[112];
      \nz.mem_633_sv2v_reg  <= w_data_i[111];
      \nz.mem_632_sv2v_reg  <= w_data_i[110];
      \nz.mem_631_sv2v_reg  <= w_data_i[109];
      \nz.mem_630_sv2v_reg  <= w_data_i[108];
      \nz.mem_629_sv2v_reg  <= w_data_i[107];
      \nz.mem_628_sv2v_reg  <= w_data_i[106];
      \nz.mem_627_sv2v_reg  <= w_data_i[105];
      \nz.mem_626_sv2v_reg  <= w_data_i[104];
      \nz.mem_625_sv2v_reg  <= w_data_i[103];
      \nz.mem_624_sv2v_reg  <= w_data_i[102];
      \nz.mem_623_sv2v_reg  <= w_data_i[101];
      \nz.mem_622_sv2v_reg  <= w_data_i[100];
      \nz.mem_621_sv2v_reg  <= w_data_i[99];
      \nz.mem_620_sv2v_reg  <= w_data_i[98];
      \nz.mem_619_sv2v_reg  <= w_data_i[97];
      \nz.mem_618_sv2v_reg  <= w_data_i[96];
      \nz.mem_617_sv2v_reg  <= w_data_i[95];
      \nz.mem_616_sv2v_reg  <= w_data_i[94];
      \nz.mem_615_sv2v_reg  <= w_data_i[93];
      \nz.mem_614_sv2v_reg  <= w_data_i[92];
      \nz.mem_613_sv2v_reg  <= w_data_i[91];
      \nz.mem_612_sv2v_reg  <= w_data_i[90];
      \nz.mem_611_sv2v_reg  <= w_data_i[89];
      \nz.mem_610_sv2v_reg  <= w_data_i[88];
      \nz.mem_609_sv2v_reg  <= w_data_i[87];
      \nz.mem_608_sv2v_reg  <= w_data_i[86];
      \nz.mem_607_sv2v_reg  <= w_data_i[85];
      \nz.mem_606_sv2v_reg  <= w_data_i[84];
      \nz.mem_605_sv2v_reg  <= w_data_i[83];
      \nz.mem_604_sv2v_reg  <= w_data_i[82];
      \nz.mem_603_sv2v_reg  <= w_data_i[81];
      \nz.mem_602_sv2v_reg  <= w_data_i[80];
      \nz.mem_601_sv2v_reg  <= w_data_i[79];
      \nz.mem_600_sv2v_reg  <= w_data_i[78];
      \nz.mem_599_sv2v_reg  <= w_data_i[77];
      \nz.mem_598_sv2v_reg  <= w_data_i[76];
      \nz.mem_597_sv2v_reg  <= w_data_i[75];
      \nz.mem_522_sv2v_reg  <= w_data_i[0];
    end 
    if(N41) begin
      \nz.mem_596_sv2v_reg  <= w_data_i[74];
      \nz.mem_595_sv2v_reg  <= w_data_i[73];
      \nz.mem_594_sv2v_reg  <= w_data_i[72];
      \nz.mem_593_sv2v_reg  <= w_data_i[71];
      \nz.mem_592_sv2v_reg  <= w_data_i[70];
      \nz.mem_591_sv2v_reg  <= w_data_i[69];
      \nz.mem_590_sv2v_reg  <= w_data_i[68];
      \nz.mem_589_sv2v_reg  <= w_data_i[67];
      \nz.mem_588_sv2v_reg  <= w_data_i[66];
      \nz.mem_587_sv2v_reg  <= w_data_i[65];
      \nz.mem_586_sv2v_reg  <= w_data_i[64];
      \nz.mem_585_sv2v_reg  <= w_data_i[63];
      \nz.mem_584_sv2v_reg  <= w_data_i[62];
      \nz.mem_583_sv2v_reg  <= w_data_i[61];
      \nz.mem_582_sv2v_reg  <= w_data_i[60];
      \nz.mem_581_sv2v_reg  <= w_data_i[59];
      \nz.mem_580_sv2v_reg  <= w_data_i[58];
      \nz.mem_579_sv2v_reg  <= w_data_i[57];
      \nz.mem_578_sv2v_reg  <= w_data_i[56];
      \nz.mem_577_sv2v_reg  <= w_data_i[55];
      \nz.mem_576_sv2v_reg  <= w_data_i[54];
      \nz.mem_575_sv2v_reg  <= w_data_i[53];
      \nz.mem_574_sv2v_reg  <= w_data_i[52];
      \nz.mem_573_sv2v_reg  <= w_data_i[51];
      \nz.mem_572_sv2v_reg  <= w_data_i[50];
      \nz.mem_571_sv2v_reg  <= w_data_i[49];
      \nz.mem_570_sv2v_reg  <= w_data_i[48];
      \nz.mem_569_sv2v_reg  <= w_data_i[47];
      \nz.mem_568_sv2v_reg  <= w_data_i[46];
      \nz.mem_567_sv2v_reg  <= w_data_i[45];
      \nz.mem_566_sv2v_reg  <= w_data_i[44];
      \nz.mem_565_sv2v_reg  <= w_data_i[43];
      \nz.mem_564_sv2v_reg  <= w_data_i[42];
      \nz.mem_563_sv2v_reg  <= w_data_i[41];
      \nz.mem_562_sv2v_reg  <= w_data_i[40];
      \nz.mem_561_sv2v_reg  <= w_data_i[39];
      \nz.mem_560_sv2v_reg  <= w_data_i[38];
      \nz.mem_559_sv2v_reg  <= w_data_i[37];
      \nz.mem_558_sv2v_reg  <= w_data_i[36];
      \nz.mem_557_sv2v_reg  <= w_data_i[35];
      \nz.mem_556_sv2v_reg  <= w_data_i[34];
      \nz.mem_555_sv2v_reg  <= w_data_i[33];
      \nz.mem_554_sv2v_reg  <= w_data_i[32];
      \nz.mem_553_sv2v_reg  <= w_data_i[31];
      \nz.mem_552_sv2v_reg  <= w_data_i[30];
      \nz.mem_551_sv2v_reg  <= w_data_i[29];
      \nz.mem_550_sv2v_reg  <= w_data_i[28];
      \nz.mem_549_sv2v_reg  <= w_data_i[27];
      \nz.mem_548_sv2v_reg  <= w_data_i[26];
      \nz.mem_547_sv2v_reg  <= w_data_i[25];
      \nz.mem_546_sv2v_reg  <= w_data_i[24];
      \nz.mem_545_sv2v_reg  <= w_data_i[23];
      \nz.mem_544_sv2v_reg  <= w_data_i[22];
      \nz.mem_543_sv2v_reg  <= w_data_i[21];
      \nz.mem_542_sv2v_reg  <= w_data_i[20];
      \nz.mem_541_sv2v_reg  <= w_data_i[19];
      \nz.mem_540_sv2v_reg  <= w_data_i[18];
      \nz.mem_539_sv2v_reg  <= w_data_i[17];
      \nz.mem_538_sv2v_reg  <= w_data_i[16];
      \nz.mem_537_sv2v_reg  <= w_data_i[15];
      \nz.mem_536_sv2v_reg  <= w_data_i[14];
      \nz.mem_535_sv2v_reg  <= w_data_i[13];
      \nz.mem_534_sv2v_reg  <= w_data_i[12];
      \nz.mem_533_sv2v_reg  <= w_data_i[11];
      \nz.mem_532_sv2v_reg  <= w_data_i[10];
      \nz.mem_531_sv2v_reg  <= w_data_i[9];
      \nz.mem_530_sv2v_reg  <= w_data_i[8];
      \nz.mem_529_sv2v_reg  <= w_data_i[7];
      \nz.mem_528_sv2v_reg  <= w_data_i[6];
      \nz.mem_527_sv2v_reg  <= w_data_i[5];
      \nz.mem_526_sv2v_reg  <= w_data_i[4];
      \nz.mem_525_sv2v_reg  <= w_data_i[3];
      \nz.mem_524_sv2v_reg  <= w_data_i[2];
      \nz.mem_523_sv2v_reg  <= w_data_i[1];
    end 
    if(N38) begin
      \nz.mem_521_sv2v_reg  <= w_data_i[173];
      \nz.mem_520_sv2v_reg  <= w_data_i[172];
      \nz.mem_519_sv2v_reg  <= w_data_i[171];
      \nz.mem_518_sv2v_reg  <= w_data_i[170];
      \nz.mem_517_sv2v_reg  <= w_data_i[169];
      \nz.mem_516_sv2v_reg  <= w_data_i[168];
      \nz.mem_515_sv2v_reg  <= w_data_i[167];
      \nz.mem_514_sv2v_reg  <= w_data_i[166];
      \nz.mem_513_sv2v_reg  <= w_data_i[165];
      \nz.mem_512_sv2v_reg  <= w_data_i[164];
      \nz.mem_511_sv2v_reg  <= w_data_i[163];
      \nz.mem_510_sv2v_reg  <= w_data_i[162];
      \nz.mem_509_sv2v_reg  <= w_data_i[161];
      \nz.mem_508_sv2v_reg  <= w_data_i[160];
      \nz.mem_507_sv2v_reg  <= w_data_i[159];
      \nz.mem_506_sv2v_reg  <= w_data_i[158];
      \nz.mem_505_sv2v_reg  <= w_data_i[157];
      \nz.mem_504_sv2v_reg  <= w_data_i[156];
      \nz.mem_503_sv2v_reg  <= w_data_i[155];
      \nz.mem_502_sv2v_reg  <= w_data_i[154];
      \nz.mem_501_sv2v_reg  <= w_data_i[153];
      \nz.mem_500_sv2v_reg  <= w_data_i[152];
      \nz.mem_499_sv2v_reg  <= w_data_i[151];
      \nz.mem_498_sv2v_reg  <= w_data_i[150];
      \nz.mem_497_sv2v_reg  <= w_data_i[149];
      \nz.mem_496_sv2v_reg  <= w_data_i[148];
      \nz.mem_495_sv2v_reg  <= w_data_i[147];
      \nz.mem_494_sv2v_reg  <= w_data_i[146];
      \nz.mem_493_sv2v_reg  <= w_data_i[145];
      \nz.mem_492_sv2v_reg  <= w_data_i[144];
      \nz.mem_491_sv2v_reg  <= w_data_i[143];
      \nz.mem_490_sv2v_reg  <= w_data_i[142];
      \nz.mem_489_sv2v_reg  <= w_data_i[141];
      \nz.mem_488_sv2v_reg  <= w_data_i[140];
      \nz.mem_487_sv2v_reg  <= w_data_i[139];
      \nz.mem_486_sv2v_reg  <= w_data_i[138];
      \nz.mem_485_sv2v_reg  <= w_data_i[137];
      \nz.mem_484_sv2v_reg  <= w_data_i[136];
      \nz.mem_483_sv2v_reg  <= w_data_i[135];
      \nz.mem_482_sv2v_reg  <= w_data_i[134];
      \nz.mem_481_sv2v_reg  <= w_data_i[133];
      \nz.mem_480_sv2v_reg  <= w_data_i[132];
      \nz.mem_479_sv2v_reg  <= w_data_i[131];
      \nz.mem_478_sv2v_reg  <= w_data_i[130];
      \nz.mem_477_sv2v_reg  <= w_data_i[129];
      \nz.mem_476_sv2v_reg  <= w_data_i[128];
      \nz.mem_475_sv2v_reg  <= w_data_i[127];
      \nz.mem_474_sv2v_reg  <= w_data_i[126];
      \nz.mem_473_sv2v_reg  <= w_data_i[125];
      \nz.mem_472_sv2v_reg  <= w_data_i[124];
      \nz.mem_471_sv2v_reg  <= w_data_i[123];
      \nz.mem_470_sv2v_reg  <= w_data_i[122];
      \nz.mem_469_sv2v_reg  <= w_data_i[121];
      \nz.mem_468_sv2v_reg  <= w_data_i[120];
      \nz.mem_467_sv2v_reg  <= w_data_i[119];
      \nz.mem_466_sv2v_reg  <= w_data_i[118];
      \nz.mem_465_sv2v_reg  <= w_data_i[117];
      \nz.mem_464_sv2v_reg  <= w_data_i[116];
      \nz.mem_463_sv2v_reg  <= w_data_i[115];
      \nz.mem_462_sv2v_reg  <= w_data_i[114];
      \nz.mem_461_sv2v_reg  <= w_data_i[113];
      \nz.mem_460_sv2v_reg  <= w_data_i[112];
      \nz.mem_459_sv2v_reg  <= w_data_i[111];
      \nz.mem_458_sv2v_reg  <= w_data_i[110];
      \nz.mem_457_sv2v_reg  <= w_data_i[109];
      \nz.mem_456_sv2v_reg  <= w_data_i[108];
      \nz.mem_455_sv2v_reg  <= w_data_i[107];
      \nz.mem_454_sv2v_reg  <= w_data_i[106];
      \nz.mem_453_sv2v_reg  <= w_data_i[105];
      \nz.mem_452_sv2v_reg  <= w_data_i[104];
      \nz.mem_451_sv2v_reg  <= w_data_i[103];
      \nz.mem_450_sv2v_reg  <= w_data_i[102];
      \nz.mem_449_sv2v_reg  <= w_data_i[101];
      \nz.mem_448_sv2v_reg  <= w_data_i[100];
      \nz.mem_447_sv2v_reg  <= w_data_i[99];
      \nz.mem_446_sv2v_reg  <= w_data_i[98];
      \nz.mem_445_sv2v_reg  <= w_data_i[97];
      \nz.mem_444_sv2v_reg  <= w_data_i[96];
      \nz.mem_443_sv2v_reg  <= w_data_i[95];
      \nz.mem_442_sv2v_reg  <= w_data_i[94];
      \nz.mem_441_sv2v_reg  <= w_data_i[93];
      \nz.mem_440_sv2v_reg  <= w_data_i[92];
      \nz.mem_439_sv2v_reg  <= w_data_i[91];
      \nz.mem_438_sv2v_reg  <= w_data_i[90];
      \nz.mem_437_sv2v_reg  <= w_data_i[89];
      \nz.mem_436_sv2v_reg  <= w_data_i[88];
      \nz.mem_435_sv2v_reg  <= w_data_i[87];
      \nz.mem_434_sv2v_reg  <= w_data_i[86];
      \nz.mem_433_sv2v_reg  <= w_data_i[85];
      \nz.mem_432_sv2v_reg  <= w_data_i[84];
      \nz.mem_431_sv2v_reg  <= w_data_i[83];
      \nz.mem_430_sv2v_reg  <= w_data_i[82];
      \nz.mem_429_sv2v_reg  <= w_data_i[81];
      \nz.mem_428_sv2v_reg  <= w_data_i[80];
      \nz.mem_427_sv2v_reg  <= w_data_i[79];
      \nz.mem_426_sv2v_reg  <= w_data_i[78];
      \nz.mem_425_sv2v_reg  <= w_data_i[77];
      \nz.mem_424_sv2v_reg  <= w_data_i[76];
      \nz.mem_423_sv2v_reg  <= w_data_i[75];
      \nz.mem_348_sv2v_reg  <= w_data_i[0];
    end 
    if(N39) begin
      \nz.mem_422_sv2v_reg  <= w_data_i[74];
      \nz.mem_421_sv2v_reg  <= w_data_i[73];
      \nz.mem_420_sv2v_reg  <= w_data_i[72];
      \nz.mem_419_sv2v_reg  <= w_data_i[71];
      \nz.mem_418_sv2v_reg  <= w_data_i[70];
      \nz.mem_417_sv2v_reg  <= w_data_i[69];
      \nz.mem_416_sv2v_reg  <= w_data_i[68];
      \nz.mem_415_sv2v_reg  <= w_data_i[67];
      \nz.mem_414_sv2v_reg  <= w_data_i[66];
      \nz.mem_413_sv2v_reg  <= w_data_i[65];
      \nz.mem_412_sv2v_reg  <= w_data_i[64];
      \nz.mem_411_sv2v_reg  <= w_data_i[63];
      \nz.mem_410_sv2v_reg  <= w_data_i[62];
      \nz.mem_409_sv2v_reg  <= w_data_i[61];
      \nz.mem_408_sv2v_reg  <= w_data_i[60];
      \nz.mem_407_sv2v_reg  <= w_data_i[59];
      \nz.mem_406_sv2v_reg  <= w_data_i[58];
      \nz.mem_405_sv2v_reg  <= w_data_i[57];
      \nz.mem_404_sv2v_reg  <= w_data_i[56];
      \nz.mem_403_sv2v_reg  <= w_data_i[55];
      \nz.mem_402_sv2v_reg  <= w_data_i[54];
      \nz.mem_401_sv2v_reg  <= w_data_i[53];
      \nz.mem_400_sv2v_reg  <= w_data_i[52];
      \nz.mem_399_sv2v_reg  <= w_data_i[51];
      \nz.mem_398_sv2v_reg  <= w_data_i[50];
      \nz.mem_397_sv2v_reg  <= w_data_i[49];
      \nz.mem_396_sv2v_reg  <= w_data_i[48];
      \nz.mem_395_sv2v_reg  <= w_data_i[47];
      \nz.mem_394_sv2v_reg  <= w_data_i[46];
      \nz.mem_393_sv2v_reg  <= w_data_i[45];
      \nz.mem_392_sv2v_reg  <= w_data_i[44];
      \nz.mem_391_sv2v_reg  <= w_data_i[43];
      \nz.mem_390_sv2v_reg  <= w_data_i[42];
      \nz.mem_389_sv2v_reg  <= w_data_i[41];
      \nz.mem_388_sv2v_reg  <= w_data_i[40];
      \nz.mem_387_sv2v_reg  <= w_data_i[39];
      \nz.mem_386_sv2v_reg  <= w_data_i[38];
      \nz.mem_385_sv2v_reg  <= w_data_i[37];
      \nz.mem_384_sv2v_reg  <= w_data_i[36];
      \nz.mem_383_sv2v_reg  <= w_data_i[35];
      \nz.mem_382_sv2v_reg  <= w_data_i[34];
      \nz.mem_381_sv2v_reg  <= w_data_i[33];
      \nz.mem_380_sv2v_reg  <= w_data_i[32];
      \nz.mem_379_sv2v_reg  <= w_data_i[31];
      \nz.mem_378_sv2v_reg  <= w_data_i[30];
      \nz.mem_377_sv2v_reg  <= w_data_i[29];
      \nz.mem_376_sv2v_reg  <= w_data_i[28];
      \nz.mem_375_sv2v_reg  <= w_data_i[27];
      \nz.mem_374_sv2v_reg  <= w_data_i[26];
      \nz.mem_373_sv2v_reg  <= w_data_i[25];
      \nz.mem_372_sv2v_reg  <= w_data_i[24];
      \nz.mem_371_sv2v_reg  <= w_data_i[23];
      \nz.mem_370_sv2v_reg  <= w_data_i[22];
      \nz.mem_369_sv2v_reg  <= w_data_i[21];
      \nz.mem_368_sv2v_reg  <= w_data_i[20];
      \nz.mem_367_sv2v_reg  <= w_data_i[19];
      \nz.mem_366_sv2v_reg  <= w_data_i[18];
      \nz.mem_365_sv2v_reg  <= w_data_i[17];
      \nz.mem_364_sv2v_reg  <= w_data_i[16];
      \nz.mem_363_sv2v_reg  <= w_data_i[15];
      \nz.mem_362_sv2v_reg  <= w_data_i[14];
      \nz.mem_361_sv2v_reg  <= w_data_i[13];
      \nz.mem_360_sv2v_reg  <= w_data_i[12];
      \nz.mem_359_sv2v_reg  <= w_data_i[11];
      \nz.mem_358_sv2v_reg  <= w_data_i[10];
      \nz.mem_357_sv2v_reg  <= w_data_i[9];
      \nz.mem_356_sv2v_reg  <= w_data_i[8];
      \nz.mem_355_sv2v_reg  <= w_data_i[7];
      \nz.mem_354_sv2v_reg  <= w_data_i[6];
      \nz.mem_353_sv2v_reg  <= w_data_i[5];
      \nz.mem_352_sv2v_reg  <= w_data_i[4];
      \nz.mem_351_sv2v_reg  <= w_data_i[3];
      \nz.mem_350_sv2v_reg  <= w_data_i[2];
      \nz.mem_349_sv2v_reg  <= w_data_i[1];
    end 
    if(N36) begin
      \nz.mem_347_sv2v_reg  <= w_data_i[173];
      \nz.mem_346_sv2v_reg  <= w_data_i[172];
      \nz.mem_345_sv2v_reg  <= w_data_i[171];
      \nz.mem_344_sv2v_reg  <= w_data_i[170];
      \nz.mem_343_sv2v_reg  <= w_data_i[169];
      \nz.mem_342_sv2v_reg  <= w_data_i[168];
      \nz.mem_341_sv2v_reg  <= w_data_i[167];
      \nz.mem_340_sv2v_reg  <= w_data_i[166];
      \nz.mem_339_sv2v_reg  <= w_data_i[165];
      \nz.mem_338_sv2v_reg  <= w_data_i[164];
      \nz.mem_337_sv2v_reg  <= w_data_i[163];
      \nz.mem_336_sv2v_reg  <= w_data_i[162];
      \nz.mem_335_sv2v_reg  <= w_data_i[161];
      \nz.mem_334_sv2v_reg  <= w_data_i[160];
      \nz.mem_333_sv2v_reg  <= w_data_i[159];
      \nz.mem_332_sv2v_reg  <= w_data_i[158];
      \nz.mem_331_sv2v_reg  <= w_data_i[157];
      \nz.mem_330_sv2v_reg  <= w_data_i[156];
      \nz.mem_329_sv2v_reg  <= w_data_i[155];
      \nz.mem_328_sv2v_reg  <= w_data_i[154];
      \nz.mem_327_sv2v_reg  <= w_data_i[153];
      \nz.mem_326_sv2v_reg  <= w_data_i[152];
      \nz.mem_325_sv2v_reg  <= w_data_i[151];
      \nz.mem_324_sv2v_reg  <= w_data_i[150];
      \nz.mem_323_sv2v_reg  <= w_data_i[149];
      \nz.mem_322_sv2v_reg  <= w_data_i[148];
      \nz.mem_321_sv2v_reg  <= w_data_i[147];
      \nz.mem_320_sv2v_reg  <= w_data_i[146];
      \nz.mem_319_sv2v_reg  <= w_data_i[145];
      \nz.mem_318_sv2v_reg  <= w_data_i[144];
      \nz.mem_317_sv2v_reg  <= w_data_i[143];
      \nz.mem_316_sv2v_reg  <= w_data_i[142];
      \nz.mem_315_sv2v_reg  <= w_data_i[141];
      \nz.mem_314_sv2v_reg  <= w_data_i[140];
      \nz.mem_313_sv2v_reg  <= w_data_i[139];
      \nz.mem_312_sv2v_reg  <= w_data_i[138];
      \nz.mem_311_sv2v_reg  <= w_data_i[137];
      \nz.mem_310_sv2v_reg  <= w_data_i[136];
      \nz.mem_309_sv2v_reg  <= w_data_i[135];
      \nz.mem_308_sv2v_reg  <= w_data_i[134];
      \nz.mem_307_sv2v_reg  <= w_data_i[133];
      \nz.mem_306_sv2v_reg  <= w_data_i[132];
      \nz.mem_305_sv2v_reg  <= w_data_i[131];
      \nz.mem_304_sv2v_reg  <= w_data_i[130];
      \nz.mem_303_sv2v_reg  <= w_data_i[129];
      \nz.mem_302_sv2v_reg  <= w_data_i[128];
      \nz.mem_301_sv2v_reg  <= w_data_i[127];
      \nz.mem_300_sv2v_reg  <= w_data_i[126];
      \nz.mem_299_sv2v_reg  <= w_data_i[125];
      \nz.mem_298_sv2v_reg  <= w_data_i[124];
      \nz.mem_297_sv2v_reg  <= w_data_i[123];
      \nz.mem_296_sv2v_reg  <= w_data_i[122];
      \nz.mem_295_sv2v_reg  <= w_data_i[121];
      \nz.mem_294_sv2v_reg  <= w_data_i[120];
      \nz.mem_293_sv2v_reg  <= w_data_i[119];
      \nz.mem_292_sv2v_reg  <= w_data_i[118];
      \nz.mem_291_sv2v_reg  <= w_data_i[117];
      \nz.mem_290_sv2v_reg  <= w_data_i[116];
      \nz.mem_289_sv2v_reg  <= w_data_i[115];
      \nz.mem_288_sv2v_reg  <= w_data_i[114];
      \nz.mem_287_sv2v_reg  <= w_data_i[113];
      \nz.mem_286_sv2v_reg  <= w_data_i[112];
      \nz.mem_285_sv2v_reg  <= w_data_i[111];
      \nz.mem_284_sv2v_reg  <= w_data_i[110];
      \nz.mem_283_sv2v_reg  <= w_data_i[109];
      \nz.mem_282_sv2v_reg  <= w_data_i[108];
      \nz.mem_281_sv2v_reg  <= w_data_i[107];
      \nz.mem_280_sv2v_reg  <= w_data_i[106];
      \nz.mem_279_sv2v_reg  <= w_data_i[105];
      \nz.mem_278_sv2v_reg  <= w_data_i[104];
      \nz.mem_277_sv2v_reg  <= w_data_i[103];
      \nz.mem_276_sv2v_reg  <= w_data_i[102];
      \nz.mem_275_sv2v_reg  <= w_data_i[101];
      \nz.mem_274_sv2v_reg  <= w_data_i[100];
      \nz.mem_273_sv2v_reg  <= w_data_i[99];
      \nz.mem_272_sv2v_reg  <= w_data_i[98];
      \nz.mem_271_sv2v_reg  <= w_data_i[97];
      \nz.mem_270_sv2v_reg  <= w_data_i[96];
      \nz.mem_269_sv2v_reg  <= w_data_i[95];
      \nz.mem_268_sv2v_reg  <= w_data_i[94];
      \nz.mem_267_sv2v_reg  <= w_data_i[93];
      \nz.mem_266_sv2v_reg  <= w_data_i[92];
      \nz.mem_265_sv2v_reg  <= w_data_i[91];
      \nz.mem_264_sv2v_reg  <= w_data_i[90];
      \nz.mem_263_sv2v_reg  <= w_data_i[89];
      \nz.mem_262_sv2v_reg  <= w_data_i[88];
      \nz.mem_261_sv2v_reg  <= w_data_i[87];
      \nz.mem_260_sv2v_reg  <= w_data_i[86];
      \nz.mem_259_sv2v_reg  <= w_data_i[85];
      \nz.mem_258_sv2v_reg  <= w_data_i[84];
      \nz.mem_257_sv2v_reg  <= w_data_i[83];
      \nz.mem_256_sv2v_reg  <= w_data_i[82];
      \nz.mem_255_sv2v_reg  <= w_data_i[81];
      \nz.mem_254_sv2v_reg  <= w_data_i[80];
      \nz.mem_253_sv2v_reg  <= w_data_i[79];
      \nz.mem_252_sv2v_reg  <= w_data_i[78];
      \nz.mem_251_sv2v_reg  <= w_data_i[77];
      \nz.mem_250_sv2v_reg  <= w_data_i[76];
      \nz.mem_249_sv2v_reg  <= w_data_i[75];
      \nz.mem_174_sv2v_reg  <= w_data_i[0];
    end 
    if(N37) begin
      \nz.mem_248_sv2v_reg  <= w_data_i[74];
      \nz.mem_247_sv2v_reg  <= w_data_i[73];
      \nz.mem_246_sv2v_reg  <= w_data_i[72];
      \nz.mem_245_sv2v_reg  <= w_data_i[71];
      \nz.mem_244_sv2v_reg  <= w_data_i[70];
      \nz.mem_243_sv2v_reg  <= w_data_i[69];
      \nz.mem_242_sv2v_reg  <= w_data_i[68];
      \nz.mem_241_sv2v_reg  <= w_data_i[67];
      \nz.mem_240_sv2v_reg  <= w_data_i[66];
      \nz.mem_239_sv2v_reg  <= w_data_i[65];
      \nz.mem_238_sv2v_reg  <= w_data_i[64];
      \nz.mem_237_sv2v_reg  <= w_data_i[63];
      \nz.mem_236_sv2v_reg  <= w_data_i[62];
      \nz.mem_235_sv2v_reg  <= w_data_i[61];
      \nz.mem_234_sv2v_reg  <= w_data_i[60];
      \nz.mem_233_sv2v_reg  <= w_data_i[59];
      \nz.mem_232_sv2v_reg  <= w_data_i[58];
      \nz.mem_231_sv2v_reg  <= w_data_i[57];
      \nz.mem_230_sv2v_reg  <= w_data_i[56];
      \nz.mem_229_sv2v_reg  <= w_data_i[55];
      \nz.mem_228_sv2v_reg  <= w_data_i[54];
      \nz.mem_227_sv2v_reg  <= w_data_i[53];
      \nz.mem_226_sv2v_reg  <= w_data_i[52];
      \nz.mem_225_sv2v_reg  <= w_data_i[51];
      \nz.mem_224_sv2v_reg  <= w_data_i[50];
      \nz.mem_223_sv2v_reg  <= w_data_i[49];
      \nz.mem_222_sv2v_reg  <= w_data_i[48];
      \nz.mem_221_sv2v_reg  <= w_data_i[47];
      \nz.mem_220_sv2v_reg  <= w_data_i[46];
      \nz.mem_219_sv2v_reg  <= w_data_i[45];
      \nz.mem_218_sv2v_reg  <= w_data_i[44];
      \nz.mem_217_sv2v_reg  <= w_data_i[43];
      \nz.mem_216_sv2v_reg  <= w_data_i[42];
      \nz.mem_215_sv2v_reg  <= w_data_i[41];
      \nz.mem_214_sv2v_reg  <= w_data_i[40];
      \nz.mem_213_sv2v_reg  <= w_data_i[39];
      \nz.mem_212_sv2v_reg  <= w_data_i[38];
      \nz.mem_211_sv2v_reg  <= w_data_i[37];
      \nz.mem_210_sv2v_reg  <= w_data_i[36];
      \nz.mem_209_sv2v_reg  <= w_data_i[35];
      \nz.mem_208_sv2v_reg  <= w_data_i[34];
      \nz.mem_207_sv2v_reg  <= w_data_i[33];
      \nz.mem_206_sv2v_reg  <= w_data_i[32];
      \nz.mem_205_sv2v_reg  <= w_data_i[31];
      \nz.mem_204_sv2v_reg  <= w_data_i[30];
      \nz.mem_203_sv2v_reg  <= w_data_i[29];
      \nz.mem_202_sv2v_reg  <= w_data_i[28];
      \nz.mem_201_sv2v_reg  <= w_data_i[27];
      \nz.mem_200_sv2v_reg  <= w_data_i[26];
      \nz.mem_199_sv2v_reg  <= w_data_i[25];
      \nz.mem_198_sv2v_reg  <= w_data_i[24];
      \nz.mem_197_sv2v_reg  <= w_data_i[23];
      \nz.mem_196_sv2v_reg  <= w_data_i[22];
      \nz.mem_195_sv2v_reg  <= w_data_i[21];
      \nz.mem_194_sv2v_reg  <= w_data_i[20];
      \nz.mem_193_sv2v_reg  <= w_data_i[19];
      \nz.mem_192_sv2v_reg  <= w_data_i[18];
      \nz.mem_191_sv2v_reg  <= w_data_i[17];
      \nz.mem_190_sv2v_reg  <= w_data_i[16];
      \nz.mem_189_sv2v_reg  <= w_data_i[15];
      \nz.mem_188_sv2v_reg  <= w_data_i[14];
      \nz.mem_187_sv2v_reg  <= w_data_i[13];
      \nz.mem_186_sv2v_reg  <= w_data_i[12];
      \nz.mem_185_sv2v_reg  <= w_data_i[11];
      \nz.mem_184_sv2v_reg  <= w_data_i[10];
      \nz.mem_183_sv2v_reg  <= w_data_i[9];
      \nz.mem_182_sv2v_reg  <= w_data_i[8];
      \nz.mem_181_sv2v_reg  <= w_data_i[7];
      \nz.mem_180_sv2v_reg  <= w_data_i[6];
      \nz.mem_179_sv2v_reg  <= w_data_i[5];
      \nz.mem_178_sv2v_reg  <= w_data_i[4];
      \nz.mem_177_sv2v_reg  <= w_data_i[3];
      \nz.mem_176_sv2v_reg  <= w_data_i[2];
      \nz.mem_175_sv2v_reg  <= w_data_i[1];
    end 
    if(N34) begin
      \nz.mem_173_sv2v_reg  <= w_data_i[173];
      \nz.mem_172_sv2v_reg  <= w_data_i[172];
      \nz.mem_171_sv2v_reg  <= w_data_i[171];
      \nz.mem_170_sv2v_reg  <= w_data_i[170];
      \nz.mem_169_sv2v_reg  <= w_data_i[169];
      \nz.mem_168_sv2v_reg  <= w_data_i[168];
      \nz.mem_167_sv2v_reg  <= w_data_i[167];
      \nz.mem_166_sv2v_reg  <= w_data_i[166];
      \nz.mem_165_sv2v_reg  <= w_data_i[165];
      \nz.mem_164_sv2v_reg  <= w_data_i[164];
      \nz.mem_163_sv2v_reg  <= w_data_i[163];
      \nz.mem_162_sv2v_reg  <= w_data_i[162];
      \nz.mem_161_sv2v_reg  <= w_data_i[161];
      \nz.mem_160_sv2v_reg  <= w_data_i[160];
      \nz.mem_159_sv2v_reg  <= w_data_i[159];
      \nz.mem_158_sv2v_reg  <= w_data_i[158];
      \nz.mem_157_sv2v_reg  <= w_data_i[157];
      \nz.mem_156_sv2v_reg  <= w_data_i[156];
      \nz.mem_155_sv2v_reg  <= w_data_i[155];
      \nz.mem_154_sv2v_reg  <= w_data_i[154];
      \nz.mem_153_sv2v_reg  <= w_data_i[153];
      \nz.mem_152_sv2v_reg  <= w_data_i[152];
      \nz.mem_151_sv2v_reg  <= w_data_i[151];
      \nz.mem_150_sv2v_reg  <= w_data_i[150];
      \nz.mem_149_sv2v_reg  <= w_data_i[149];
      \nz.mem_148_sv2v_reg  <= w_data_i[148];
      \nz.mem_147_sv2v_reg  <= w_data_i[147];
      \nz.mem_146_sv2v_reg  <= w_data_i[146];
      \nz.mem_145_sv2v_reg  <= w_data_i[145];
      \nz.mem_144_sv2v_reg  <= w_data_i[144];
      \nz.mem_143_sv2v_reg  <= w_data_i[143];
      \nz.mem_142_sv2v_reg  <= w_data_i[142];
      \nz.mem_141_sv2v_reg  <= w_data_i[141];
      \nz.mem_140_sv2v_reg  <= w_data_i[140];
      \nz.mem_139_sv2v_reg  <= w_data_i[139];
      \nz.mem_138_sv2v_reg  <= w_data_i[138];
      \nz.mem_137_sv2v_reg  <= w_data_i[137];
      \nz.mem_136_sv2v_reg  <= w_data_i[136];
      \nz.mem_135_sv2v_reg  <= w_data_i[135];
      \nz.mem_134_sv2v_reg  <= w_data_i[134];
      \nz.mem_133_sv2v_reg  <= w_data_i[133];
      \nz.mem_132_sv2v_reg  <= w_data_i[132];
      \nz.mem_131_sv2v_reg  <= w_data_i[131];
      \nz.mem_130_sv2v_reg  <= w_data_i[130];
      \nz.mem_129_sv2v_reg  <= w_data_i[129];
      \nz.mem_128_sv2v_reg  <= w_data_i[128];
      \nz.mem_127_sv2v_reg  <= w_data_i[127];
      \nz.mem_126_sv2v_reg  <= w_data_i[126];
      \nz.mem_125_sv2v_reg  <= w_data_i[125];
      \nz.mem_124_sv2v_reg  <= w_data_i[124];
      \nz.mem_123_sv2v_reg  <= w_data_i[123];
      \nz.mem_122_sv2v_reg  <= w_data_i[122];
      \nz.mem_121_sv2v_reg  <= w_data_i[121];
      \nz.mem_120_sv2v_reg  <= w_data_i[120];
      \nz.mem_119_sv2v_reg  <= w_data_i[119];
      \nz.mem_118_sv2v_reg  <= w_data_i[118];
      \nz.mem_117_sv2v_reg  <= w_data_i[117];
      \nz.mem_116_sv2v_reg  <= w_data_i[116];
      \nz.mem_115_sv2v_reg  <= w_data_i[115];
      \nz.mem_114_sv2v_reg  <= w_data_i[114];
      \nz.mem_113_sv2v_reg  <= w_data_i[113];
      \nz.mem_112_sv2v_reg  <= w_data_i[112];
      \nz.mem_111_sv2v_reg  <= w_data_i[111];
      \nz.mem_110_sv2v_reg  <= w_data_i[110];
      \nz.mem_109_sv2v_reg  <= w_data_i[109];
      \nz.mem_108_sv2v_reg  <= w_data_i[108];
      \nz.mem_107_sv2v_reg  <= w_data_i[107];
      \nz.mem_106_sv2v_reg  <= w_data_i[106];
      \nz.mem_105_sv2v_reg  <= w_data_i[105];
      \nz.mem_104_sv2v_reg  <= w_data_i[104];
      \nz.mem_103_sv2v_reg  <= w_data_i[103];
      \nz.mem_102_sv2v_reg  <= w_data_i[102];
      \nz.mem_101_sv2v_reg  <= w_data_i[101];
      \nz.mem_100_sv2v_reg  <= w_data_i[100];
      \nz.mem_99_sv2v_reg  <= w_data_i[99];
      \nz.mem_98_sv2v_reg  <= w_data_i[98];
      \nz.mem_97_sv2v_reg  <= w_data_i[97];
      \nz.mem_96_sv2v_reg  <= w_data_i[96];
      \nz.mem_95_sv2v_reg  <= w_data_i[95];
      \nz.mem_94_sv2v_reg  <= w_data_i[94];
      \nz.mem_93_sv2v_reg  <= w_data_i[93];
      \nz.mem_92_sv2v_reg  <= w_data_i[92];
      \nz.mem_91_sv2v_reg  <= w_data_i[91];
      \nz.mem_90_sv2v_reg  <= w_data_i[90];
      \nz.mem_89_sv2v_reg  <= w_data_i[89];
      \nz.mem_88_sv2v_reg  <= w_data_i[88];
      \nz.mem_87_sv2v_reg  <= w_data_i[87];
      \nz.mem_86_sv2v_reg  <= w_data_i[86];
      \nz.mem_85_sv2v_reg  <= w_data_i[85];
      \nz.mem_84_sv2v_reg  <= w_data_i[84];
      \nz.mem_83_sv2v_reg  <= w_data_i[83];
      \nz.mem_82_sv2v_reg  <= w_data_i[82];
      \nz.mem_81_sv2v_reg  <= w_data_i[81];
      \nz.mem_80_sv2v_reg  <= w_data_i[80];
      \nz.mem_79_sv2v_reg  <= w_data_i[79];
      \nz.mem_78_sv2v_reg  <= w_data_i[78];
      \nz.mem_77_sv2v_reg  <= w_data_i[77];
      \nz.mem_76_sv2v_reg  <= w_data_i[76];
      \nz.mem_75_sv2v_reg  <= w_data_i[75];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
    if(N35) begin
      \nz.mem_74_sv2v_reg  <= w_data_i[74];
      \nz.mem_73_sv2v_reg  <= w_data_i[73];
      \nz.mem_72_sv2v_reg  <= w_data_i[72];
      \nz.mem_71_sv2v_reg  <= w_data_i[71];
      \nz.mem_70_sv2v_reg  <= w_data_i[70];
      \nz.mem_69_sv2v_reg  <= w_data_i[69];
      \nz.mem_68_sv2v_reg  <= w_data_i[68];
      \nz.mem_67_sv2v_reg  <= w_data_i[67];
      \nz.mem_66_sv2v_reg  <= w_data_i[66];
      \nz.mem_65_sv2v_reg  <= w_data_i[65];
      \nz.mem_64_sv2v_reg  <= w_data_i[64];
      \nz.mem_63_sv2v_reg  <= w_data_i[63];
      \nz.mem_62_sv2v_reg  <= w_data_i[62];
      \nz.mem_61_sv2v_reg  <= w_data_i[61];
      \nz.mem_60_sv2v_reg  <= w_data_i[60];
      \nz.mem_59_sv2v_reg  <= w_data_i[59];
      \nz.mem_58_sv2v_reg  <= w_data_i[58];
      \nz.mem_57_sv2v_reg  <= w_data_i[57];
      \nz.mem_56_sv2v_reg  <= w_data_i[56];
      \nz.mem_55_sv2v_reg  <= w_data_i[55];
      \nz.mem_54_sv2v_reg  <= w_data_i[54];
      \nz.mem_53_sv2v_reg  <= w_data_i[53];
      \nz.mem_52_sv2v_reg  <= w_data_i[52];
      \nz.mem_51_sv2v_reg  <= w_data_i[51];
      \nz.mem_50_sv2v_reg  <= w_data_i[50];
      \nz.mem_49_sv2v_reg  <= w_data_i[49];
      \nz.mem_48_sv2v_reg  <= w_data_i[48];
      \nz.mem_47_sv2v_reg  <= w_data_i[47];
      \nz.mem_46_sv2v_reg  <= w_data_i[46];
      \nz.mem_45_sv2v_reg  <= w_data_i[45];
      \nz.mem_44_sv2v_reg  <= w_data_i[44];
      \nz.mem_43_sv2v_reg  <= w_data_i[43];
      \nz.mem_42_sv2v_reg  <= w_data_i[42];
      \nz.mem_41_sv2v_reg  <= w_data_i[41];
      \nz.mem_40_sv2v_reg  <= w_data_i[40];
      \nz.mem_39_sv2v_reg  <= w_data_i[39];
      \nz.mem_38_sv2v_reg  <= w_data_i[38];
      \nz.mem_37_sv2v_reg  <= w_data_i[37];
      \nz.mem_36_sv2v_reg  <= w_data_i[36];
      \nz.mem_35_sv2v_reg  <= w_data_i[35];
      \nz.mem_34_sv2v_reg  <= w_data_i[34];
      \nz.mem_33_sv2v_reg  <= w_data_i[33];
      \nz.mem_32_sv2v_reg  <= w_data_i[32];
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
    end 
  end


endmodule



module bsg_mem_1r1w_000000ae_00000008
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [2:0] w_addr_i;
  input [173:0] w_data_i;
  input [2:0] r_addr_i;
  output [173:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [173:0] r_data_o;

  bsg_mem_1r1w_synth_000000ae_00000008_0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bp_be_instr_decoder_00
(
  preissue_pkt_i,
  decode_info_i,
  decode_o,
  illegal_instr_o,
  ecall_m_o,
  ecall_s_o,
  ecall_u_o,
  ebreak_o,
  dbreak_o,
  dret_o,
  mret_o,
  sret_o,
  wfi_o,
  sfence_vma_o,
  fencei_o,
  csrw_o,
  imm_o
);

  input [38:0] preissue_pkt_i;
  input [12:0] decode_info_i;
  output [53:0] decode_o;
  output [63:0] imm_o;
  output illegal_instr_o;
  output ecall_m_o;
  output ecall_s_o;
  output ecall_u_o;
  output ebreak_o;
  output dbreak_o;
  output dret_o;
  output mret_o;
  output sret_o;
  output wfi_o;
  output sfence_vma_o;
  output fencei_o;
  output csrw_o;
  wire [53:0] decode_o;
  wire [63:0] imm_o;
  wire illegal_instr_o,ecall_m_o,ecall_s_o,ecall_u_o,ebreak_o,dbreak_o,dret_o,mret_o,
  sret_o,wfi_o,sfence_vma_o,fencei_o,csrw_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,
  N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,
  N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,
  N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,
  N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,
  N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,
  N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,
  N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,
  N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,
  N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,
  decode_o_45_,decode_o_44_,decode_o_43_,decode_o_42_,decode_o_41_,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,
  N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,
  N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,
  N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,
  N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,
  N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,
  N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,
  N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
  N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,
  N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
  N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,
  N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,
  N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,
  N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,
  N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,
  N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,
  N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,
  N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,
  N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,
  N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,
  N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,
  N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,
  N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,
  N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,
  N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,
  N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,
  N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,
  N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,
  N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,
  N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,
  N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,
  N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,
  N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,
  N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
  N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,
  N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,
  N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,
  N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,
  N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,
  N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,
  N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,
  N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,
  N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,
  N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,
  N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,
  N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,
  N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,
  N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,
  N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,
  N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,
  N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,
  N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,
  N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,
  N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,
  N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,
  N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,
  N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,
  N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,
  N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,
  N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,
  N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,
  N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,
  N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,
  N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,
  N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,
  N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,
  N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,
  N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,
  N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,
  N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,
  N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,
  N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,
  N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,
  N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,
  N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,
  N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,
  N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,
  N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,
  N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,
  N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,
  N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,
  N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,
  N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,
  N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
  N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,
  N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,
  N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,
  N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,
  N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,
  N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,
  N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,
  N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,
  N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,
  N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,
  N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,
  N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,
  N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,
  N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,
  N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,
  N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,
  N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,
  N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,
  N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,
  N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,
  N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,
  N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,
  N1754,N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,
  N1767,N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,
  N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,
  N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,
  N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,
  N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,
  N1834,N1835,N1836,N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,
  N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,
  N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,
  N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,
  N1887,N1888,N1889,N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,
  N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,
  N1914,N1915,N1916,N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,
  N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,
  N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,
  N1954,N1955,N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,
  N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,
  N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,
  N1994,N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,
  N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,
  N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,
  N2034,N2035,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,
  N2047,N2048,N2049,N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,
  N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,
  N2074,N2075,N2076,N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,
  N2087,N2088,N2089,N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,
  N2100,N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,
  N2114,N2115,N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,
  N2127,N2128,N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,
  N2140,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,
  N2154,N2155,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,
  N2167,N2168,N2169,N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,
  N2180,N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,
  N2194,N2195,N2196,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,
  N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,
  N2220,N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,
  N2234,N2235,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,
  N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,
  N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,
  N2274,N2275,N2276,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,
  N2287,N2288,N2289,N2290,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,
  N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,
  N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,
  N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,
  N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,
  N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,
  N2367,N2368,N2369,N2370,N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,
  N2380,N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,
  N2394,N2395,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,
  N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,
  N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,
  N2434,N2435,N2436,N2437,N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,
  N2447,N2448,N2449,N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,
  N2460,N2461,N2462,N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,
  N2474,N2475,N2476,N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,
  N2487,N2488,N2489,N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,
  N2500,N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,
  N2514,N2515,N2516,N2517,N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,
  N2527,N2528,N2529,N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,
  N2540,N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,
  N2554,N2555,N2556,N2557,N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,
  N2567,N2568,N2569,N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,
  N2580,N2581,N2582,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,
  N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,
  N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,
  N2620,N2621,N2622,N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,
  N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,
  N2647,N2648,N2649,N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,
  N2660,N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,
  N2674,N2675,N2676,N2677,N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,
  N2687,N2688,N2689,N2690,N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,
  N2700,N2701,N2702,N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,
  N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,
  N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,
  N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,
  N2754,N2755,N2756,N2757,N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,
  N2767,N2768,N2769,N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,
  N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,
  N2794,N2795,N2796,N2797,N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,
  N2807,N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,N2819,
  N2820,N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,
  N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,
  N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,N2859,
  N2860,N2861,N2862,N2863,N2864,N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,
  N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,
  N2887,N2888,N2889,N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,
  N2900,N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908;
  assign decode_o[7] = 1'b0;
  assign decode_o[19] = 1'b0;
  assign decode_o[31] = 1'b0;
  assign decode_o_45_ = preissue_pkt_i[38];
  assign decode_o[45] = decode_o_45_;
  assign decode_o_44_ = preissue_pkt_i[37];
  assign decode_o[44] = decode_o_44_;
  assign decode_o_43_ = preissue_pkt_i[36];
  assign decode_o[43] = decode_o_43_;
  assign decode_o_42_ = preissue_pkt_i[35];
  assign decode_o[42] = decode_o_42_;
  assign decode_o_41_ = preissue_pkt_i[34];
  assign decode_o[41] = decode_o_41_;
  assign N173 = preissue_pkt_i[3] & preissue_pkt_i[2];
  assign N175 = N188 | preissue_pkt_i[4];
  assign N176 = N187 | N183;
  assign N177 = N176 | preissue_pkt_i[4];
  assign N179 = preissue_pkt_i[8] | preissue_pkt_i[7];
  assign N180 = N203 | preissue_pkt_i[5];
  assign N181 = N179 | N180;
  assign N182 = N181 | preissue_pkt_i[4];
  assign N183 = N203 | N204;
  assign N184 = N179 | N183;
  assign N185 = N184 | preissue_pkt_i[4];
  assign N187 = preissue_pkt_i[8] | N202;
  assign N188 = N187 | N180;
  assign N189 = N188 | N205;
  assign N191 = N181 | N205;
  assign N193 = N197 | N235;
  assign N194 = N193 | N205;
  assign N195 = N198 | N205;
  assign N197 = N201 | N202;
  assign N198 = N197 | N212;
  assign N199 = N198 | preissue_pkt_i[4];
  assign N206 = N201 & N202;
  assign N207 = N203 & N204;
  assign N208 = N206 & N207;
  assign N209 = N208 & N205;
  assign N210 = N2568 | N205;
  assign N212 = preissue_pkt_i[6] | preissue_pkt_i[5];
  assign N213 = N187 | N212;
  assign N214 = N213 | preissue_pkt_i[4];
  assign N216 = N213 | N205;
  assign N218 = N179 | N235;
  assign N219 = N218 | N205;
  assign N221 = N197 | N180;
  assign N222 = N221 | preissue_pkt_i[4];
  assign N224 = N201 | preissue_pkt_i[7];
  assign N225 = N224 | N180;
  assign N226 = N225 | preissue_pkt_i[4];
  assign N228 = N224 | N212;
  assign N229 = N228 | preissue_pkt_i[4];
  assign N230 = N228 | N205;
  assign N231 = N224 | N235;
  assign N232 = N231 | preissue_pkt_i[4];
  assign N233 = N231 | N205;
  assign N235 = preissue_pkt_i[6] | N204;
  assign N236 = N187 | N235;
  assign N237 = N236 | N205;
  assign N239 = preissue_pkt_i[6] & preissue_pkt_i[5];
  assign N240 = N239 & preissue_pkt_i[4];
  assign N241 = preissue_pkt_i[8] & preissue_pkt_i[6];
  assign N242 = N241 & preissue_pkt_i[4];
  assign N243 = N241 & preissue_pkt_i[5];
  assign N244 = preissue_pkt_i[7] & N203;
  assign N245 = preissue_pkt_i[5] & N205;
  assign N246 = N244 & N245;
  assign N247 = N201 & N203;
  assign N248 = N247 & N245;
  assign N250 = preissue_pkt_i[16] | N526;
  assign N251 = preissue_pkt_i[15] | N250;
  assign N252 = preissue_pkt_i[14] | N251;
  assign N253 = preissue_pkt_i[8] | N252;
  assign N254 = N1328 | N253;
  assign N255 = N394 | N254;
  assign N256 = preissue_pkt_i[5] | N255;
  assign N257 = preissue_pkt_i[4] | N256;
  assign N258 = N395 | N257;
  assign N259 = N396 | N258;
  assign N260 = ~N259;
  assign N261 = N1329 | N255;
  assign N262 = preissue_pkt_i[4] | N261;
  assign N263 = N395 | N262;
  assign N264 = N396 | N263;
  assign N265 = ~N264;
  assign N266 = N260 | N265;
  assign N267 = N2305 | N251;
  assign N268 = preissue_pkt_i[8] | N267;
  assign N269 = N1328 | N268;
  assign N270 = N394 | N269;
  assign N271 = preissue_pkt_i[5] | N270;
  assign N272 = preissue_pkt_i[4] | N271;
  assign N273 = N395 | N272;
  assign N274 = N396 | N273;
  assign N275 = ~N274;
  assign N276 = N394 | N483;
  assign N277 = preissue_pkt_i[5] | N276;
  assign N278 = preissue_pkt_i[4] | N277;
  assign N279 = N395 | N278;
  assign N280 = N396 | N279;
  assign N281 = ~N280;
  assign N282 = N275 | N281;
  assign N283 = N394 | N492;
  assign N284 = preissue_pkt_i[5] | N283;
  assign N285 = preissue_pkt_i[4] | N284;
  assign N286 = N395 | N285;
  assign N287 = N396 | N286;
  assign N288 = ~N287;
  assign N289 = N282 | N288;
  assign N290 = preissue_pkt_i[5] | N305;
  assign N291 = preissue_pkt_i[4] | N290;
  assign N292 = N395 | N291;
  assign N293 = N396 | N292;
  assign N294 = ~N293;
  assign N295 = N289 | N294;
  assign N296 = preissue_pkt_i[5] | N312;
  assign N297 = preissue_pkt_i[4] | N296;
  assign N298 = N395 | N297;
  assign N299 = N396 | N298;
  assign N300 = ~N299;
  assign N301 = N295 | N300;
  assign N302 = preissue_pkt_i[14] | N506;
  assign N303 = preissue_pkt_i[8] | N302;
  assign N304 = N1328 | N303;
  assign N305 = N394 | N304;
  assign N306 = N1329 | N305;
  assign N307 = preissue_pkt_i[4] | N306;
  assign N308 = N395 | N307;
  assign N309 = N396 | N308;
  assign N310 = ~N309;
  assign N311 = N301 | N310;
  assign N312 = N394 | N509;
  assign N313 = N1329 | N312;
  assign N314 = preissue_pkt_i[4] | N313;
  assign N315 = N395 | N314;
  assign N316 = N396 | N315;
  assign N317 = ~N316;
  assign N318 = N311 | N317;
  assign N319 = preissue_pkt_i[5] | N334;
  assign N320 = preissue_pkt_i[4] | N319;
  assign N321 = N395 | N320;
  assign N322 = N396 | N321;
  assign N323 = ~N322;
  assign N324 = N318 | N323;
  assign N325 = preissue_pkt_i[5] | N341;
  assign N326 = preissue_pkt_i[4] | N325;
  assign N327 = N395 | N326;
  assign N328 = N396 | N327;
  assign N329 = ~N328;
  assign N330 = N324 | N329;
  assign N331 = preissue_pkt_i[14] | N528;
  assign N332 = preissue_pkt_i[8] | N331;
  assign N333 = N1328 | N332;
  assign N334 = N394 | N333;
  assign N335 = N1329 | N334;
  assign N336 = preissue_pkt_i[4] | N335;
  assign N337 = N395 | N336;
  assign N338 = N396 | N337;
  assign N339 = ~N338;
  assign N340 = N330 | N339;
  assign N341 = N394 | N531;
  assign N342 = N1329 | N341;
  assign N343 = preissue_pkt_i[4] | N342;
  assign N344 = N395 | N343;
  assign N345 = N396 | N344;
  assign N346 = ~N345;
  assign N347 = N340 | N346;
  assign N350 = preissue_pkt_i[16] | N402;
  assign N351 = preissue_pkt_i[15] | N350;
  assign N352 = preissue_pkt_i[14] | N351;
  assign N353 = preissue_pkt_i[8] | N352;
  assign N354 = N1328 | N353;
  assign N355 = N394 | N354;
  assign N356 = N1329 | N355;
  assign N357 = preissue_pkt_i[4] | N356;
  assign N358 = N395 | N357;
  assign N359 = N396 | N358;
  assign N360 = ~N359;
  assign N361 = preissue_pkt_i[16] | N974;
  assign N362 = N2304 | N361;
  assign N363 = preissue_pkt_i[14] | N362;
  assign N364 = preissue_pkt_i[8] | N363;
  assign N365 = N1328 | N364;
  assign N366 = N394 | N365;
  assign N367 = N1329 | N366;
  assign N368 = preissue_pkt_i[4] | N367;
  assign N369 = N395 | N368;
  assign N370 = N396 | N369;
  assign N371 = ~N370;
  assign N372 = N360 | N371;
  assign N373 = preissue_pkt_i[15] | N975;
  assign N374 = preissue_pkt_i[14] | N373;
  assign N375 = preissue_pkt_i[8] | N374;
  assign N376 = N1328 | N375;
  assign N377 = N394 | N376;
  assign N378 = N1329 | N377;
  assign N379 = preissue_pkt_i[4] | N378;
  assign N380 = N395 | N379;
  assign N381 = N396 | N380;
  assign N382 = ~N381;
  assign N383 = N372 | N382;
  assign N384 = N394 | N979;
  assign N385 = N1329 | N384;
  assign N386 = preissue_pkt_i[4] | N385;
  assign N387 = N395 | N386;
  assign N388 = N396 | N387;
  assign N389 = ~N388;
  assign N390 = N383 | N389;
  assign N393 = ~preissue_pkt_i[29];
  assign N394 = ~preissue_pkt_i[6];
  assign N395 = ~preissue_pkt_i[3];
  assign N396 = ~preissue_pkt_i[2];
  assign N397 = preissue_pkt_i[32] | preissue_pkt_i[33];
  assign N398 = preissue_pkt_i[31] | N397;
  assign N399 = preissue_pkt_i[30] | N398;
  assign N400 = N393 | N399;
  assign N401 = preissue_pkt_i[28] | N400;
  assign N402 = preissue_pkt_i[27] | N401;
  assign N403 = N1631 | N402;
  assign N404 = preissue_pkt_i[15] | N403;
  assign N405 = preissue_pkt_i[14] | N404;
  assign N406 = preissue_pkt_i[8] | N405;
  assign N407 = N1328 | N406;
  assign N408 = N394 | N407;
  assign N409 = N1329 | N408;
  assign N410 = preissue_pkt_i[4] | N409;
  assign N411 = N395 | N410;
  assign N412 = N396 | N411;
  assign N413 = ~N412;
  assign N415 = N288 | N300;
  assign N416 = N415 | N317;
  assign N417 = N416 | N329;
  assign N418 = N417 | N346;
  assign N419 = preissue_pkt_i[5] | N425;
  assign N420 = preissue_pkt_i[4] | N419;
  assign N421 = N395 | N420;
  assign N422 = N396 | N421;
  assign N423 = ~N422;
  assign N424 = N418 | N423;
  assign N425 = N394 | N860;
  assign N426 = N1329 | N425;
  assign N427 = preissue_pkt_i[4] | N426;
  assign N428 = N395 | N427;
  assign N429 = N396 | N428;
  assign N430 = ~N429;
  assign N431 = N424 | N430;
  assign N432 = N431 | N360;
  assign N433 = N432 | N371;
  assign N434 = N433 | N382;
  assign N435 = N434 | N389;
  assign N436 = N394 | N407;
  assign N437 = N1329 | N436;
  assign N438 = preissue_pkt_i[4] | N437;
  assign N439 = N395 | N438;
  assign N440 = N396 | N439;
  assign N441 = ~N440;
  assign N442 = N435 | N441;
  assign N443 = preissue_pkt_i[5] | N449;
  assign N444 = preissue_pkt_i[4] | N443;
  assign N445 = N395 | N444;
  assign N446 = N396 | N445;
  assign N447 = ~N446;
  assign N448 = N442 | N447;
  assign N449 = N394 | N914;
  assign N450 = N1329 | N449;
  assign N451 = preissue_pkt_i[4] | N450;
  assign N452 = N395 | N451;
  assign N453 = N396 | N452;
  assign N454 = ~N453;
  assign N455 = N448 | N454;
  assign N456 = preissue_pkt_i[5] | N473;
  assign N457 = preissue_pkt_i[4] | N456;
  assign N458 = N395 | N457;
  assign N459 = N396 | N458;
  assign N460 = ~N459;
  assign N461 = N455 | N460;
  assign N462 = ~preissue_pkt_i[31];
  assign N463 = N462 | N1288;
  assign N464 = preissue_pkt_i[30] | N463;
  assign N465 = preissue_pkt_i[29] | N464;
  assign N466 = preissue_pkt_i[28] | N465;
  assign N467 = preissue_pkt_i[27] | N466;
  assign N468 = preissue_pkt_i[16] | N467;
  assign N469 = preissue_pkt_i[15] | N468;
  assign N470 = N2305 | N469;
  assign N471 = preissue_pkt_i[8] | N470;
  assign N472 = N1328 | N471;
  assign N473 = N394 | N472;
  assign N474 = N1329 | N473;
  assign N475 = preissue_pkt_i[4] | N474;
  assign N476 = N395 | N475;
  assign N477 = N396 | N476;
  assign N478 = ~N477;
  assign N479 = N461 | N478;
  assign N480 = N2304 | N250;
  assign N481 = preissue_pkt_i[14] | N480;
  assign N482 = preissue_pkt_i[8] | N481;
  assign N483 = N1328 | N482;
  assign N484 = N394 | N483;
  assign N485 = preissue_pkt_i[5] | N484;
  assign N486 = preissue_pkt_i[4] | N485;
  assign N487 = N395 | N486;
  assign N488 = N396 | N487;
  assign N489 = ~N488;
  assign N490 = N2305 | N480;
  assign N491 = preissue_pkt_i[8] | N490;
  assign N492 = N1328 | N491;
  assign N493 = N394 | N492;
  assign N494 = preissue_pkt_i[5] | N493;
  assign N495 = preissue_pkt_i[4] | N494;
  assign N496 = N395 | N495;
  assign N497 = N396 | N496;
  assign N498 = ~N497;
  assign N499 = N489 | N498;
  assign N500 = preissue_pkt_i[5] | N510;
  assign N501 = preissue_pkt_i[4] | N500;
  assign N502 = N395 | N501;
  assign N503 = N396 | N502;
  assign N504 = ~N503;
  assign N505 = N499 | N504;
  assign N506 = preissue_pkt_i[15] | N527;
  assign N507 = N2305 | N506;
  assign N508 = preissue_pkt_i[8] | N507;
  assign N509 = N1328 | N508;
  assign N510 = N394 | N509;
  assign N511 = N1329 | N510;
  assign N512 = preissue_pkt_i[4] | N511;
  assign N513 = N395 | N512;
  assign N514 = N396 | N513;
  assign N515 = ~N514;
  assign N516 = N505 | N515;
  assign N517 = preissue_pkt_i[5] | N532;
  assign N518 = preissue_pkt_i[4] | N517;
  assign N519 = N395 | N518;
  assign N520 = N396 | N519;
  assign N521 = ~N520;
  assign N522 = N516 | N521;
  assign N523 = ~preissue_pkt_i[27];
  assign N524 = preissue_pkt_i[29] | N399;
  assign N525 = preissue_pkt_i[28] | N524;
  assign N526 = N523 | N525;
  assign N527 = N1631 | N526;
  assign N528 = N2304 | N527;
  assign N529 = N2305 | N528;
  assign N530 = preissue_pkt_i[8] | N529;
  assign N531 = N1328 | N530;
  assign N532 = N394 | N531;
  assign N533 = N1329 | N532;
  assign N534 = preissue_pkt_i[4] | N533;
  assign N535 = N395 | N534;
  assign N536 = N396 | N535;
  assign N537 = ~N536;
  assign N538 = N522 | N537;
  assign N539 = N2135 & N2303;
  assign N540 = N2684 & N1327;
  assign N541 = N1330 & preissue_pkt_i[3];
  assign N542 = N539 & N540;
  assign N543 = N2573 & N541;
  assign N544 = N542 & N543;
  assign N545 = N544 & preissue_pkt_i[2];
  assign N547 = N2305 & N1329;
  assign N548 = N617 & N547;
  assign N549 = N585 & N548;
  assign N550 = N2305 & preissue_pkt_i[5];
  assign N551 = N617 & N550;
  assign N552 = N585 & N551;
  assign N553 = N581 & N616;
  assign N554 = N553 & N551;
  assign N555 = preissue_pkt_i[32] & N462;
  assign N556 = N555 & N582;
  assign N557 = N617 & N584;
  assign N558 = N556 & N557;
  assign N559 = N617 & N697;
  assign N560 = N556 & N559;
  assign N561 = N585 & N619;
  assign N562 = N617 & N651;
  assign N563 = N585 & N562;
  assign N564 = N585 & N595;
  assign N565 = N1357 & N651;
  assign N566 = N585 & N565;
  assign N567 = N625 & N582;
  assign N568 = N567 & N586;
  assign N569 = N583 & N697;
  assign N570 = N567 & N569;
  assign N571 = N567 & N593;
  assign N572 = N1357 & N697;
  assign N573 = N567 & N572;
  assign N574 = N567 & N597;
  assign N575 = N1360 & N697;
  assign N576 = N567 & N575;
  assign N577 = N553 & N572;
  assign N578 = N556 & N595;
  assign N579 = N556 & N565;
  assign N581 = N1287 & N462;
  assign N582 = N393 & N523;
  assign N583 = N1631 & preissue_pkt_i[15];
  assign N584 = N2305 & N1329;
  assign N585 = N581 & N582;
  assign N586 = N583 & N584;
  assign N587 = N585 & N586;
  assign N588 = preissue_pkt_i[14] & N1329;
  assign N589 = N583 & N588;
  assign N590 = N585 & N589;
  assign N591 = preissue_pkt_i[29] & preissue_pkt_i[27];
  assign N592 = N581 & N591;
  assign N593 = N1357 & N584;
  assign N594 = N592 & N593;
  assign N595 = N1357 & N588;
  assign N596 = N592 & N595;
  assign N597 = N1360 & N584;
  assign N598 = N592 & N597;
  assign N599 = N1360 & N588;
  assign N600 = N592 & N599;
  assign N601 = N585 & N593;
  assign N602 = N556 & N593;
  assign N604 = N622 & N582;
  assign N605 = N604 & N619;
  assign N606 = N604 & N562;
  assign N607 = N604 & N595;
  assign N608 = N604 & N565;
  assign N609 = N585 & N597;
  assign N610 = N556 & N597;
  assign N612 = N585 & N599;
  assign N613 = N556 & N599;
  assign N615 = preissue_pkt_i[32] & N462;
  assign N616 = preissue_pkt_i[29] & N523;
  assign N617 = N1631 & N2304;
  assign N618 = N615 & N616;
  assign N619 = N617 & N588;
  assign N620 = N618 & N619;
  assign N621 = N618 & N595;
  assign N622 = preissue_pkt_i[32] & preissue_pkt_i[31];
  assign N623 = N622 & N616;
  assign N624 = N623 & N619;
  assign N625 = N1287 & preissue_pkt_i[31];
  assign N626 = N625 & N616;
  assign N627 = N626 & N619;
  assign N628 = N633 & N557;
  assign N629 = N633 & N559;
  assign N631 = N1287 & N462;
  assign N632 = N393 & preissue_pkt_i[27];
  assign N633 = N631 & N632;
  assign N634 = N633 & N619;
  assign N635 = N633 & N586;
  assign N636 = N633 & N589;
  assign N637 = N633 & N593;
  assign N638 = N633 & N572;
  assign N640 = N633 & N595;
  assign N641 = N633 & N565;
  assign N643 = N633 & N597;
  assign N644 = N633 & N575;
  assign N646 = N633 & N599;
  assign N647 = N1360 & N651;
  assign N648 = N633 & N647;
  assign N650 = N523 & preissue_pkt_i[15];
  assign N651 = preissue_pkt_i[14] & preissue_pkt_i[5];
  assign N652 = N650 & N651;
  assign N653 = N1287 & preissue_pkt_i[29];
  assign N654 = N523 & preissue_pkt_i[16];
  assign N655 = N653 & N654;
  assign N656 = N655 & preissue_pkt_i[14];
  assign N657 = preissue_pkt_i[16] & preissue_pkt_i[14];
  assign N658 = N2458 & N657;
  assign N659 = N1287 & preissue_pkt_i[31];
  assign N660 = N659 & N657;
  assign N661 = preissue_pkt_i[31] & preissue_pkt_i[15];
  assign N662 = N661 & preissue_pkt_i[14];
  assign N663 = N393 & preissue_pkt_i[14];
  assign N664 = N659 & N663;
  assign N665 = N583 & N651;
  assign N666 = N615 & N672;
  assign N667 = N666 & preissue_pkt_i[5];
  assign N668 = preissue_pkt_i[29] & preissue_pkt_i[14];
  assign N669 = N668 & preissue_pkt_i[5];
  assign N670 = preissue_pkt_i[27] & N1631;
  assign N671 = N670 & N651;
  assign N672 = N1631 & preissue_pkt_i[14];
  assign N673 = N591 & N672;
  assign N674 = N631 & N688;
  assign N675 = N674 & preissue_pkt_i[14];
  assign N676 = N393 & N1631;
  assign N677 = N615 & N676;
  assign N678 = N677 & preissue_pkt_i[14];
  assign N679 = preissue_pkt_i[29] & preissue_pkt_i[15];
  assign N680 = N679 & preissue_pkt_i[5];
  assign N681 = N616 & preissue_pkt_i[15];
  assign N682 = N622 & preissue_pkt_i[15];
  assign N683 = N462 & N523;
  assign N684 = preissue_pkt_i[15] & preissue_pkt_i[5];
  assign N685 = N683 & N684;
  assign N686 = preissue_pkt_i[32] & N1631;
  assign N687 = N686 & preissue_pkt_i[15];
  assign N688 = preissue_pkt_i[29] & N1631;
  assign N689 = N688 & preissue_pkt_i[15];
  assign N690 = N462 & N1631;
  assign N691 = N690 & N684;
  assign N692 = preissue_pkt_i[32] & preissue_pkt_i[16];
  assign N693 = N692 & N1410;
  assign N694 = N693 & preissue_pkt_i[5];
  assign N695 = N2458 & preissue_pkt_i[5];
  assign N696 = N462 & N393;
  assign N697 = N2305 & preissue_pkt_i[5];
  assign N698 = N696 & N654;
  assign N699 = N698 & N697;
  assign N700 = N591 & preissue_pkt_i[5];
  assign N701 = N2460 & preissue_pkt_i[5];
  assign N702 = preissue_pkt_i[31] & preissue_pkt_i[27];
  assign N703 = N616 & N584;
  assign N704 = N622 & N584;
  assign N705 = preissue_pkt_i[31] & N1631;
  assign N706 = N705 & N1410;
  assign N707 = N688 & N584;
  assign N708 = preissue_pkt_i[32] & preissue_pkt_i[27];
  assign N722 = preissue_pkt_i[16] | N2036;
  assign N723 = preissue_pkt_i[15] | N722;
  assign N724 = preissue_pkt_i[14] | N723;
  assign N725 = preissue_pkt_i[8] | N724;
  assign N726 = N1328 | N725;
  assign N727 = N394 | N726;
  assign N728 = preissue_pkt_i[5] | N727;
  assign N729 = preissue_pkt_i[4] | N728;
  assign N730 = N395 | N729;
  assign N731 = N396 | N730;
  assign N732 = ~N731;
  assign N733 = N1329 | N727;
  assign N734 = preissue_pkt_i[4] | N733;
  assign N735 = N395 | N734;
  assign N736 = N396 | N735;
  assign N737 = ~N736;
  assign N738 = N732 | N737;
  assign N739 = preissue_pkt_i[14] | N749;
  assign N740 = preissue_pkt_i[8] | N739;
  assign N741 = N1328 | N740;
  assign N742 = N394 | N741;
  assign N743 = preissue_pkt_i[5] | N742;
  assign N744 = preissue_pkt_i[4] | N743;
  assign N745 = N395 | N744;
  assign N746 = N396 | N745;
  assign N747 = ~N746;
  assign N748 = N738 | N747;
  assign N749 = N2304 | N836;
  assign N750 = N2305 | N749;
  assign N751 = preissue_pkt_i[8] | N750;
  assign N752 = N1328 | N751;
  assign N753 = N394 | N752;
  assign N754 = preissue_pkt_i[5] | N753;
  assign N755 = preissue_pkt_i[4] | N754;
  assign N756 = N395 | N755;
  assign N757 = N396 | N756;
  assign N758 = ~N757;
  assign N759 = N748 | N758;
  assign N760 = preissue_pkt_i[14] | N770;
  assign N761 = preissue_pkt_i[8] | N760;
  assign N762 = N1328 | N761;
  assign N763 = N394 | N762;
  assign N764 = preissue_pkt_i[5] | N763;
  assign N765 = preissue_pkt_i[4] | N764;
  assign N766 = N395 | N765;
  assign N767 = N396 | N766;
  assign N768 = ~N767;
  assign N769 = N759 | N768;
  assign N770 = preissue_pkt_i[15] | N792;
  assign N771 = N2305 | N770;
  assign N772 = preissue_pkt_i[8] | N771;
  assign N773 = N1328 | N772;
  assign N774 = N394 | N773;
  assign N775 = preissue_pkt_i[5] | N774;
  assign N776 = preissue_pkt_i[4] | N775;
  assign N777 = N395 | N776;
  assign N778 = N396 | N777;
  assign N779 = ~N778;
  assign N780 = N769 | N779;
  assign N781 = preissue_pkt_i[14] | N793;
  assign N782 = preissue_pkt_i[8] | N781;
  assign N783 = N1328 | N782;
  assign N784 = N394 | N783;
  assign N785 = preissue_pkt_i[5] | N784;
  assign N786 = preissue_pkt_i[4] | N785;
  assign N787 = N395 | N786;
  assign N788 = N396 | N787;
  assign N789 = ~N788;
  assign N790 = N780 | N789;
  assign N791 = N523 | N401;
  assign N792 = N1631 | N791;
  assign N793 = N2304 | N792;
  assign N794 = N2305 | N793;
  assign N795 = preissue_pkt_i[8] | N794;
  assign N796 = N1328 | N795;
  assign N797 = N394 | N796;
  assign N798 = preissue_pkt_i[5] | N797;
  assign N799 = preissue_pkt_i[4] | N798;
  assign N800 = N395 | N799;
  assign N801 = N396 | N800;
  assign N802 = ~N801;
  assign N803 = N790 | N802;
  assign N804 = N2304 | N879;
  assign N805 = N2305 | N804;
  assign N806 = preissue_pkt_i[8] | N805;
  assign N807 = N1328 | N806;
  assign N808 = N394 | N807;
  assign N809 = preissue_pkt_i[5] | N808;
  assign N810 = preissue_pkt_i[4] | N809;
  assign N811 = N395 | N810;
  assign N812 = N396 | N811;
  assign N813 = ~N812;
  assign N814 = preissue_pkt_i[14] | N804;
  assign N815 = preissue_pkt_i[8] | N814;
  assign N816 = N1328 | N815;
  assign N817 = N394 | N816;
  assign N818 = preissue_pkt_i[5] | N817;
  assign N819 = preissue_pkt_i[4] | N818;
  assign N820 = N395 | N819;
  assign N821 = N396 | N820;
  assign N822 = ~N821;
  assign N823 = N813 | N822;
  assign N824 = preissue_pkt_i[14] | N880;
  assign N825 = preissue_pkt_i[8] | N824;
  assign N826 = N1328 | N825;
  assign N827 = N394 | N826;
  assign N828 = preissue_pkt_i[5] | N827;
  assign N829 = preissue_pkt_i[4] | N828;
  assign N830 = N395 | N829;
  assign N831 = N396 | N830;
  assign N832 = ~N831;
  assign N833 = N823 | N832;
  assign N836 = preissue_pkt_i[16] | N1809;
  assign N837 = preissue_pkt_i[15] | N836;
  assign N838 = N2305 | N837;
  assign N839 = preissue_pkt_i[8] | N838;
  assign N840 = N1328 | N839;
  assign N841 = N394 | N840;
  assign N842 = preissue_pkt_i[5] | N841;
  assign N843 = preissue_pkt_i[4] | N842;
  assign N844 = N395 | N843;
  assign N845 = N396 | N844;
  assign N846 = ~N845;
  assign N847 = N1329 | N841;
  assign N848 = preissue_pkt_i[4] | N847;
  assign N849 = N395 | N848;
  assign N850 = N396 | N849;
  assign N851 = ~N850;
  assign N852 = N846 | N851;
  assign N856 = N1631 | N1809;
  assign N857 = preissue_pkt_i[15] | N856;
  assign N858 = N2305 | N857;
  assign N859 = preissue_pkt_i[8] | N858;
  assign N860 = N1328 | N859;
  assign N861 = N394 | N860;
  assign N862 = preissue_pkt_i[5] | N861;
  assign N863 = preissue_pkt_i[4] | N862;
  assign N864 = N395 | N863;
  assign N865 = N396 | N864;
  assign N866 = ~N865;
  assign N867 = N1329 | N861;
  assign N868 = preissue_pkt_i[4] | N867;
  assign N869 = N395 | N868;
  assign N870 = N396 | N869;
  assign N871 = ~N870;
  assign N872 = N866 | N871;
  assign N873 = preissue_pkt_i[5] | N884;
  assign N874 = preissue_pkt_i[4] | N873;
  assign N875 = N395 | N874;
  assign N876 = N396 | N875;
  assign N877 = ~N876;
  assign N878 = N872 | N877;
  assign N879 = N1631 | N2036;
  assign N880 = preissue_pkt_i[15] | N879;
  assign N881 = N2305 | N880;
  assign N882 = preissue_pkt_i[8] | N881;
  assign N883 = N1328 | N882;
  assign N884 = N394 | N883;
  assign N885 = N1329 | N884;
  assign N886 = preissue_pkt_i[4] | N885;
  assign N887 = N395 | N886;
  assign N888 = N396 | N887;
  assign N889 = ~N888;
  assign N890 = N878 | N889;
  assign N896 = N394 | N472;
  assign N897 = preissue_pkt_i[5] | N896;
  assign N898 = preissue_pkt_i[4] | N897;
  assign N899 = N395 | N898;
  assign N900 = N396 | N899;
  assign N901 = ~N900;
  assign N902 = N1329 | N896;
  assign N903 = preissue_pkt_i[4] | N902;
  assign N904 = N395 | N903;
  assign N905 = N396 | N904;
  assign N906 = ~N905;
  assign N907 = N901 | N906;
  assign N914 = N1328 | N1249;
  assign N915 = N394 | N914;
  assign N916 = preissue_pkt_i[5] | N915;
  assign N917 = preissue_pkt_i[4] | N916;
  assign N918 = N395 | N917;
  assign N919 = N396 | N918;
  assign N920 = ~N919;
  assign N921 = N1329 | N915;
  assign N922 = preissue_pkt_i[4] | N921;
  assign N923 = N395 | N922;
  assign N924 = N396 | N923;
  assign N925 = ~N924;
  assign N926 = N920 | N925;
  assign N933 = N395 | N410;
  assign N934 = N396 | N933;
  assign N935 = ~N934;
  assign N939 = N394 | N365;
  assign N940 = preissue_pkt_i[5] | N939;
  assign N941 = preissue_pkt_i[4] | N940;
  assign N942 = N395 | N941;
  assign N943 = N396 | N942;
  assign N944 = ~N943;
  assign N945 = N1329 | N939;
  assign N946 = preissue_pkt_i[4] | N945;
  assign N947 = N395 | N946;
  assign N948 = N396 | N947;
  assign N949 = ~N948;
  assign N950 = N944 | N949;
  assign N951 = preissue_pkt_i[5] | N957;
  assign N952 = preissue_pkt_i[4] | N951;
  assign N953 = N395 | N952;
  assign N954 = N396 | N953;
  assign N955 = ~N954;
  assign N956 = N950 | N955;
  assign N957 = N394 | N376;
  assign N958 = N1329 | N957;
  assign N959 = preissue_pkt_i[4] | N958;
  assign N960 = N395 | N959;
  assign N961 = N396 | N960;
  assign N962 = ~N961;
  assign N963 = N956 | N962;
  assign N964 = preissue_pkt_i[5] | N980;
  assign N965 = preissue_pkt_i[4] | N964;
  assign N966 = N395 | N965;
  assign N967 = N396 | N966;
  assign N968 = ~N967;
  assign N969 = N963 | N968;
  assign N970 = N462 | N397;
  assign N971 = preissue_pkt_i[30] | N970;
  assign N972 = preissue_pkt_i[29] | N971;
  assign N973 = preissue_pkt_i[28] | N972;
  assign N974 = preissue_pkt_i[27] | N973;
  assign N975 = N1631 | N974;
  assign N976 = N2304 | N975;
  assign N977 = preissue_pkt_i[14] | N976;
  assign N978 = preissue_pkt_i[8] | N977;
  assign N979 = N1328 | N978;
  assign N980 = N394 | N979;
  assign N981 = N1329 | N980;
  assign N982 = preissue_pkt_i[4] | N981;
  assign N983 = N395 | N982;
  assign N984 = N396 | N983;
  assign N985 = ~N984;
  assign N986 = N969 | N985;
  assign N991 = preissue_pkt_i[16] | N401;
  assign N992 = preissue_pkt_i[15] | N991;
  assign N993 = N2305 | N992;
  assign N994 = preissue_pkt_i[8] | N993;
  assign N995 = preissue_pkt_i[7] | N994;
  assign N996 = N394 | N995;
  assign N997 = N1329 | N996;
  assign N998 = preissue_pkt_i[4] | N997;
  assign N999 = N395 | N998;
  assign N1000 = N396 | N999;
  assign N1001 = ~N1000;
  assign N1003 = N1011 & N2339;
  assign N1004 = N1003 & N1016;
  assign N1005 = N1018 & N1004;
  assign N1006 = N1005 & N1020;
  assign N1007 = N2135 & preissue_pkt_i[32];
  assign N1008 = preissue_pkt_i[31] & N2303;
  assign N1009 = N393 & N2684;
  assign N1010 = N523 & N2685;
  assign N1011 = N2686 & preissue_pkt_i[24];
  assign N1012 = N2079 & preissue_pkt_i[22];
  assign N1013 = N1007 & N1008;
  assign N1014 = N1009 & N1010;
  assign N1015 = N1011 & N1012;
  assign N1016 = N1354 & N2384;
  assign N1017 = N1870 & N2290;
  assign N1018 = N1013 & N1014;
  assign N1019 = N1015 & N1016;
  assign N1020 = N1017 & N173;
  assign N1021 = N1018 & N1019;
  assign N1022 = N1021 & N1020;
  assign N1027 = preissue_pkt_i[6] & N1330;
  assign N1028 = N1426 & N1027;
  assign N1029 = N1028 & N173;
  assign N1031 = N1354 & N584;
  assign N1032 = N1354 & N697;
  assign N1033 = N462 & N2303;
  assign N1034 = N1973 & N1033;
  assign N1035 = N1009 & N1354;
  assign N1036 = N1034 & N1035;
  assign N1037 = N1036 & N588;
  assign N1038 = N1036 & N651;
  assign N1039 = N1034 & N1103;
  assign N1040 = N1039 & N651;
  assign N1041 = N1034 & N1055;
  assign N1042 = N1041 & N588;
  assign N1043 = N1041 & N651;
  assign N1044 = N1003 & N1069;
  assign N1045 = N1018 & N1044;
  assign N1046 = N1015 & N1069;
  assign N1047 = N1018 & N1046;
  assign N1048 = N1007 & N1033;
  assign N1049 = N1048 & N1055;
  assign N1050 = N1049 & N588;
  assign N1051 = N1049 & N651;
  assign N1053 = N1363 & N584;
  assign N1054 = N1363 & N588;
  assign N1055 = N1009 & N1357;
  assign N1056 = N1013 & N1055;
  assign N1057 = N1056 & N588;
  assign N1058 = N1009 & N654;
  assign N1059 = N1411 & preissue_pkt_i[5];
  assign N1060 = N1013 & N1058;
  assign N1061 = N1060 & N1059;
  assign N1063 = N1461 & N1069;
  assign N1064 = N1018 & N1063;
  assign N1065 = N1461 & N1072;
  assign N1066 = N1018 & N1065;
  assign N1068 = N2383 & N1012;
  assign N1069 = N1354 & N588;
  assign N1070 = N1068 & N1069;
  assign N1071 = N1018 & N1070;
  assign N1072 = N1354 & N651;
  assign N1073 = N1068 & N1072;
  assign N1074 = N1018 & N1073;
  assign N1075 = N2383 & N2339;
  assign N1076 = N1075 & N1069;
  assign N1077 = N1018 & N1076;
  assign N1078 = N1075 & N1072;
  assign N1079 = N1018 & N1078;
  assign N1081 = preissue_pkt_i[23] & preissue_pkt_i[22];
  assign N1082 = N1102 & N1010;
  assign N1083 = N1011 & N1081;
  assign N1084 = N1928 & N1082;
  assign N1085 = N1083 & N595;
  assign N1086 = N1084 & N1085;
  assign N1087 = preissue_pkt_i[27] & preissue_pkt_i[26];
  assign N1088 = preissue_pkt_i[25] & N1183;
  assign N1089 = N1102 & N1087;
  assign N1090 = N1088 & N2339;
  assign N1091 = N1099 & N1089;
  assign N1092 = N1090 & N595;
  assign N1093 = N1091 & N1092;
  assign N1094 = N1874 & N1103;
  assign N1095 = N1094 & N588;
  assign N1096 = N1102 & N1357;
  assign N1097 = N1874 & N1096;
  assign N1098 = N1097 & N588;
  assign N1099 = N1007 & N2005;
  assign N1100 = N1099 & N1103;
  assign N1101 = N1100 & N588;
  assign N1102 = preissue_pkt_i[29] & N2684;
  assign N1103 = N1102 & N1354;
  assign N1104 = N1928 & N1103;
  assign N1105 = N1104 & N588;
  assign N1132 = preissue_pkt_i[26] | N467;
  assign N1133 = preissue_pkt_i[25] | N1132;
  assign N1134 = preissue_pkt_i[24] | N1133;
  assign N1135 = preissue_pkt_i[23] | N1134;
  assign N1136 = N2035 | N1135;
  assign N1137 = preissue_pkt_i[16] | N1136;
  assign N1138 = preissue_pkt_i[15] | N1137;
  assign N1139 = N2305 | N1138;
  assign N1140 = preissue_pkt_i[8] | N1139;
  assign N1141 = preissue_pkt_i[7] | N1140;
  assign N1142 = N394 | N1141;
  assign N1143 = preissue_pkt_i[5] | N1142;
  assign N1144 = preissue_pkt_i[4] | N1143;
  assign N1145 = N395 | N1144;
  assign N1146 = N396 | N1145;
  assign N1147 = ~N1146;
  assign N1148 = N1329 | N1142;
  assign N1149 = preissue_pkt_i[4] | N1148;
  assign N1150 = N395 | N1149;
  assign N1151 = N396 | N1150;
  assign N1152 = ~N1151;
  assign N1153 = N1147 | N1152;
  assign N1154 = N1280 | N1001;
  assign N1155 = N2079 | N1134;
  assign N1156 = preissue_pkt_i[22] | N1155;
  assign N1157 = preissue_pkt_i[16] | N1156;
  assign N1158 = preissue_pkt_i[15] | N1157;
  assign N1159 = N2305 | N1158;
  assign N1160 = preissue_pkt_i[8] | N1159;
  assign N1161 = preissue_pkt_i[7] | N1160;
  assign N1162 = N394 | N1161;
  assign N1163 = N1329 | N1162;
  assign N1164 = preissue_pkt_i[4] | N1163;
  assign N1165 = N395 | N1164;
  assign N1166 = N396 | N1165;
  assign N1167 = ~N1166;
  assign N1168 = N1154 | N1167;
  assign N1169 = preissue_pkt_i[22] | N1135;
  assign N1170 = preissue_pkt_i[16] | N1169;
  assign N1171 = preissue_pkt_i[15] | N1170;
  assign N1172 = N2305 | N1171;
  assign N1173 = preissue_pkt_i[8] | N1172;
  assign N1174 = preissue_pkt_i[7] | N1173;
  assign N1175 = N394 | N1174;
  assign N1176 = N1329 | N1175;
  assign N1177 = preissue_pkt_i[4] | N1176;
  assign N1178 = N395 | N1177;
  assign N1179 = N396 | N1178;
  assign N1180 = ~N1179;
  assign N1181 = N1168 | N1180;
  assign N1182 = N1181 | N1152;
  assign N1183 = ~preissue_pkt_i[24];
  assign N1184 = N1183 | N1133;
  assign N1185 = preissue_pkt_i[23] | N1184;
  assign N1186 = preissue_pkt_i[22] | N1185;
  assign N1187 = preissue_pkt_i[16] | N1186;
  assign N1188 = preissue_pkt_i[15] | N1187;
  assign N1189 = N2305 | N1188;
  assign N1190 = preissue_pkt_i[8] | N1189;
  assign N1191 = preissue_pkt_i[7] | N1190;
  assign N1192 = N394 | N1191;
  assign N1193 = preissue_pkt_i[5] | N1192;
  assign N1194 = preissue_pkt_i[4] | N1193;
  assign N1195 = N395 | N1194;
  assign N1196 = N396 | N1195;
  assign N1197 = ~N1196;
  assign N1198 = N2035 | N1185;
  assign N1199 = preissue_pkt_i[16] | N1198;
  assign N1200 = preissue_pkt_i[15] | N1199;
  assign N1201 = N2305 | N1200;
  assign N1202 = preissue_pkt_i[8] | N1201;
  assign N1203 = preissue_pkt_i[7] | N1202;
  assign N1204 = N394 | N1203;
  assign N1205 = preissue_pkt_i[5] | N1204;
  assign N1206 = preissue_pkt_i[4] | N1205;
  assign N1207 = N395 | N1206;
  assign N1208 = N396 | N1207;
  assign N1209 = ~N1208;
  assign N1210 = N1197 | N1209;
  assign N1213 = preissue_pkt_i[16] | N525;
  assign N1214 = preissue_pkt_i[15] | N1213;
  assign N1215 = N2305 | N1214;
  assign N1216 = preissue_pkt_i[8] | N1215;
  assign N1217 = preissue_pkt_i[7] | N1216;
  assign N1218 = N394 | N1217;
  assign N1219 = preissue_pkt_i[5] | N1218;
  assign N1220 = preissue_pkt_i[4] | N1219;
  assign N1221 = N395 | N1220;
  assign N1222 = N396 | N1221;
  assign N1223 = ~N1222;
  assign N1224 = N1329 | N1218;
  assign N1225 = preissue_pkt_i[4] | N1224;
  assign N1226 = N395 | N1225;
  assign N1227 = N396 | N1226;
  assign N1228 = ~N1227;
  assign N1229 = N1223 | N1228;
  assign N1230 = N1229 | N1001;
  assign N1235 = N1631 | N466;
  assign N1236 = preissue_pkt_i[15] | N1235;
  assign N1237 = N2305 | N1236;
  assign N1238 = preissue_pkt_i[8] | N1237;
  assign N1239 = preissue_pkt_i[7] | N1238;
  assign N1240 = N394 | N1239;
  assign N1241 = preissue_pkt_i[5] | N1240;
  assign N1242 = preissue_pkt_i[4] | N1241;
  assign N1243 = N395 | N1242;
  assign N1244 = N396 | N1243;
  assign N1245 = ~N1244;
  assign N1246 = N1631 | N467;
  assign N1247 = preissue_pkt_i[15] | N1246;
  assign N1248 = N2305 | N1247;
  assign N1249 = preissue_pkt_i[8] | N1248;
  assign N1250 = preissue_pkt_i[7] | N1249;
  assign N1251 = N394 | N1250;
  assign N1252 = N1329 | N1251;
  assign N1253 = preissue_pkt_i[4] | N1252;
  assign N1254 = N395 | N1253;
  assign N1255 = N396 | N1254;
  assign N1256 = ~N1255;
  assign N1257 = N1245 | N1256;
  assign N1264 = N1631 | N525;
  assign N1265 = preissue_pkt_i[15] | N1264;
  assign N1266 = N2305 | N1265;
  assign N1267 = preissue_pkt_i[8] | N1266;
  assign N1268 = preissue_pkt_i[7] | N1267;
  assign N1269 = N394 | N1268;
  assign N1270 = preissue_pkt_i[5] | N1269;
  assign N1271 = preissue_pkt_i[4] | N1270;
  assign N1272 = N395 | N1271;
  assign N1273 = N396 | N1272;
  assign N1274 = ~N1273;
  assign N1275 = N1329 | N1269;
  assign N1276 = preissue_pkt_i[4] | N1275;
  assign N1277 = N395 | N1276;
  assign N1278 = N396 | N1277;
  assign N1279 = ~N1278;
  assign N1280 = N1274 | N1279;
  assign N1281 = preissue_pkt_i[5] | N1298;
  assign N1282 = preissue_pkt_i[4] | N1281;
  assign N1283 = N395 | N1282;
  assign N1284 = N396 | N1283;
  assign N1285 = ~N1284;
  assign N1286 = N1280 | N1285;
  assign N1287 = ~preissue_pkt_i[32];
  assign N1288 = N1287 | preissue_pkt_i[33];
  assign N1289 = preissue_pkt_i[31] | N1288;
  assign N1290 = preissue_pkt_i[30] | N1289;
  assign N1291 = preissue_pkt_i[29] | N1290;
  assign N1292 = preissue_pkt_i[28] | N1291;
  assign N1293 = N1631 | N1292;
  assign N1294 = preissue_pkt_i[15] | N1293;
  assign N1295 = N2305 | N1294;
  assign N1296 = preissue_pkt_i[8] | N1295;
  assign N1297 = preissue_pkt_i[7] | N1296;
  assign N1298 = N394 | N1297;
  assign N1299 = N1329 | N1298;
  assign N1300 = preissue_pkt_i[4] | N1299;
  assign N1301 = N395 | N1300;
  assign N1302 = N396 | N1301;
  assign N1303 = ~N1302;
  assign N1304 = N1286 | N1303;
  assign N1311 = N394 | N1389;
  assign N1312 = preissue_pkt_i[5] | N1311;
  assign N1313 = preissue_pkt_i[4] | N1312;
  assign N1314 = N395 | N1313;
  assign N1315 = N396 | N1314;
  assign N1316 = ~N1315;
  assign N1317 = N2305 | N1386;
  assign N1318 = preissue_pkt_i[8] | N1317;
  assign N1319 = preissue_pkt_i[7] | N1318;
  assign N1320 = N394 | N1319;
  assign N1321 = preissue_pkt_i[5] | N1320;
  assign N1322 = preissue_pkt_i[4] | N1321;
  assign N1323 = N395 | N1322;
  assign N1324 = N396 | N1323;
  assign N1325 = ~N1324;
  assign N1326 = N1316 | N1325;
  assign N1327 = ~preissue_pkt_i[8];
  assign N1328 = ~preissue_pkt_i[7];
  assign N1329 = ~preissue_pkt_i[5];
  assign N1330 = ~preissue_pkt_i[4];
  assign N1331 = N1328 | N1327;
  assign N1332 = preissue_pkt_i[6] | N1331;
  assign N1333 = N1329 | N1332;
  assign N1334 = N1330 | N1333;
  assign N1335 = N395 | N1334;
  assign N1336 = N396 | N1335;
  assign N1337 = ~N1336;
  assign N1338 = preissue_pkt_i[15] | preissue_pkt_i[16];
  assign N1339 = preissue_pkt_i[14] | N1338;
  assign N1340 = N1327 | N1339;
  assign N1341 = N1328 | N1340;
  assign N1342 = preissue_pkt_i[6] | N1341;
  assign N1343 = preissue_pkt_i[5] | N1342;
  assign N1344 = N1330 | N1343;
  assign N1345 = N395 | N1344;
  assign N1346 = N396 | N1345;
  assign N1347 = ~N1346;
  assign N1348 = N1337 | N1347;
  assign N1350 = preissue_pkt_i[4] | N395;
  assign N1351 = N1350 | N396;
  assign N1352 = N2553 | N1351;
  assign N1354 = N1631 & N2304;
  assign N1355 = N1354 & N2305;
  assign N1356 = N1354 & preissue_pkt_i[14];
  assign N1357 = preissue_pkt_i[16] & N2304;
  assign N1358 = N1357 & N2305;
  assign N1359 = N1357 & preissue_pkt_i[14];
  assign N1360 = preissue_pkt_i[16] & preissue_pkt_i[15];
  assign N1361 = N1360 & N2305;
  assign N1362 = N1360 & preissue_pkt_i[14];
  assign N1363 = N1631 & preissue_pkt_i[15];
  assign N1374 = N2568 | N1351;
  assign N1376 = N1363 & N2305;
  assign N1377 = N1363 & preissue_pkt_i[14];
  assign N1386 = N2304 | preissue_pkt_i[16];
  assign N1387 = preissue_pkt_i[14] | N1386;
  assign N1388 = preissue_pkt_i[8] | N1387;
  assign N1389 = preissue_pkt_i[7] | N1388;
  assign N1390 = preissue_pkt_i[6] | N1389;
  assign N1391 = preissue_pkt_i[5] | N1390;
  assign N1392 = N1330 | N1391;
  assign N1393 = N395 | N1392;
  assign N1394 = N396 | N1393;
  assign N1395 = ~N1394;
  assign N1396 = preissue_pkt_i[4] & preissue_pkt_i[3];
  assign N1397 = N1363 & N1426;
  assign N1398 = N2561 & N1396;
  assign N1399 = N1397 & N1398;
  assign N1400 = N1399 & preissue_pkt_i[2];
  assign N1404 = N1631 & N1327;
  assign N1405 = preissue_pkt_i[7] & N394;
  assign N1406 = N1404 & N1405;
  assign N1407 = N2290 & N173;
  assign N1408 = N1406 & N1407;
  assign N1410 = N2304 & N2305;
  assign N1411 = N2304 & preissue_pkt_i[14];
  assign N1412 = preissue_pkt_i[15] & N2305;
  assign N1413 = preissue_pkt_i[15] & preissue_pkt_i[14];
  assign N1419 = N1327 & preissue_pkt_i[7];
  assign N1420 = N1363 & N1419;
  assign N1421 = N1420 & N1398;
  assign N1422 = N1421 & preissue_pkt_i[2];
  assign N1426 = N1327 & N1328;
  assign N1427 = N1426 & N173;
  assign N1429 = N2305 & N394;
  assign N1430 = N1354 & N1429;
  assign N1431 = N1430 & N2295;
  assign N1432 = preissue_pkt_i[14] & N394;
  assign N1433 = N1354 & N1432;
  assign N1434 = N1433 & N2295;
  assign N1435 = N1075 & N1442;
  assign N1436 = N1449 & N1435;
  assign N1437 = N1436 & N1467;
  assign N1438 = N1068 & N1442;
  assign N1439 = N1449 & N1438;
  assign N1440 = N1439 & N1467;
  assign N1441 = preissue_pkt_i[14] & N1589;
  assign N1442 = N1360 & N1441;
  assign N1443 = N1461 & N1442;
  assign N1444 = N1449 & N1443;
  assign N1445 = N1444 & N1467;
  assign N1446 = N1003 & N1462;
  assign N1447 = N1449 & N1446;
  assign N1448 = N1447 & N1467;
  assign N1449 = N1976 & N1014;
  assign N1450 = N1068 & N1462;
  assign N1451 = N1449 & N1450;
  assign N1452 = N1451 & N1467;
  assign N1453 = N1075 & N1462;
  assign N1454 = N1465 & N1453;
  assign N1455 = N1454 & N1467;
  assign N1456 = preissue_pkt_i[23] & N2035;
  assign N1457 = N2305 & N1589;
  assign N1458 = N1590 & N1591;
  assign N1459 = N1592 & N1593;
  assign N1460 = N2666 & N1010;
  assign N1461 = N2383 & N1456;
  assign N1462 = N1363 & N1457;
  assign N1463 = N1458 & N1459;
  assign N1464 = N2575 & preissue_pkt_i[4];
  assign N1465 = N1976 & N1460;
  assign N1466 = N1461 & N1462;
  assign N1467 = N1463 & N1464;
  assign N1468 = N1465 & N1466;
  assign N1469 = N1468 & N1467;
  assign N1470 = N2035 & preissue_pkt_i[16];
  assign N1471 = N1470 & N1412;
  assign N1472 = N1474 & N1471;
  assign N1473 = N1472 & N1484;
  assign N1474 = N1880 & N1881;
  assign N1475 = N1474 & N1480;
  assign N1476 = N1475 & N1484;
  assign N1477 = preissue_pkt_i[22] & preissue_pkt_i[16];
  assign N1478 = N1593 & preissue_pkt_i[6];
  assign N1479 = N1880 & N1886;
  assign N1480 = N1477 & N1412;
  assign N1481 = N1594 & N1595;
  assign N1482 = N1478 & N2290;
  assign N1483 = N1479 & N1480;
  assign N1484 = N1481 & N1482;
  assign N1485 = N1483 & N1484;
  assign N1516 = N2548 | N2542;
  assign N1517 = N1516 | N1351;
  assign N1524 = N1519 & N1520;
  assign N1525 = N1521 & N1522;
  assign N1526 = N1523 & N1631;
  assign N1527 = N1524 & N1525;
  assign N1528 = N1526 & N1410;
  assign N1529 = N1075 & N1527;
  assign N1530 = N1528 & N1481;
  assign N1531 = N1465 & N1529;
  assign N1532 = N1530 & N1593;
  assign N1533 = N1531 & N1532;
  assign N1534 = preissue_pkt_i[31] | preissue_pkt_i[30];
  assign N1535 = N1564 | N1534;
  assign N1536 = N1557 | N1569;
  assign N1537 = N1535 | N1577;
  assign N1538 = N1536 | N1579;
  assign N1539 = N1537 | N1538;
  assign N1540 = N1539 | N1586;
  assign N1542 = preissue_pkt_i[33] | N1287;
  assign N1543 = N393 | preissue_pkt_i[28];
  assign N1544 = N523 | N2685;
  assign N1545 = N1542 | N1551;
  assign N1546 = N1543 | N1544;
  assign N1547 = N1545 | N1546;
  assign N1548 = N1547 | N1560;
  assign N1549 = N1548 | N1586;
  assign N1551 = N462 | N2303;
  assign N1552 = N1564 | N1551;
  assign N1553 = N1552 | N1577;
  assign N1554 = N1553 | N1560;
  assign N1555 = N1554 | N1586;
  assign N1557 = preissue_pkt_i[25] | preissue_pkt_i[24];
  assign N1558 = N2079 | preissue_pkt_i[22];
  assign N1559 = N1557 | N1558;
  assign N1560 = N1559 | N1579;
  assign N1561 = N1582 | N1560;
  assign N1562 = N1561 | N1586;
  assign N1564 = preissue_pkt_i[33] | preissue_pkt_i[32];
  assign N1565 = preissue_pkt_i[31] | N2303;
  assign N1566 = preissue_pkt_i[29] | preissue_pkt_i[28];
  assign N1567 = preissue_pkt_i[27] | preissue_pkt_i[26];
  assign N1568 = preissue_pkt_i[25] | N1183;
  assign N1569 = preissue_pkt_i[23] | N2035;
  assign N1570 = preissue_pkt_i[21] | preissue_pkt_i[20];
  assign N1571 = preissue_pkt_i[19] | preissue_pkt_i[18];
  assign N1572 = preissue_pkt_i[17] | preissue_pkt_i[16];
  assign N1573 = preissue_pkt_i[15] | preissue_pkt_i[14];
  assign N1574 = preissue_pkt_i[13] | preissue_pkt_i[12];
  assign N1575 = preissue_pkt_i[11] | preissue_pkt_i[10];
  assign N1576 = N1564 | N1565;
  assign N1577 = N1566 | N1567;
  assign N1578 = N1568 | N1569;
  assign N1579 = N1570 | N1571;
  assign N1580 = N1572 | N1573;
  assign N1581 = N1574 | N1575;
  assign N1582 = N1576 | N1577;
  assign N1583 = N1578 | N1579;
  assign N1584 = N1580 | N1581;
  assign N1585 = N1582 | N1583;
  assign N1586 = N1584 | preissue_pkt_i[9];
  assign N1587 = N1585 | N1586;
  assign N1594 = N1589 & N1590;
  assign N1595 = N1591 & N1592;
  assign N1596 = N1973 & N1986;
  assign N1597 = N2666 & N670;
  assign N1598 = N1410 & N1594;
  assign N1599 = N1595 & N1593;
  assign N1600 = N1596 & N1597;
  assign N1601 = N1598 & N1599;
  assign N1602 = N1600 & N1601;
  assign N1622 = N2305 | N1338;
  assign N1623 = N1327 | N1622;
  assign N1624 = N1328 | N1623;
  assign N1625 = N394 | N1624;
  assign N1626 = preissue_pkt_i[5] | N1625;
  assign N1627 = preissue_pkt_i[4] | N1626;
  assign N1628 = N395 | N1627;
  assign N1629 = N396 | N1628;
  assign N1630 = ~N1629;
  assign N1631 = ~preissue_pkt_i[16];
  assign N1632 = preissue_pkt_i[15] | N1631;
  assign N1633 = N2305 | N1632;
  assign N1634 = N1327 | N1633;
  assign N1635 = N1328 | N1634;
  assign N1636 = N394 | N1635;
  assign N1637 = preissue_pkt_i[5] | N1636;
  assign N1638 = preissue_pkt_i[4] | N1637;
  assign N1639 = N395 | N1638;
  assign N1640 = N396 | N1639;
  assign N1641 = ~N1640;
  assign N1642 = N1630 | N1641;
  assign N1644 = N2079 | N2035;
  assign N1645 = N1557 | N1644;
  assign N1646 = N1537 | N1645;
  assign N1647 = N1537 | N1536;
  assign N1648 = N1537 | N1559;
  assign N1650 = N1654 | N1659;
  assign N1652 = N2135 | N1287;
  assign N1653 = N1652 | N1534;
  assign N1654 = N1653 | N1577;
  assign N1655 = N1654 | N1559;
  assign N1657 = preissue_pkt_i[23] | preissue_pkt_i[22];
  assign N1658 = N1543 | N1567;
  assign N1659 = N1557 | N1657;
  assign N1660 = N1576 | N1658;
  assign N1661 = N1660 | N1659;
  assign N1706 = preissue_pkt_i[15] | N361;
  assign N1707 = preissue_pkt_i[14] | N1706;
  assign N1708 = N1327 | N1707;
  assign N1709 = preissue_pkt_i[7] | N1708;
  assign N1710 = N394 | N1709;
  assign N1711 = preissue_pkt_i[5] | N1710;
  assign N1712 = preissue_pkt_i[4] | N1711;
  assign N1713 = N395 | N1712;
  assign N1714 = N396 | N1713;
  assign N1715 = ~N1714;
  assign N1716 = N2305 | N1706;
  assign N1717 = N1327 | N1716;
  assign N1718 = preissue_pkt_i[7] | N1717;
  assign N1719 = N394 | N1718;
  assign N1720 = preissue_pkt_i[5] | N1719;
  assign N1721 = preissue_pkt_i[4] | N1720;
  assign N1722 = N395 | N1721;
  assign N1723 = N396 | N1722;
  assign N1724 = ~N1723;
  assign N1725 = N1715 | N1724;
  assign N1726 = N1327 | N363;
  assign N1727 = preissue_pkt_i[7] | N1726;
  assign N1728 = N394 | N1727;
  assign N1729 = preissue_pkt_i[5] | N1728;
  assign N1730 = preissue_pkt_i[4] | N1729;
  assign N1731 = N395 | N1730;
  assign N1732 = N396 | N1731;
  assign N1733 = ~N1732;
  assign N1734 = N1725 | N1733;
  assign N1735 = preissue_pkt_i[14] | N1749;
  assign N1736 = N1327 | N1735;
  assign N1737 = preissue_pkt_i[7] | N1736;
  assign N1738 = N394 | N1737;
  assign N1739 = preissue_pkt_i[5] | N1738;
  assign N1740 = preissue_pkt_i[4] | N1739;
  assign N1741 = N395 | N1740;
  assign N1742 = N396 | N1741;
  assign N1743 = ~N1742;
  assign N1744 = N1734 | N1743;
  assign N1745 = N393 | N971;
  assign N1746 = preissue_pkt_i[28] | N1745;
  assign N1747 = preissue_pkt_i[27] | N1746;
  assign N1748 = preissue_pkt_i[16] | N1747;
  assign N1749 = preissue_pkt_i[15] | N1748;
  assign N1750 = N2305 | N1749;
  assign N1751 = N1327 | N1750;
  assign N1752 = preissue_pkt_i[7] | N1751;
  assign N1753 = N394 | N1752;
  assign N1754 = preissue_pkt_i[5] | N1753;
  assign N1755 = preissue_pkt_i[4] | N1754;
  assign N1756 = N395 | N1755;
  assign N1757 = N396 | N1756;
  assign N1758 = ~N1757;
  assign N1759 = N1744 | N1758;
  assign N1760 = N2304 | N1787;
  assign N1761 = preissue_pkt_i[14] | N1760;
  assign N1762 = N1327 | N1761;
  assign N1763 = preissue_pkt_i[7] | N1762;
  assign N1764 = N394 | N1763;
  assign N1765 = preissue_pkt_i[5] | N1764;
  assign N1766 = preissue_pkt_i[4] | N1765;
  assign N1767 = N395 | N1766;
  assign N1768 = N396 | N1767;
  assign N1769 = ~N1768;
  assign N1770 = N1759 | N1769;
  assign N1771 = N2305 | N1788;
  assign N1772 = N1327 | N1771;
  assign N1773 = preissue_pkt_i[7] | N1772;
  assign N1774 = N394 | N1773;
  assign N1775 = preissue_pkt_i[5] | N1774;
  assign N1776 = preissue_pkt_i[4] | N1775;
  assign N1777 = N395 | N1776;
  assign N1778 = N396 | N1777;
  assign N1779 = ~N1778;
  assign N1780 = N1770 | N1779;
  assign N1781 = preissue_pkt_i[32] | N2135;
  assign N1782 = N462 | N1781;
  assign N1783 = preissue_pkt_i[30] | N1782;
  assign N1784 = preissue_pkt_i[29] | N1783;
  assign N1785 = preissue_pkt_i[28] | N1784;
  assign N1786 = preissue_pkt_i[27] | N1785;
  assign N1787 = preissue_pkt_i[16] | N1786;
  assign N1788 = preissue_pkt_i[15] | N1787;
  assign N1789 = preissue_pkt_i[14] | N1788;
  assign N1790 = N1327 | N1789;
  assign N1791 = preissue_pkt_i[7] | N1790;
  assign N1792 = N394 | N1791;
  assign N1793 = preissue_pkt_i[5] | N1792;
  assign N1794 = preissue_pkt_i[4] | N1793;
  assign N1795 = N395 | N1794;
  assign N1796 = N396 | N1795;
  assign N1797 = ~N1796;
  assign N1798 = N1780 | N1797;
  assign N1799 = N2305 | N2220;
  assign N1800 = N1327 | N1799;
  assign N1801 = preissue_pkt_i[7] | N1800;
  assign N1802 = N394 | N1801;
  assign N1803 = preissue_pkt_i[5] | N1802;
  assign N1804 = preissue_pkt_i[4] | N1803;
  assign N1805 = N395 | N1804;
  assign N1806 = N396 | N1805;
  assign N1807 = ~N1806;
  assign N1808 = N1798 | N1807;
  assign N1809 = preissue_pkt_i[27] | N525;
  assign N1810 = N1327 | N1809;
  assign N1811 = preissue_pkt_i[7] | N1810;
  assign N1812 = N394 | N1811;
  assign N1813 = preissue_pkt_i[5] | N1812;
  assign N1814 = preissue_pkt_i[4] | N1813;
  assign N1815 = N395 | N1814;
  assign N1816 = N396 | N1815;
  assign N1817 = ~N1816;
  assign N1818 = N1808 | N1817;
  assign N1819 = N1327 | N402;
  assign N1820 = preissue_pkt_i[7] | N1819;
  assign N1821 = N394 | N1820;
  assign N1822 = preissue_pkt_i[5] | N1821;
  assign N1823 = preissue_pkt_i[4] | N1822;
  assign N1824 = N395 | N1823;
  assign N1825 = N396 | N1824;
  assign N1826 = ~N1825;
  assign N1827 = N1818 | N1826;
  assign N1828 = preissue_pkt_i[28] | N2307;
  assign N1829 = preissue_pkt_i[27] | N1828;
  assign N1830 = N1327 | N1829;
  assign N1831 = preissue_pkt_i[7] | N1830;
  assign N1832 = N394 | N1831;
  assign N1833 = preissue_pkt_i[5] | N1832;
  assign N1834 = preissue_pkt_i[4] | N1833;
  assign N1835 = N395 | N1834;
  assign N1836 = N396 | N1835;
  assign N1837 = ~N1836;
  assign N1838 = N1827 | N1837;
  assign N1839 = N393 | N2306;
  assign N1840 = preissue_pkt_i[28] | N1839;
  assign N1841 = preissue_pkt_i[27] | N1840;
  assign N1842 = N1327 | N1841;
  assign N1843 = preissue_pkt_i[7] | N1842;
  assign N1844 = N394 | N1843;
  assign N1845 = preissue_pkt_i[5] | N1844;
  assign N1846 = preissue_pkt_i[4] | N1845;
  assign N1847 = N395 | N1846;
  assign N1848 = N396 | N1847;
  assign N1849 = ~N1848;
  assign N1850 = N1838 | N1849;
  assign N1851 = N2303 | N1289;
  assign N1852 = N393 | N1851;
  assign N1853 = preissue_pkt_i[28] | N1852;
  assign N1854 = preissue_pkt_i[27] | N1853;
  assign N1855 = preissue_pkt_i[26] | N1854;
  assign N1856 = preissue_pkt_i[25] | N1855;
  assign N1857 = preissue_pkt_i[24] | N1856;
  assign N1858 = preissue_pkt_i[23] | N1857;
  assign N1859 = preissue_pkt_i[22] | N1858;
  assign N1860 = N1327 | N1859;
  assign N1861 = preissue_pkt_i[7] | N1860;
  assign N1862 = N394 | N1861;
  assign N1863 = preissue_pkt_i[5] | N1862;
  assign N1864 = preissue_pkt_i[4] | N1863;
  assign N1865 = N395 | N1864;
  assign N1866 = N396 | N1865;
  assign N1867 = ~N1866;
  assign N1868 = N1850 | N1867;
  assign N1869 = N2684 & preissue_pkt_i[8];
  assign N1870 = N1328 & preissue_pkt_i[6];
  assign N1871 = N1869 & N1870;
  assign N1872 = N1871 & N1407;
  assign N1874 = N1007 & N1974;
  assign N1875 = N1874 & N1882;
  assign N1876 = N1875 & N1894;
  assign N1877 = N1874 & N1889;
  assign N1878 = N1877 & N1883;
  assign N1880 = N2685 & N2686;
  assign N1881 = N1183 & N2079;
  assign N1882 = N1975 & N1880;
  assign N1883 = N1881 & N2035;
  assign N1884 = N2446 & N1882;
  assign N1885 = N1884 & N1883;
  assign N1886 = N1183 & preissue_pkt_i[23];
  assign N1887 = N1886 & N2035;
  assign N1888 = N1884 & N1887;
  assign N1889 = N1978 & N1880;
  assign N1890 = N2446 & N1889;
  assign N1891 = N1890 & N1883;
  assign N1892 = N1890 & N1887;
  assign N1894 = N1881 & preissue_pkt_i[22];
  assign N1895 = N1884 & N1894;
  assign N1896 = N1886 & preissue_pkt_i[22];
  assign N1897 = N1884 & N1896;
  assign N1898 = N1890 & N1894;
  assign N1899 = N1890 & N1896;
  assign N1901 = N2445 & N1986;
  assign N1902 = N1901 & N1882;
  assign N1903 = N1902 & N1883;
  assign N1904 = N1902 & N1887;
  assign N1905 = N1901 & N1889;
  assign N1906 = N1905 & N1883;
  assign N1907 = N1905 & N1887;
  assign N1909 = N1902 & N1894;
  assign N1910 = N1902 & N1896;
  assign N1911 = N1905 & N1894;
  assign N1912 = N1905 & N1896;
  assign N1914 = N2035 & N1631;
  assign N1915 = N1881 & N1914;
  assign N1916 = N2451 & N1882;
  assign N1917 = N1915 & N1410;
  assign N1918 = N1916 & N1917;
  assign N1919 = N2451 & N1889;
  assign N1920 = N1919 & N1917;
  assign N1922 = N2445 & N2457;
  assign N1923 = N1922 & N1882;
  assign N1924 = N1923 & N1917;
  assign N1925 = N1922 & N1889;
  assign N1926 = N1925 & N1917;
  assign N1928 = N1973 & N2005;
  assign N1929 = N1975 & N1354;
  assign N1930 = N1928 & N1929;
  assign N1931 = N1930 & N2305;
  assign N1932 = N1978 & N1354;
  assign N1933 = N1928 & N1932;
  assign N1934 = N1933 & N2305;
  assign N1936 = N1930 & preissue_pkt_i[14];
  assign N1937 = N1933 & preissue_pkt_i[14];
  assign N1939 = N1975 & N1363;
  assign N1940 = N1928 & N1939;
  assign N1941 = N1940 & N2305;
  assign N1942 = N1978 & N1363;
  assign N1943 = N1928 & N1942;
  assign N1944 = N1943 & N2305;
  assign N1946 = N616 & N1354;
  assign N1947 = N1928 & N1946;
  assign N1948 = N1947 & N2305;
  assign N1949 = N591 & N1354;
  assign N1950 = N1928 & N1949;
  assign N1951 = N1950 & N2305;
  assign N1953 = N1947 & preissue_pkt_i[14];
  assign N1954 = N1950 & preissue_pkt_i[14];
  assign N1956 = N2440 & N1939;
  assign N1957 = N1956 & N2305;
  assign N1958 = N2440 & N1942;
  assign N1959 = N1958 & N2305;
  assign N1961 = N2440 & N1929;
  assign N1962 = N1961 & preissue_pkt_i[14];
  assign N1963 = N2440 & N1932;
  assign N1964 = N1963 & preissue_pkt_i[14];
  assign N1966 = N1961 & N2305;
  assign N1967 = N1963 & N2305;
  assign N1969 = N1915 & N1411;
  assign N1970 = N1916 & N1969;
  assign N1971 = N1919 & N1969;
  assign N1973 = N2135 & N1287;
  assign N1974 = N462 & N2303;
  assign N1975 = N393 & N523;
  assign N1976 = N1973 & N1974;
  assign N1977 = N1976 & N1975;
  assign N1978 = N393 & preissue_pkt_i[27];
  assign N1979 = N1976 & N1978;
  assign N1981 = N1976 & N616;
  assign N1982 = N2135 & N1287;
  assign N1983 = N1982 & N1974;
  assign N1984 = N1983 & N591;
  assign N1986 = N462 & preissue_pkt_i[30];
  assign N1987 = N1982 & N1986;
  assign N1988 = N1987 & N1975;
  assign N1989 = N1987 & N1978;
  assign N1991 = N1987 & N616;
  assign N1992 = N1987 & N591;
  assign N1994 = N2002 & N1986;
  assign N1995 = N616 & N1880;
  assign N1996 = N1994 & N1995;
  assign N1997 = N1996 & N1883;
  assign N1998 = N591 & N1880;
  assign N1999 = N1994 & N1998;
  assign N2000 = N1999 & N1883;
  assign N2002 = N2135 & preissue_pkt_i[32];
  assign N2003 = preissue_pkt_i[27] & preissue_pkt_i[22];
  assign N2004 = N2002 & N2003;
  assign N2005 = preissue_pkt_i[31] & N2303;
  assign N2006 = N2002 & N2005;
  assign N2007 = N2006 & preissue_pkt_i[27];
  assign N2008 = preissue_pkt_i[32] & preissue_pkt_i[26];
  assign N2009 = preissue_pkt_i[32] & preissue_pkt_i[25];
  assign N2010 = preissue_pkt_i[32] & preissue_pkt_i[24];
  assign N2011 = preissue_pkt_i[30] & preissue_pkt_i[22];
  assign N2012 = N2002 & N2011;
  assign N2013 = N2460 & preissue_pkt_i[22];
  assign N2014 = N2460 & preissue_pkt_i[23];
  assign N2015 = N622 & preissue_pkt_i[29];
  assign N2016 = N2002 & N2463;
  assign N2017 = N2457 & preissue_pkt_i[14];
  assign N2018 = preissue_pkt_i[32] & N2303;
  assign N2019 = N2018 & preissue_pkt_i[29];
  assign N2020 = N622 & preissue_pkt_i[22];
  assign N2021 = N2002 & preissue_pkt_i[23];
  assign N2022 = N2303 & N523;
  assign N2023 = N2002 & N2022;
  assign N2024 = N2023 & N2035;
  assign N2025 = N622 & preissue_pkt_i[23];
  assign N2026 = N2458 & preissue_pkt_i[15];
  assign N2027 = preissue_pkt_i[33] & N1287;
  assign N2028 = N2027 & N462;
  assign N2029 = N2027 & preissue_pkt_i[30];
  assign N2030 = N2027 & preissue_pkt_i[16];
  assign N2031 = N2027 & N1413;
  assign N2032 = N659 & preissue_pkt_i[30];
  assign N2033 = preissue_pkt_i[31] & preissue_pkt_i[16];
  assign N2035 = ~preissue_pkt_i[22];
  assign N2036 = preissue_pkt_i[27] | N1292;
  assign N2037 = preissue_pkt_i[26] | N2036;
  assign N2038 = preissue_pkt_i[25] | N2037;
  assign N2039 = preissue_pkt_i[24] | N2038;
  assign N2040 = preissue_pkt_i[23] | N2039;
  assign N2041 = N2035 | N2040;
  assign N2042 = N1327 | N2041;
  assign N2043 = preissue_pkt_i[7] | N2042;
  assign N2044 = N394 | N2043;
  assign N2045 = preissue_pkt_i[5] | N2044;
  assign N2046 = preissue_pkt_i[4] | N2045;
  assign N2047 = N395 | N2046;
  assign N2048 = N396 | N2047;
  assign N2049 = N523 | N1292;
  assign N2050 = preissue_pkt_i[26] | N2049;
  assign N2051 = preissue_pkt_i[25] | N2050;
  assign N2052 = preissue_pkt_i[24] | N2051;
  assign N2053 = preissue_pkt_i[23] | N2052;
  assign N2054 = preissue_pkt_i[22] | N2053;
  assign N2055 = N1327 | N2054;
  assign N2056 = preissue_pkt_i[7] | N2055;
  assign N2057 = N394 | N2056;
  assign N2058 = preissue_pkt_i[5] | N2057;
  assign N2059 = preissue_pkt_i[4] | N2058;
  assign N2060 = N395 | N2059;
  assign N2061 = N396 | N2060;
  assign N2062 = preissue_pkt_i[30] | N2137;
  assign N2063 = preissue_pkt_i[29] | N2062;
  assign N2064 = preissue_pkt_i[28] | N2063;
  assign N2065 = preissue_pkt_i[27] | N2064;
  assign N2066 = preissue_pkt_i[26] | N2065;
  assign N2067 = preissue_pkt_i[25] | N2066;
  assign N2068 = preissue_pkt_i[24] | N2067;
  assign N2069 = preissue_pkt_i[23] | N2068;
  assign N2070 = preissue_pkt_i[22] | N2069;
  assign N2071 = N1327 | N2070;
  assign N2072 = preissue_pkt_i[7] | N2071;
  assign N2073 = N394 | N2072;
  assign N2074 = preissue_pkt_i[5] | N2073;
  assign N2075 = preissue_pkt_i[4] | N2074;
  assign N2076 = N395 | N2075;
  assign N2077 = N396 | N2076;
  assign N2078 = ~N2077;
  assign N2079 = ~preissue_pkt_i[23];
  assign N2080 = N2079 | N2068;
  assign N2081 = preissue_pkt_i[22] | N2080;
  assign N2082 = N1327 | N2081;
  assign N2083 = preissue_pkt_i[7] | N2082;
  assign N2084 = N394 | N2083;
  assign N2085 = preissue_pkt_i[5] | N2084;
  assign N2086 = preissue_pkt_i[4] | N2085;
  assign N2087 = N395 | N2086;
  assign N2088 = N396 | N2087;
  assign N2089 = ~N2088;
  assign N2090 = N2078 | N2089;
  assign N2091 = N523 | N2064;
  assign N2092 = preissue_pkt_i[26] | N2091;
  assign N2093 = preissue_pkt_i[25] | N2092;
  assign N2094 = preissue_pkt_i[24] | N2093;
  assign N2095 = preissue_pkt_i[23] | N2094;
  assign N2096 = preissue_pkt_i[22] | N2095;
  assign N2097 = N1327 | N2096;
  assign N2098 = preissue_pkt_i[7] | N2097;
  assign N2099 = N394 | N2098;
  assign N2100 = preissue_pkt_i[5] | N2099;
  assign N2101 = preissue_pkt_i[4] | N2100;
  assign N2102 = N395 | N2101;
  assign N2103 = N396 | N2102;
  assign N2104 = ~N2103;
  assign N2105 = N2078 | N2104;
  assign N2106 = N2035 | N2069;
  assign N2107 = N1327 | N2106;
  assign N2108 = preissue_pkt_i[7] | N2107;
  assign N2109 = N394 | N2108;
  assign N2110 = preissue_pkt_i[5] | N2109;
  assign N2111 = preissue_pkt_i[4] | N2110;
  assign N2112 = N395 | N2111;
  assign N2113 = N396 | N2112;
  assign N2114 = ~N2113;
  assign N2115 = N2035 | N2080;
  assign N2116 = N1327 | N2115;
  assign N2117 = preissue_pkt_i[7] | N2116;
  assign N2118 = N394 | N2117;
  assign N2119 = preissue_pkt_i[5] | N2118;
  assign N2120 = preissue_pkt_i[4] | N2119;
  assign N2121 = N395 | N2120;
  assign N2122 = N396 | N2121;
  assign N2123 = ~N2122;
  assign N2124 = N2114 | N2123;
  assign N2125 = N2035 | N2095;
  assign N2126 = N1327 | N2125;
  assign N2127 = preissue_pkt_i[7] | N2126;
  assign N2128 = N394 | N2127;
  assign N2129 = preissue_pkt_i[5] | N2128;
  assign N2130 = preissue_pkt_i[4] | N2129;
  assign N2131 = N395 | N2130;
  assign N2132 = N396 | N2131;
  assign N2133 = ~N2132;
  assign N2134 = N2114 | N2133;
  assign N2135 = ~preissue_pkt_i[33];
  assign N2136 = N1287 | N2135;
  assign N2137 = preissue_pkt_i[31] | N2136;
  assign N2138 = N2303 | N2137;
  assign N2139 = preissue_pkt_i[29] | N2138;
  assign N2140 = preissue_pkt_i[28] | N2139;
  assign N2141 = preissue_pkt_i[27] | N2140;
  assign N2142 = preissue_pkt_i[26] | N2141;
  assign N2143 = preissue_pkt_i[25] | N2142;
  assign N2144 = preissue_pkt_i[24] | N2143;
  assign N2145 = preissue_pkt_i[23] | N2144;
  assign N2146 = preissue_pkt_i[22] | N2145;
  assign N2147 = N1327 | N2146;
  assign N2148 = preissue_pkt_i[7] | N2147;
  assign N2149 = N394 | N2148;
  assign N2150 = preissue_pkt_i[5] | N2149;
  assign N2151 = preissue_pkt_i[4] | N2150;
  assign N2152 = N395 | N2151;
  assign N2153 = N396 | N2152;
  assign N2154 = ~N2153;
  assign N2155 = N523 | N2140;
  assign N2156 = preissue_pkt_i[26] | N2155;
  assign N2157 = preissue_pkt_i[25] | N2156;
  assign N2158 = preissue_pkt_i[24] | N2157;
  assign N2159 = preissue_pkt_i[23] | N2158;
  assign N2160 = preissue_pkt_i[22] | N2159;
  assign N2161 = N1327 | N2160;
  assign N2162 = preissue_pkt_i[7] | N2161;
  assign N2163 = N394 | N2162;
  assign N2164 = preissue_pkt_i[5] | N2163;
  assign N2165 = preissue_pkt_i[4] | N2164;
  assign N2166 = N395 | N2165;
  assign N2167 = N396 | N2166;
  assign N2168 = ~N2167;
  assign N2169 = N2154 | N2168;
  assign N2170 = N2079 | N2144;
  assign N2171 = preissue_pkt_i[22] | N2170;
  assign N2172 = N1327 | N2171;
  assign N2173 = preissue_pkt_i[7] | N2172;
  assign N2174 = N394 | N2173;
  assign N2175 = preissue_pkt_i[5] | N2174;
  assign N2176 = preissue_pkt_i[4] | N2175;
  assign N2177 = N395 | N2176;
  assign N2178 = N396 | N2177;
  assign N2179 = ~N2178;
  assign N2180 = N2154 | N2179;
  assign N2181 = N2035 | N2145;
  assign N2182 = N1327 | N2181;
  assign N2183 = preissue_pkt_i[7] | N2182;
  assign N2184 = N394 | N2183;
  assign N2185 = preissue_pkt_i[5] | N2184;
  assign N2186 = preissue_pkt_i[4] | N2185;
  assign N2187 = N395 | N2186;
  assign N2188 = N396 | N2187;
  assign N2189 = ~N2188;
  assign N2190 = N2035 | N2159;
  assign N2191 = N1327 | N2190;
  assign N2192 = preissue_pkt_i[7] | N2191;
  assign N2193 = N394 | N2192;
  assign N2194 = preissue_pkt_i[5] | N2193;
  assign N2195 = preissue_pkt_i[4] | N2194;
  assign N2196 = N395 | N2195;
  assign N2197 = N396 | N2196;
  assign N2198 = ~N2197;
  assign N2199 = N2189 | N2198;
  assign N2200 = N2035 | N2170;
  assign N2201 = N1327 | N2200;
  assign N2202 = preissue_pkt_i[7] | N2201;
  assign N2203 = N394 | N2202;
  assign N2204 = preissue_pkt_i[5] | N2203;
  assign N2205 = preissue_pkt_i[4] | N2204;
  assign N2206 = N395 | N2205;
  assign N2207 = N396 | N2206;
  assign N2208 = ~N2207;
  assign N2209 = N2189 | N2208;
  assign N2210 = preissue_pkt_i[30] | N2230;
  assign N2211 = preissue_pkt_i[29] | N2210;
  assign N2212 = preissue_pkt_i[28] | N2211;
  assign N2213 = preissue_pkt_i[27] | N2212;
  assign N2214 = preissue_pkt_i[26] | N2213;
  assign N2215 = preissue_pkt_i[25] | N2214;
  assign N2216 = preissue_pkt_i[24] | N2215;
  assign N2217 = preissue_pkt_i[23] | N2216;
  assign N2218 = preissue_pkt_i[22] | N2217;
  assign N2219 = preissue_pkt_i[16] | N2218;
  assign N2220 = preissue_pkt_i[15] | N2219;
  assign N2221 = preissue_pkt_i[14] | N2220;
  assign N2222 = N1327 | N2221;
  assign N2223 = preissue_pkt_i[7] | N2222;
  assign N2224 = N394 | N2223;
  assign N2225 = preissue_pkt_i[5] | N2224;
  assign N2226 = preissue_pkt_i[4] | N2225;
  assign N2227 = N395 | N2226;
  assign N2228 = N396 | N2227;
  assign N2229 = ~N2228;
  assign N2230 = N462 | N2136;
  assign N2231 = N2303 | N2230;
  assign N2232 = preissue_pkt_i[29] | N2231;
  assign N2233 = preissue_pkt_i[28] | N2232;
  assign N2234 = preissue_pkt_i[27] | N2233;
  assign N2235 = preissue_pkt_i[26] | N2234;
  assign N2236 = preissue_pkt_i[25] | N2235;
  assign N2237 = preissue_pkt_i[24] | N2236;
  assign N2238 = preissue_pkt_i[23] | N2237;
  assign N2239 = preissue_pkt_i[22] | N2238;
  assign N2240 = preissue_pkt_i[16] | N2239;
  assign N2241 = preissue_pkt_i[15] | N2240;
  assign N2242 = preissue_pkt_i[14] | N2241;
  assign N2243 = N1327 | N2242;
  assign N2244 = preissue_pkt_i[7] | N2243;
  assign N2245 = N394 | N2244;
  assign N2246 = preissue_pkt_i[5] | N2245;
  assign N2247 = preissue_pkt_i[4] | N2246;
  assign N2248 = N395 | N2247;
  assign N2249 = N396 | N2248;
  assign N2250 = ~N2249;
  assign N2286 = N394 & preissue_pkt_i[3];
  assign N2287 = N2577 & N2286;
  assign N2288 = N2287 & preissue_pkt_i[2];
  assign N2290 = N1329 & N1330;
  assign N2291 = preissue_pkt_i[5] | N1330;
  assign N2293 = N1329 | preissue_pkt_i[4];
  assign N2295 = preissue_pkt_i[5] & preissue_pkt_i[4];
  assign N2303 = ~preissue_pkt_i[30];
  assign N2304 = ~preissue_pkt_i[15];
  assign N2305 = ~preissue_pkt_i[14];
  assign N2306 = N2303 | N398;
  assign N2307 = preissue_pkt_i[29] | N2306;
  assign N2308 = preissue_pkt_i[26] | N2307;
  assign N2309 = preissue_pkt_i[25] | N2308;
  assign N2310 = preissue_pkt_i[24] | N2309;
  assign N2311 = preissue_pkt_i[23] | N2310;
  assign N2312 = preissue_pkt_i[22] | N2311;
  assign N2313 = preissue_pkt_i[16] | N2312;
  assign N2314 = N2304 | N2313;
  assign N2315 = N2305 | N2314;
  assign N2316 = preissue_pkt_i[8] | N2315;
  assign N2317 = N1328 | N2316;
  assign N2318 = preissue_pkt_i[6] | N2317;
  assign N2319 = N1329 | N2318;
  assign N2320 = N1330 | N2319;
  assign N2321 = N395 | N2320;
  assign N2322 = N396 | N2321;
  assign N2323 = ~N2322;
  assign N2324 = preissue_pkt_i[14] | N2314;
  assign N2325 = preissue_pkt_i[8] | N2324;
  assign N2326 = N1328 | N2325;
  assign N2327 = preissue_pkt_i[6] | N2326;
  assign N2328 = N1329 | N2327;
  assign N2329 = N1330 | N2328;
  assign N2330 = N395 | N2329;
  assign N2331 = N396 | N2330;
  assign N2332 = ~N2331;
  assign N2333 = N2323 | N2332;
  assign N2335 = N2575 & N1396;
  assign N2336 = N1420 & N2335;
  assign N2337 = N2336 & preissue_pkt_i[2];
  assign N2339 = N2079 & N2035;
  assign N2340 = N2339 & preissue_pkt_i[14];
  assign N2341 = N2389 & N2340;
  assign N2342 = N2339 & N2305;
  assign N2343 = N2389 & N2342;
  assign N2344 = N1987 & N668;
  assign N2345 = preissue_pkt_i[29] & N2305;
  assign N2346 = N1987 & N2345;
  assign N2347 = N1983 & N668;
  assign N2348 = N1983 & N2345;
  assign N2349 = N393 & preissue_pkt_i[14];
  assign N2350 = N1983 & N2349;
  assign N2351 = N393 & N2305;
  assign N2352 = N1983 & N2351;
  assign N2353 = N2425 & N2349;
  assign N2354 = N2425 & N2351;
  assign N2355 = N2006 & N2349;
  assign N2356 = N2006 & N2351;
  assign N2357 = N2420 & N2349;
  assign N2358 = N2420 & N2351;
  assign N2359 = N2435 & N2349;
  assign N2360 = N2435 & N2351;
  assign N2361 = N2440 & N2349;
  assign N2362 = N2440 & N2351;
  assign N2363 = N2446 & N2349;
  assign N2364 = N2446 & N2351;
  assign N2365 = N2451 & N2349;
  assign N2366 = N2451 & N2351;
  assign N2382 = N393 & N2685;
  assign N2383 = N2686 & N1183;
  assign N2384 = preissue_pkt_i[14] & N1327;
  assign N2385 = N2382 & N2383;
  assign N2386 = N2339 & N1363;
  assign N2387 = N2384 & N1405;
  assign N2388 = N2295 & N173;
  assign N2389 = N1987 & N2385;
  assign N2390 = N2386 & N2387;
  assign N2391 = N2389 & N2390;
  assign N2392 = N2391 & N2388;
  assign N2393 = N2305 & N1327;
  assign N2394 = N2393 & N1405;
  assign N2395 = N2386 & N2394;
  assign N2396 = N2389 & N2395;
  assign N2397 = N2396 & N2388;
  assign N2398 = N688 & N1413;
  assign N2399 = N1419 & N2575;
  assign N2400 = N1396 & preissue_pkt_i[2];
  assign N2401 = N1987 & N2398;
  assign N2402 = N2399 & N2400;
  assign N2403 = N2401 & N2402;
  assign N2404 = N688 & N1412;
  assign N2405 = N1987 & N2404;
  assign N2406 = N2405 & N2402;
  assign N2408 = N1983 & N2398;
  assign N2409 = N2408 & N2402;
  assign N2410 = N1983 & N2404;
  assign N2411 = N2410 & N2402;
  assign N2413 = N393 & N1631;
  assign N2414 = N2413 & N1413;
  assign N2415 = N2006 & N2414;
  assign N2416 = N2415 & N2402;
  assign N2417 = N2413 & N1412;
  assign N2418 = N2006 & N2417;
  assign N2419 = N2418 & N2402;
  assign N2420 = N2002 & N1974;
  assign N2421 = N2420 & N2414;
  assign N2422 = N2421 & N2402;
  assign N2423 = N2420 & N2417;
  assign N2424 = N2423 & N2402;
  assign N2425 = N1982 & N2005;
  assign N2426 = N2425 & N2414;
  assign N2427 = N2426 & N2402;
  assign N2428 = N2425 & N2417;
  assign N2429 = N2428 & N2402;
  assign N2431 = N1983 & N2414;
  assign N2432 = N2431 & N2402;
  assign N2433 = N1983 & N2417;
  assign N2434 = N2433 & N2402;
  assign N2435 = N2027 & N1974;
  assign N2436 = N2435 & N2414;
  assign N2437 = N2436 & N2402;
  assign N2438 = N2435 & N2417;
  assign N2439 = N2438 & N2402;
  assign N2440 = N2027 & N2005;
  assign N2441 = N2440 & N2414;
  assign N2442 = N2441 & N2402;
  assign N2443 = N2440 & N2417;
  assign N2444 = N2443 & N2402;
  assign N2445 = preissue_pkt_i[33] & preissue_pkt_i[32];
  assign N2446 = N2445 & N1974;
  assign N2447 = N2446 & N2414;
  assign N2448 = N2447 & N2402;
  assign N2449 = N2446 & N2417;
  assign N2450 = N2449 & N2402;
  assign N2451 = N2445 & N2005;
  assign N2452 = N2451 & N2414;
  assign N2453 = N2452 & N2402;
  assign N2454 = N2451 & N2417;
  assign N2455 = N2454 & N2402;
  assign N2457 = preissue_pkt_i[31] & preissue_pkt_i[30];
  assign N2458 = preissue_pkt_i[31] & preissue_pkt_i[29];
  assign N2459 = preissue_pkt_i[33] & preissue_pkt_i[29];
  assign N2460 = preissue_pkt_i[32] & preissue_pkt_i[29];
  assign N2461 = preissue_pkt_i[32] & preissue_pkt_i[30];
  assign N2462 = preissue_pkt_i[33] & preissue_pkt_i[30];
  assign N2463 = preissue_pkt_i[30] & N393;
  assign N2464 = N2463 & preissue_pkt_i[26];
  assign N2465 = N2463 & preissue_pkt_i[25];
  assign N2466 = N2463 & preissue_pkt_i[24];
  assign N2467 = N2463 & preissue_pkt_i[23];
  assign N2468 = N2463 & preissue_pkt_i[22];
  assign N2541 = preissue_pkt_i[8] | N1328;
  assign N2542 = N394 | preissue_pkt_i[5];
  assign N2543 = N2541 | N2542;
  assign N2544 = N2543 | N1330;
  assign N2545 = N179 | N2542;
  assign N2546 = N2545 | N1330;
  assign N2548 = N1327 | N1328;
  assign N2549 = preissue_pkt_i[6] | N1329;
  assign N2550 = N2548 | N2549;
  assign N2551 = N2550 | N1330;
  assign N2553 = N2548 | N212;
  assign N2554 = N2553 | preissue_pkt_i[4];
  assign N2556 = N2541 | N212;
  assign N2557 = N2556 | preissue_pkt_i[4];
  assign N2558 = N2556 | N1330;
  assign N2560 = N2553 | N1330;
  assign N2561 = N394 & N1329;
  assign N2562 = N1426 & N2561;
  assign N2563 = N2562 & N1330;
  assign N2564 = N2545 | preissue_pkt_i[4];
  assign N2565 = N394 | N1329;
  assign N2566 = N179 | N2565;
  assign N2567 = N2566 | preissue_pkt_i[4];
  assign N2568 = N179 | N212;
  assign N2569 = N2568 | N1330;
  assign N2571 = N1327 & preissue_pkt_i[5];
  assign N2572 = N2571 & preissue_pkt_i[4];
  assign N2573 = preissue_pkt_i[7] & preissue_pkt_i[6];
  assign N2574 = N2573 & N1330;
  assign N2575 = N394 & preissue_pkt_i[5];
  assign N2576 = N2575 & N1330;
  assign N2577 = preissue_pkt_i[8] & N1328;
  assign N2643 = N1363 & N2393;
  assign N2644 = N2643 & N1017;
  assign N2645 = N2644 & N173;
  assign N2646 = N1363 & N2384;
  assign N2647 = N2646 & N1017;
  assign N2648 = N2647 & N173;
  assign N2650 = N523 & N1631;
  assign N2651 = N2666 & N2650;
  assign N2652 = N2425 & N2651;
  assign N2653 = N2652 & N2672;
  assign N2654 = N2653 & preissue_pkt_i[2];
  assign N2655 = N2652 & N2676;
  assign N2656 = N2655 & preissue_pkt_i[2];
  assign N2658 = N1410 & N1419;
  assign N2659 = N2658 & N2670;
  assign N2660 = N2671 & N2659;
  assign N2661 = N2660 & preissue_pkt_i[2];
  assign N2662 = N2658 & N2675;
  assign N2663 = N2671 & N2662;
  assign N2664 = N2663 & preissue_pkt_i[2];
  assign N2666 = N393 & N2684;
  assign N2667 = preissue_pkt_i[6] & N1329;
  assign N2668 = N2666 & N654;
  assign N2669 = N1412 & N1419;
  assign N2670 = N2667 & N541;
  assign N2671 = N2425 & N2668;
  assign N2672 = N2669 & N2670;
  assign N2673 = N2671 & N2672;
  assign N2674 = N2673 & preissue_pkt_i[2];
  assign N2675 = N239 & N541;
  assign N2676 = N2669 & N2675;
  assign N2677 = N2671 & N2676;
  assign N2678 = N2677 & preissue_pkt_i[2];
  assign N2704 = preissue_pkt_i[12] | preissue_pkt_i[13];
  assign N2705 = preissue_pkt_i[11] | N2704;
  assign N2706 = preissue_pkt_i[10] | N2705;
  assign N2707 = preissue_pkt_i[9] | N2706;
  assign N2708 = preissue_pkt_i[27] | preissue_pkt_i[28];
  assign N2709 = ~N2708;
  assign N2710 = N1328 | preissue_pkt_i[8];
  assign N2711 = N394 | N2710;
  assign N2712 = N1329 | N2711;
  assign N2713 = preissue_pkt_i[4] | N2712;
  assign N2714 = N395 | N2713;
  assign N2715 = N396 | N2714;
  assign N2716 = ~N2715;
  assign N2717 = preissue_pkt_i[7] | preissue_pkt_i[8];
  assign N2718 = N394 | N2717;
  assign N2719 = N1329 | N2718;
  assign N2720 = preissue_pkt_i[4] | N2719;
  assign N2721 = N395 | N2720;
  assign N2722 = N396 | N2721;
  assign N2723 = ~N2722;
  assign N2724 = preissue_pkt_i[20] | preissue_pkt_i[21];
  assign N2725 = preissue_pkt_i[19] | N2724;
  assign N2726 = preissue_pkt_i[18] | N2725;
  assign N2727 = preissue_pkt_i[17] | N2726;
  assign N349 = ~N348;
  assign N391 = ~N390;
  assign N392 = (N0)? N391 : 
                (N1)? 1'b0 : 1'b0;
  assign N0 = N2716;
  assign N1 = N2715;
  assign N414 = (N2)? 1'b0 : 
                (N3)? N2716 : 1'b0;
  assign N2 = N413;
  assign N3 = N412;
  assign { N714, N713, N712, N711, N710 } = (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                            (N5)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                            (N6)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                            (N7)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                                            (N8)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                            (N9)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                                            (N10)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                                            (N11)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                            (N12)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                            (N13)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                            (N14)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                            (N15)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                            (N16)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                            (N17)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                            (N18)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                            (N19)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                            (N20)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                            (N21)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                            (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                            (N23)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                            (N24)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                            (N25)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                            (N26)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N4 = N580;
  assign N5 = N587;
  assign N6 = N590;
  assign N7 = N594;
  assign N8 = N596;
  assign N9 = N598;
  assign N10 = N600;
  assign N11 = N603;
  assign N12 = N611;
  assign N13 = N614;
  assign N14 = N620;
  assign N15 = N621;
  assign N16 = N624;
  assign N17 = N627;
  assign N18 = N630;
  assign N19 = N634;
  assign N20 = N635;
  assign N21 = N636;
  assign N22 = N639;
  assign N23 = N642;
  assign N24 = N645;
  assign N25 = N649;
  assign N26 = N709;
  assign N715 = (N4)? 1'b0 : 
                (N5)? 1'b0 : 
                (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N8)? 1'b0 : 
                (N9)? 1'b0 : 
                (N10)? 1'b0 : 
                (N11)? 1'b0 : 
                (N12)? 1'b0 : 
                (N13)? 1'b0 : 
                (N14)? 1'b0 : 
                (N15)? 1'b0 : 
                (N16)? 1'b0 : 
                (N17)? 1'b0 : 
                (N18)? 1'b0 : 
                (N19)? 1'b0 : 
                (N20)? 1'b0 : 
                (N21)? 1'b0 : 
                (N22)? 1'b0 : 
                (N23)? 1'b0 : 
                (N24)? 1'b0 : 
                (N25)? 1'b0 : 
                (N26)? 1'b1 : 1'b0;
  assign { N720, N719, N718, N717, N716 } = (N27)? { N714, N713, N712, N711, N710 } : 
                                            (N546)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N27 = N545;
  assign N721 = (N27)? N715 : 
                (N546)? 1'b1 : 1'b0;
  assign N835 = (N28)? 1'b1 : 
                (N834)? N803 : 1'b0;
  assign N28 = N833;
  assign { N855, N854 } = (N29)? { 1'b1, 1'b0 } : 
                          (N853)? { N835, N835 } : 1'b0;
  assign N29 = N852;
  assign { N895, N894, N893, N892 } = (N30)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                      (N891)? { N852, N852, N855, N854 } : 1'b0;
  assign N30 = N890;
  assign { N913, N912, N911, N910, N909 } = (N31)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                            (N908)? { N895, N894, N890, N893, N892 } : 1'b0;
  assign N31 = N907;
  assign { N932, N931, N930, N929, N928 } = (N32)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                            (N927)? { N913, N912, N911, N910, N909 } : 1'b0;
  assign N32 = N926;
  assign { N938, N937, N936 } = (N33)? { 1'b0, 1'b1, 1'b0 } : 
                                (N34)? { N930, N929, N928 } : 1'b0;
  assign N33 = N935;
  assign N34 = N934;
  assign { N990, N989, N988 } = (N35)? { 1'b0, 1'b1, 1'b1 } : 
                                (N987)? { N926, N932, N931 } : 1'b0;
  assign N35 = N986;
  assign N1002 = (N36)? N1000 : 
                 (N37)? 1'b0 : 1'b0;
  assign N36 = N2723;
  assign N37 = N2722;
  assign { N1026, N1025 } = (N38)? { 1'b1, 1'b1 } : 
                            (N39)? { 1'b1, 1'b0 } : 
                            (N1024)? { 1'b0, N2723 } : 1'b0;
  assign N38 = N1006;
  assign N39 = N1022;
  assign { N1124, N1123, N1122, N1121, N1120 } = (N40)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                 (N41)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                                 (N42)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                 (N43)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                                 (N44)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                                 (N45)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                 (N46)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                                 (N47)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                                                 (N48)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                                 (N49)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                 (N50)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                 (N51)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                                 (N52)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                                 (N53)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                                 (N1119)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N40 = N1052;
  assign N41 = N1053;
  assign N42 = N1054;
  assign N43 = N593;
  assign N44 = N1062;
  assign N45 = N599;
  assign N46 = N1067;
  assign N47 = N1080;
  assign N48 = N1086;
  assign N49 = N1093;
  assign N50 = N1095;
  assign N51 = N1098;
  assign N52 = N1101;
  assign N53 = N1105;
  assign N1125 = (N40)? 1'b0 : 
                 (N41)? 1'b0 : 
                 (N42)? 1'b0 : 
                 (N43)? 1'b0 : 
                 (N44)? 1'b0 : 
                 (N45)? 1'b0 : 
                 (N46)? 1'b0 : 
                 (N47)? 1'b0 : 
                 (N48)? 1'b0 : 
                 (N49)? 1'b0 : 
                 (N50)? 1'b0 : 
                 (N51)? 1'b0 : 
                 (N52)? 1'b0 : 
                 (N53)? 1'b0 : 
                 (N1119)? 1'b1 : 1'b0;
  assign { N1130, N1129, N1128, N1127, N1126 } = (N54)? { N1124, N1123, N1122, N1121, N1120 } : 
                                                 (N1030)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N54 = N1029;
  assign N1131 = (N54)? N1125 : 
                 (N1030)? 1'b1 : 1'b0;
  assign N1212 = (N55)? 1'b1 : 
                 (N1211)? N1182 : 1'b0;
  assign N55 = N1210;
  assign { N1234, N1233, N1232 } = (N56)? { 1'b0, 1'b1, 1'b1 } : 
                                   (N1231)? { N1153, N1153, N1212 } : 1'b0;
  assign N56 = N1230;
  assign { N1263, N1262, N1261, N1260, N1259 } = (N57)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                                 (N1258)? { N1182, N1234, N1230, N1233, N1232 } : 1'b0;
  assign N57 = N1257;
  assign { N1310, N1309, N1308, N1307, N1306 } = (N58)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                                                 (N1305)? { N1262, N1261, N1260, N1257, N1259 } : 1'b0;
  assign N58 = N1304;
  assign { N1367, N1366, N1365, N1364 } = (N59)? { 1'b1, 1'b1, 1'b0, 1'b0 } : 
                                          (N60)? { 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                          (N61)? { 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                          (N62)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                                          (N63)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                          (N64)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                          (N65)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N59 = N1355;
  assign N60 = N1356;
  assign N61 = N1358;
  assign N62 = N1359;
  assign N63 = N1361;
  assign N64 = N1362;
  assign N65 = N1363;
  assign N1368 = (N59)? 1'b0 : 
                 (N60)? 1'b0 : 
                 (N61)? 1'b0 : 
                 (N62)? 1'b0 : 
                 (N63)? 1'b0 : 
                 (N64)? 1'b0 : 
                 (N65)? 1'b1 : 1'b0;
  assign { N1372, N1371, N1370, N1369 } = (N66)? { N1367, N1366, N1365, N1364 } : 
                                          (N67)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N66 = N1353;
  assign N67 = N1352;
  assign N1373 = (N66)? N1368 : 
                 (N67)? 1'b1 : 1'b0;
  assign { N1380, N1379, N1378 } = (N59)? { 1'b0, 1'b0, 1'b0 } : 
                                   (N60)? { 1'b0, 1'b0, 1'b1 } : 
                                   (N68)? { 1'b0, 1'b1, 1'b0 } : 
                                   (N61)? { 1'b1, 1'b0, 1'b0 } : 
                                   (N62)? { 1'b1, 1'b0, 1'b1 } : 
                                   (N63)? { 1'b1, 1'b1, 1'b0 } : 
                                   (N69)? { 1'b0, 1'b1, 1'b1 } : 
                                   (N64)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N68 = N1376;
  assign N69 = N1377;
  assign N1381 = (N59)? 1'b0 : 
                 (N60)? 1'b0 : 
                 (N68)? 1'b0 : 
                 (N61)? 1'b0 : 
                 (N62)? 1'b0 : 
                 (N63)? 1'b0 : 
                 (N69)? 1'b0 : 
                 (N64)? 1'b1 : 1'b0;
  assign { N1384, N1383, N1382 } = (N70)? { N1380, N1379, N1378 } : 
                                   (N71)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N70 = N1375;
  assign N71 = N1374;
  assign N1385 = (N70)? N1381 : 
                 (N71)? 1'b1 : 1'b0;
  assign N1402 = (N72)? preissue_pkt_i[14] : 
                 (N1401)? 1'b0 : 1'b0;
  assign N72 = N1400;
  assign N1403 = (N72)? N2302 : 
                 (N1401)? 1'b1 : 1'b0;
  assign { N1415, N1414 } = (N73)? { 1'b0, 1'b0 } : 
                            (N74)? { 1'b0, 1'b1 } : 
                            (N75)? { 1'b1, 1'b0 } : 
                            (N76)? { 1'b1, 1'b1 } : 1'b0;
  assign N73 = N1410;
  assign N74 = N1411;
  assign N75 = N1412;
  assign N76 = N1413;
  assign { N1417, N1416 } = (N77)? { N1415, N1414 } : 
                            (N1409)? { 1'b0, 1'b0 } : 1'b0;
  assign N77 = N1408;
  assign N1418 = ~N1408;
  assign N1424 = (N78)? preissue_pkt_i[14] : 
                 (N1423)? 1'b0 : 1'b0;
  assign N78 = N1422;
  assign N1425 = (N78)? N2302 : 
                 (N1423)? 1'b1 : 1'b0;
  assign { N1503, N1502, N1501, N1500, N1499, N1498, N1497 } = (N79)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N80)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                                               (N81)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                                                               (N82)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                                               (N83)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                               (N84)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N85)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                                               (N86)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                                               (N87)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                                               (N88)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N89)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N90)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N91)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N79 = N1431;
  assign N80 = N1434;
  assign N81 = N1437;
  assign N82 = N1440;
  assign N83 = N1445;
  assign N84 = N1448;
  assign N85 = N1452;
  assign N86 = N1455;
  assign N87 = N1469;
  assign N88 = N1473;
  assign N89 = N1476;
  assign N90 = N1485;
  assign N91 = N1505;
  assign N1504 = (N79)? 1'b0 : 
                 (N80)? 1'b1 : 
                 (N81)? 1'b0 : 
                 (N82)? 1'b0 : 
                 (N83)? 1'b0 : 
                 (N84)? 1'b0 : 
                 (N85)? 1'b0 : 
                 (N86)? 1'b0 : 
                 (N87)? 1'b0 : 
                 (N88)? 1'b0 : 
                 (N89)? 1'b0 : 
                 (N90)? 1'b0 : 
                 (N91)? 1'b0 : 1'b0;
  assign N1505 = ~N1496;
  assign N1506 = (N92)? N1504 : 
                 (N1428)? 1'b0 : 1'b0;
  assign N92 = N1427;
  assign N1507 = (N92)? N1505 : 
                 (N1428)? 1'b1 : 1'b0;
  assign { N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508 } = (N92)? { N1503, N1448, N1502, N1501, N1500, N1499, N1498, N1497 } : 
                                                                      (N1428)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1675 = (N93)? N2302 : 
                 (N2688)? N1663 : 
                 (N2690)? N1664 : 
                 (N2692)? N1665 : 
                 (N2694)? N1621 : 
                 (N2697)? decode_info_i[12] : 
                 (N2700)? N1666 : 
                 (N2703)? N1666 : 
                 (N1674)? 1'b0 : 1'b0;
  assign N93 = N1649;
  assign N1676 = (N94)? decode_info_i[10] : 
                 (N95)? 1'b0 : 
                 (N96)? 1'b0 : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N94 = N1533;
  assign N95 = N1541;
  assign N96 = N1550;
  assign N97 = N1556;
  assign N98 = N1563;
  assign N99 = N1588;
  assign N100 = N1602;
  assign N101 = N1603;
  assign N1677 = (N94)? decode_info_i[11] : 
                 (N95)? 1'b0 : 
                 (N96)? 1'b0 : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N1678 = (N94)? decode_info_i[12] : 
                 (N95)? 1'b0 : 
                 (N96)? 1'b0 : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N1679 = (N94)? 1'b0 : 
                 (N95)? N1612 : 
                 (N96)? 1'b0 : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N1680 = (N94)? 1'b0 : 
                 (N95)? N1613 : 
                 (N96)? 1'b0 : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N1681 = (N94)? 1'b0 : 
                 (N95)? 1'b0 : 
                 (N96)? N1614 : 
                 (N97)? N1666 : 
                 (N98)? N1616 : 
                 (N99)? decode_info_i[7] : 
                 (N100)? N1619 : 
                 (N101)? N1675 : 
                 (N1611)? 1'b1 : 1'b0;
  assign N1682 = (N94)? 1'b0 : 
                 (N95)? 1'b0 : 
                 (N96)? decode_info_i[9] : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N1683 = (N94)? 1'b0 : 
                 (N95)? 1'b0 : 
                 (N96)? 1'b0 : 
                 (N97)? N1615 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N1684 = (N94)? 1'b0 : 
                 (N95)? 1'b0 : 
                 (N96)? 1'b0 : 
                 (N97)? 1'b0 : 
                 (N98)? N1617 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N1685 = (N94)? 1'b0 : 
                 (N95)? 1'b0 : 
                 (N96)? 1'b0 : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? N1618 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign { N1689, N1688, N1687, N1686 } = (N94)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                          (N95)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                          (N96)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                          (N97)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                          (N98)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                          (N99)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                          (N100)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                          (N101)? { N2707, 1'b0, N1621, N1643 } : 
                                          (N1611)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1690 = (N94)? 1'b0 : 
                 (N95)? 1'b0 : 
                 (N96)? 1'b0 : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? N1620 : 
                 (N101)? 1'b0 : 
                 (N1611)? 1'b0 : 1'b0;
  assign N1691 = (N102)? N1690 : 
                 (N103)? 1'b0 : 1'b0;
  assign N102 = N1518;
  assign N103 = N1517;
  assign N1692 = (N102)? N1676 : 
                 (N103)? 1'b0 : 1'b0;
  assign N1693 = (N102)? N1677 : 
                 (N103)? 1'b0 : 1'b0;
  assign N1694 = (N102)? N1678 : 
                 (N103)? 1'b0 : 1'b0;
  assign N1695 = (N102)? N1679 : 
                 (N103)? 1'b0 : 1'b0;
  assign N1696 = (N102)? N1680 : 
                 (N103)? 1'b0 : 1'b0;
  assign N1697 = (N102)? N1681 : 
                 (N103)? 1'b1 : 1'b0;
  assign N1698 = (N102)? N1682 : 
                 (N103)? 1'b0 : 1'b0;
  assign N1699 = (N102)? N1683 : 
                 (N103)? 1'b0 : 1'b0;
  assign N1700 = (N102)? N1684 : 
                 (N103)? 1'b0 : 1'b0;
  assign N1701 = (N102)? N1685 : 
                 (N103)? 1'b0 : 1'b0;
  assign { N1705, N1704, N1703, N1702 } = (N102)? { N1689, N1688, N1687, N1686 } : 
                                          (N103)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2256, N2255, N2254, N2253, N2252, N2251 } = (N104)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, N2048, 1'b0, 1'b0, 1'b0, 1'b0, N2061, 1'b0 } : 
                                                                                                                (N105)? { 1'b1, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, N2090, 1'b0, 1'b0, 1'b0, 1'b1, N1868, N2105 } : 
                                                                                                                (N106)? { 1'b1, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, N2124, 1'b0, 1'b0, 1'b1, 1'b1, N1868, N2134 } : 
                                                                                                                (N107)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, N2169, N1868, 1'b0, 1'b0, 1'b1, 1'b0, N2180, 1'b0 } : 
                                                                                                                (N108)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, N2199, N1868, 1'b0, 1'b1, 1'b0, 1'b0, N2209, 1'b0 } : 
                                                                                                                (N109)? { 1'b1, 1'b0, N2707, 1'b0, 1'b0, 1'b1, 1'b0, N2229, 1'b0, 1'b1, 1'b1, 1'b0, N1868, N2229 } : 
                                                                                                                (N110)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, N2250, N1868, 1'b0, 1'b1, 1'b0, 1'b1, N2250, 1'b0 } : 
                                                                                                                (N111)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, N1868, 1'b0, 1'b1, 1'b1, 1'b1, N1868, 1'b0 } : 
                                                                                                                (N112)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, N1868, 1'b1, 1'b0, 1'b0, 1'b0, N1868, 1'b0 } : 
                                                                                                                (N113)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, N1868, 1'b1, 1'b0, 1'b0, 1'b1, N1868, 1'b0 } : 
                                                                                                                (N114)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, N1868, 1'b1, 1'b1, 1'b1, 1'b0, N1868, 1'b0 } : 
                                                                                                                (N115)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, N1868, 1'b1, 1'b1, 1'b0, 1'b1, N1868, 1'b0 } : 
                                                                                                                (N116)? { 1'b1, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, N1868, 1'b1, 1'b0, 1'b1, 1'b0, N1868, 1'b0 } : 
                                                                                                                (N117)? { 1'b1, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, N1868, 1'b1, 1'b0, 1'b1, 1'b1, N1868, 1'b0 } : 
                                                                                                                (N118)? { 1'b1, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, N1868, 1'b1, 1'b1, 1'b0, 1'b0, N1868, 1'b0 } : 
                                                                                                                (N119)? { 1'b1, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, N1868, 1'b1, 1'b1, 1'b1, 1'b1, N1868, 1'b0 } : 
                                                                                                                (N120)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, N1868, 1'b0, 1'b0, 1'b0, 1'b0, N1868, 1'b0 } : 
                                                                                                                (N121)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, N1868, 1'b0, 1'b0, 1'b0, 1'b1, N1868, 1'b0 } : 
                                                                                                                (N122)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, N1868, 1'b0, 1'b0, 1'b1, 1'b0, N1868, 1'b0 } : 
                                                                                                                (N123)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, N1868, 1'b1, 1'b0, 1'b0, 1'b0, N1868, 1'b0 } : 
                                                                                                                (N124)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, N1868, 1'b1, 1'b0, 1'b0, 1'b1, N1868, 1'b0 } : 
                                                                                                                (N125)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1868, 1'b0, 1'b0, 1'b0, 1'b0, N1868, 1'b0 } : 1'b0;
  assign N104 = N1879;
  assign N105 = N1893;
  assign N106 = N1900;
  assign N107 = N1908;
  assign N108 = N1913;
  assign N109 = N1921;
  assign N110 = N1927;
  assign N111 = N1935;
  assign N112 = N1938;
  assign N113 = N1945;
  assign N114 = N1952;
  assign N115 = N1955;
  assign N116 = N1960;
  assign N117 = N1965;
  assign N118 = N1968;
  assign N119 = N1972;
  assign N120 = N1980;
  assign N121 = N1985;
  assign N122 = N1990;
  assign N123 = N1993;
  assign N124 = N2001;
  assign N125 = N2034;
  assign N2259 = (N104)? N2048 : 
                 (N2258)? N1868 : 1'b0;
  assign N2268 = (N104)? N2302 : 
                 (N105)? N2302 : 
                 (N106)? N2302 : 
                 (N107)? N2302 : 
                 (N108)? N2302 : 
                 (N109)? N2302 : 
                 (N110)? N2302 : 
                 (N111)? N2302 : 
                 (N112)? N2302 : 
                 (N113)? N2302 : 
                 (N114)? N2302 : 
                 (N115)? N2302 : 
                 (N116)? N2302 : 
                 (N117)? N2302 : 
                 (N118)? N2302 : 
                 (N119)? N2302 : 
                 (N120)? N2302 : 
                 (N121)? N2302 : 
                 (N122)? N2302 : 
                 (N123)? N2302 : 
                 (N124)? N2302 : 
                 (N125)? 1'b1 : 1'b0;
  assign { N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269 } = (N126)? { N2267, N2266, N2265, N2264, N2263, N2262, N1913, N2261, N2260, N2259, N2256, N2255, N2254, N2253, N2252, N2251 } : 
                                                                                                                              (N1873)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1868, N1868, 1'b0, 1'b0, 1'b0, 1'b0, N1868, 1'b0 } : 1'b0;
  assign N126 = N1872;
  assign N2285 = (N126)? N2268 : 
                 (N1873)? 1'b1 : 1'b0;
  assign { N2298, N2297, N2296 } = (N127)? { 1'b0, 1'b1, 1'b1 } : 
                                   (N128)? { 1'b1, 1'b0, 1'b0 } : 
                                   (N129)? { 1'b1, 1'b0, 1'b1 } : 
                                   (N130)? { 1'b1, 1'b1, 1'b0 } : 1'b0;
  assign N127 = N2290;
  assign N128 = N2292;
  assign N129 = N2294;
  assign N130 = N2295;
  assign { N2301, N2300, N2299 } = (N131)? { N2298, N2297, N2296 } : 
                                   (N2289)? { 1'b0, 1'b1, 1'b1 } : 1'b0;
  assign N131 = N2288;
  assign { N2373, N2372, N2371, N2370, N2369, N2368 } = (N132)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                                                        (N133)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                        (N134)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                                        (N135)? { 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                                                        (N136)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                                                        (N137)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N138)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                                                        (N139)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                                        (N140)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                                        (N141)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                                        (N142)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                                                        (N143)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                        (N144)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                                                        (N145)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                                        (N146)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                                        (N147)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                                        (N148)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                        (N149)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                                        (N150)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N151)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                        (N152)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                                        (N153)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                                        (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N132 = N2341;
  assign N133 = N2343;
  assign N134 = N2344;
  assign N135 = N2346;
  assign N136 = N2347;
  assign N137 = N2348;
  assign N138 = N2350;
  assign N139 = N2352;
  assign N140 = N2353;
  assign N141 = N2354;
  assign N142 = N2355;
  assign N143 = N2356;
  assign N144 = N2357;
  assign N145 = N2358;
  assign N146 = N2359;
  assign N147 = N2360;
  assign N148 = N2361;
  assign N149 = N2362;
  assign N150 = N2363;
  assign N151 = N2364;
  assign N152 = N2365;
  assign N153 = N2366;
  assign N154 = N2367;
  assign N2374 = (N132)? 1'b0 : 
                 (N133)? 1'b0 : 
                 (N134)? 1'b0 : 
                 (N135)? 1'b0 : 
                 (N136)? 1'b0 : 
                 (N137)? 1'b0 : 
                 (N138)? 1'b0 : 
                 (N139)? 1'b0 : 
                 (N140)? 1'b0 : 
                 (N141)? 1'b0 : 
                 (N142)? 1'b0 : 
                 (N143)? 1'b0 : 
                 (N144)? 1'b0 : 
                 (N145)? 1'b0 : 
                 (N146)? 1'b0 : 
                 (N147)? 1'b0 : 
                 (N148)? 1'b0 : 
                 (N149)? 1'b0 : 
                 (N150)? 1'b0 : 
                 (N151)? 1'b0 : 
                 (N152)? 1'b0 : 
                 (N153)? 1'b0 : 
                 (N154)? 1'b1 : 1'b0;
  assign { N2380, N2379, N2378, N2377, N2376, N2375 } = (N155)? { N2373, N2372, N2371, N2370, N2369, N2368 } : 
                                                        (N2338)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N155 = N2337;
  assign N2381 = (N155)? N2374 : 
                 (N2338)? 1'b1 : 1'b0;
  assign N2470 = (N156)? 1'b0 : 
                 (N157)? 1'b0 : 
                 (N158)? 1'b0 : 
                 (N159)? 1'b0 : 
                 (N160)? N2381 : 1'b0;
  assign N156 = N2407;
  assign N157 = N2412;
  assign N158 = N2430;
  assign N159 = N2456;
  assign N160 = N2469;
  assign { N2527, N2526, N2519, N2518, N2517, N2516, N2509, N2508, N2507, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2489, N2488, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471 } = (N178)? { N349, 1'b0, 1'b0, N347, N2707, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N347, 1'b0, 1'b0, N803, N479, N413, N414, 1'b0, 1'b0, N720, N719, 1'b0, N718, N717, N716, 1'b0, N392, N990, N989, N988, N938, N937, N936 } : 
                                                                                                                                                                                                                                                     (N186)? { 1'b1, 1'b0, 1'b0, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1326, N1263, N1026, N1025, 1'b0, 1'b0, N1130, N1129, 1'b0, N1128, N1127, N1126, 1'b0, N1002, N1310, N1309, N1308, N1307, N1306, 1'b0 } : 
                                                                                                                                                                                                                                                     (N190)? { 1'b1, 1'b0, 1'b0, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N192)? { 1'b1, 1'b0, 1'b0, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N196)? { 1'b1, 1'b0, 1'b0, 1'b0, N2707, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N200)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1372, N1371, N1370, N1369, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                                                                     (N161)? { 1'b0, 1'b1, 1'b0, 1'b0, N2707, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1384, N1383, N1382, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N211)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1400, 1'b0, 1'b0, 1'b0, N1400, N1402, N1395, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N215)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1408, 1'b0, N1417, N1416, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N217)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1422, 1'b0, 1'b0, N1422, 1'b0, N1424, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N220)? { 1'b0, N1512, 1'b0, 1'b0, 1'b0, 1'b0, N1515, 1'b0, N1514, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1512, N1512, N1511, N1510, N1509, N1508, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N223)? { 1'b0, 1'b0, 1'b0, 1'b0, N1705, 1'b0, N1704, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N227)? { 1'b0, 1'b0, N2283, N2280, N2282, N2281, 1'b0, 1'b0, 1'b0, 1'b0, N2280, 1'b0, N2279, 1'b0, N2278, 1'b0, N2277, N2276, N2275, 1'b0, 1'b0, N2274, N2273, N2272, N2271, N2270, N2269, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N234)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N2709, N2709, 1'b0, 1'b0, 1'b0, N2301, N2300, N2299, N2709, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N238)? { 1'b0, 1'b1, 1'b0, 1'b0, N2707, 1'b0, 1'b0, N2333, N2334, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N2380, N2379, N2378, N2377, N2376, N2375, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                     (N249)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N161 = N209;
  assign N2487 = (N234)? N2709 : 
                 (N2486)? 1'b0 : 1'b0;
  assign { N2520, N2493, N2492 } = (N178)? { N266, N538, N392 } : 
                                   (N2491)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N2521, N2504, N2503 } = (N223)? { 1'b1, N1703, N1702 } : 
                                   (N2502)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2506 = (N220)? N1513 : 
                 (N2505)? 1'b0 : 1'b0;
  assign { N2513, N2512 } = (N196)? { N1337, N1347 } : 
                            (N2511)? { 1'b0, 1'b0 } : 1'b0;
  assign N2515 = (N200)? 1'b1 : 
                 (N2514)? 1'b0 : 1'b0;
  assign N2523 = (N211)? 1'b1 : 
                 (N2522)? 1'b0 : 1'b0;
  assign N2525 = (N227)? N2284 : 
                 (N2524)? 1'b0 : 1'b0;
  assign N2528 = (N178)? N721 : 
                 (N186)? N1131 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? N1349 : 
                 (N200)? N1373 : 
                 (N161)? N1385 : 
                 (N211)? N1403 : 
                 (N215)? N1418 : 
                 (N217)? N1425 : 
                 (N220)? N1507 : 
                 (N223)? N1697 : 
                 (N227)? N2285 : 
                 (N234)? N2302 : 
                 (N238)? N2470 : 
                 (N249)? 1'b1 : 1'b0;
  assign N2529 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? N1506 : 
                 (N223)? 1'b0 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2530 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1700 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2531 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1701 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2532 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1691 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2533 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1703 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2534 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1692 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2535 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1693 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2536 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1694 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2537 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1695 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2538 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1696 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2539 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1698 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign N2540 = (N178)? 1'b0 : 
                 (N186)? 1'b0 : 
                 (N190)? 1'b0 : 
                 (N192)? 1'b0 : 
                 (N196)? 1'b0 : 
                 (N200)? 1'b0 : 
                 (N161)? 1'b0 : 
                 (N211)? 1'b0 : 
                 (N215)? 1'b0 : 
                 (N217)? 1'b0 : 
                 (N220)? 1'b0 : 
                 (N223)? N1699 : 
                 (N227)? 1'b0 : 
                 (N234)? 1'b0 : 
                 (N238)? 1'b0 : 
                 (N249)? 1'b0 : 1'b0;
  assign dret_o = (N162)? N2539 : 
                  (N174)? 1'b0 : 1'b0;
  assign N162 = N173;
  assign mret_o = (N162)? N2540 : 
                  (N174)? 1'b0 : 1'b0;
  assign { decode_o[53:46], decode_o[40:32], decode_o[30:20], decode_o[18:8], decode_o[6:0] } = (N162)? { N2527, N2526, N2525, N2523, N2521, N2520, N2519, N2518, N2517, N2516, N2515, N2513, N2512, N2509, N2508, N2507, N2506, N2504, N2503, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2489, N2488, N2487, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471 } : 
                                                                                                (N174)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign illegal_instr_o = (N162)? N2528 : 
                           (N174)? 1'b1 : 1'b0;
  assign fencei_o = (N162)? N2529 : 
                    (N174)? 1'b0 : 1'b0;
  assign sret_o = (N162)? N2530 : 
                  (N174)? 1'b0 : 1'b0;
  assign wfi_o = (N162)? N2531 : 
                 (N174)? 1'b0 : 1'b0;
  assign sfence_vma_o = (N162)? N2532 : 
                        (N174)? 1'b0 : 1'b0;
  assign csrw_o = (N162)? N2533 : 
                  (N174)? 1'b0 : 1'b0;
  assign ecall_m_o = (N162)? N2534 : 
                     (N174)? 1'b0 : 1'b0;
  assign ecall_s_o = (N162)? N2535 : 
                     (N174)? 1'b0 : 1'b0;
  assign ecall_u_o = (N162)? N2536 : 
                     (N174)? 1'b0 : 1'b0;
  assign dbreak_o = (N162)? N2537 : 
                    (N174)? 1'b0 : 1'b0;
  assign ebreak_o = (N162)? N2538 : 
                    (N174)? 1'b0 : 1'b0;
  assign { N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579 } = (N163)? { preissue_pkt_i[33:14], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                              (N164)? { preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[21:14], preissue_pkt_i[22:22], preissue_pkt_i[32:23], 1'b0 } : 
                                                                                                                                                                                                                                              (N165)? { preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[9:9], preissue_pkt_i[32:27], preissue_pkt_i[13:10], 1'b0 } : 
                                                                                                                                                                                                                                              (N166)? { preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:27], preissue_pkt_i[13:9] } : 
                                                                                                                                                                                                                                              (N167)? { preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:33], preissue_pkt_i[33:22] } : 
                                                                                                                                                                                                                                              (N168)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N163 = N2547;
  assign N164 = N2552;
  assign N165 = N2555;
  assign N166 = N2559;
  assign N167 = N2570;
  assign N168 = N2578;
  assign { N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611 } = (N162)? { N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579 } : 
                                                                                                                                                                                                                                              (N174)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign imm_o = (N169)? { N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N2135, N1287, N462, N2303, N393, N2684, N523, N2685, N2686, N1183, N2079, N2035 } : 
                 (N170)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                 (N171)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                 (N172)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                 (N2683)? { N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611 } : 1'b0;
  assign N169 = N2649;
  assign N170 = N2657;
  assign N171 = N2665;
  assign N172 = N2679;
  assign N174 = ~N173;
  assign N178 = N2728 | N2729;
  assign N2728 = ~N175;
  assign N2729 = ~N177;
  assign N186 = N2730 | N2731;
  assign N2730 = ~N182;
  assign N2731 = ~N185;
  assign N190 = ~N189;
  assign N192 = ~N191;
  assign N196 = N2732 | N2733;
  assign N2732 = ~N194;
  assign N2733 = ~N195;
  assign N200 = ~N199;
  assign N201 = ~preissue_pkt_i[8];
  assign N202 = ~preissue_pkt_i[7];
  assign N203 = ~preissue_pkt_i[6];
  assign N204 = ~preissue_pkt_i[5];
  assign N205 = ~preissue_pkt_i[4];
  assign N211 = ~N210;
  assign N215 = ~N214;
  assign N217 = ~N216;
  assign N220 = ~N219;
  assign N223 = ~N222;
  assign N227 = ~N226;
  assign N234 = N2738 | N2739;
  assign N2738 = N2736 | N2737;
  assign N2736 = N2734 | N2735;
  assign N2734 = ~N229;
  assign N2735 = ~N230;
  assign N2737 = ~N232;
  assign N2739 = ~N233;
  assign N238 = ~N237;
  assign N249 = N240 | N2742;
  assign N2742 = N242 | N2741;
  assign N2741 = N243 | N2740;
  assign N2740 = N246 | N248;
  assign N348 = N347 | N266;
  assign N546 = ~N545;
  assign N580 = N2758 | N579;
  assign N2758 = N2757 | N578;
  assign N2757 = N2756 | N577;
  assign N2756 = N2755 | N576;
  assign N2755 = N2754 | N574;
  assign N2754 = N2753 | N573;
  assign N2753 = N2752 | N571;
  assign N2752 = N2751 | N570;
  assign N2751 = N2750 | N568;
  assign N2750 = N2749 | N566;
  assign N2749 = N2748 | N564;
  assign N2748 = N2747 | N563;
  assign N2747 = N2746 | N561;
  assign N2746 = N2745 | N560;
  assign N2745 = N2744 | N558;
  assign N2744 = N2743 | N554;
  assign N2743 = N549 | N552;
  assign N603 = N601 | N602;
  assign N611 = N2762 | N610;
  assign N2762 = N2761 | N609;
  assign N2761 = N2760 | N608;
  assign N2760 = N2759 | N607;
  assign N2759 = N605 | N606;
  assign N614 = N612 | N613;
  assign N630 = N628 | N629;
  assign N639 = N637 | N638;
  assign N642 = N640 | N641;
  assign N645 = N643 | N644;
  assign N649 = N646 | N648;
  assign N709 = N652 | N2791;
  assign N2791 = N656 | N2790;
  assign N2790 = N658 | N2789;
  assign N2789 = N660 | N2788;
  assign N2788 = N662 | N2787;
  assign N2787 = N664 | N2786;
  assign N2786 = N665 | N2785;
  assign N2785 = N667 | N2784;
  assign N2784 = N669 | N2783;
  assign N2783 = N671 | N2782;
  assign N2782 = N673 | N2781;
  assign N2781 = N675 | N2780;
  assign N2780 = N678 | N2779;
  assign N2779 = N680 | N2778;
  assign N2778 = N681 | N2777;
  assign N2777 = N682 | N2776;
  assign N2776 = N685 | N2775;
  assign N2775 = N687 | N2774;
  assign N2774 = N689 | N2773;
  assign N2773 = N691 | N2772;
  assign N2772 = N694 | N2771;
  assign N2771 = N695 | N2770;
  assign N2770 = N699 | N2769;
  assign N2769 = N700 | N2768;
  assign N2768 = N701 | N2767;
  assign N2767 = N702 | N2766;
  assign N2766 = N703 | N2765;
  assign N2765 = N704 | N2764;
  assign N2764 = N706 | N2763;
  assign N2763 = N707 | N708;
  assign N834 = ~N833;
  assign N853 = ~N852;
  assign N891 = ~N890;
  assign N908 = ~N907;
  assign N927 = ~N926;
  assign N987 = ~N986;
  assign N1023 = N1022 | N1006;
  assign N1024 = ~N1023;
  assign N1030 = ~N1029;
  assign N1052 = N2800 | N1051;
  assign N2800 = N2799 | N1050;
  assign N2799 = N2798 | N1047;
  assign N2798 = N2797 | N1045;
  assign N2797 = N2796 | N1043;
  assign N2796 = N2795 | N1042;
  assign N2795 = N2794 | N1040;
  assign N2794 = N2793 | N1038;
  assign N2793 = N2792 | N1037;
  assign N2792 = N1031 | N1032;
  assign N1062 = N2801 | N597;
  assign N2801 = N1057 | N1061;
  assign N1067 = N1064 | N1066;
  assign N1080 = N2803 | N1079;
  assign N2803 = N2802 | N1077;
  assign N2802 = N1071 | N1074;
  assign N1106 = N1053 | N1052;
  assign N1107 = N1054 | N1106;
  assign N1108 = N593 | N1107;
  assign N1109 = N1062 | N1108;
  assign N1110 = N599 | N1109;
  assign N1111 = N1067 | N1110;
  assign N1112 = N1080 | N1111;
  assign N1113 = N1086 | N1112;
  assign N1114 = N1093 | N1113;
  assign N1115 = N1095 | N1114;
  assign N1116 = N1098 | N1115;
  assign N1117 = N1101 | N1116;
  assign N1118 = N1105 | N1117;
  assign N1119 = ~N1118;
  assign N1211 = ~N1210;
  assign N1231 = ~N1230;
  assign N1258 = ~N1257;
  assign N1305 = ~N1304;
  assign N1349 = ~N1348;
  assign N1353 = ~N1352;
  assign N1375 = ~N1374;
  assign N1401 = ~N1400;
  assign N1409 = ~N1408;
  assign N1423 = ~N1422;
  assign N1428 = ~N1427;
  assign N1486 = N1434 | N1431;
  assign N1487 = N1437 | N1486;
  assign N1488 = N1440 | N1487;
  assign N1489 = N1445 | N1488;
  assign N1490 = N1448 | N1489;
  assign N1491 = N1452 | N1490;
  assign N1492 = N1455 | N1491;
  assign N1493 = N1469 | N1492;
  assign N1494 = N1473 | N1493;
  assign N1495 = N1476 | N1494;
  assign N1496 = N1485 | N1495;
  assign N1518 = ~N1517;
  assign N1519 = ~preissue_pkt_i[21];
  assign N1520 = ~preissue_pkt_i[20];
  assign N1521 = ~preissue_pkt_i[19];
  assign N1522 = ~preissue_pkt_i[18];
  assign N1523 = ~preissue_pkt_i[17];
  assign N1541 = ~N1540;
  assign N1550 = ~N1549;
  assign N1556 = ~N1555;
  assign N1563 = ~N1562;
  assign N1588 = ~N1587;
  assign N1589 = ~preissue_pkt_i[13];
  assign N1590 = ~preissue_pkt_i[12];
  assign N1591 = ~preissue_pkt_i[11];
  assign N1592 = ~preissue_pkt_i[10];
  assign N1593 = ~preissue_pkt_i[9];
  assign N1603 = N2807 | N1362;
  assign N2807 = N2806 | N1377;
  assign N2806 = N2805 | N1361;
  assign N2805 = N2804 | N1376;
  assign N2804 = N1356 | N1359;
  assign N1604 = N1541 | N1533;
  assign N1605 = N1550 | N1604;
  assign N1606 = N1556 | N1605;
  assign N1607 = N1563 | N1606;
  assign N1608 = N1588 | N1607;
  assign N1609 = N1602 | N1608;
  assign N1610 = N1603 | N1609;
  assign N1611 = ~N1610;
  assign N1612 = N2811 | N2812;
  assign N2811 = N2809 | N2810;
  assign N2809 = decode_info_i[9] | N2808;
  assign N2808 = decode_info_i[5] & decode_info_i[10];
  assign N2810 = decode_info_i[4] & decode_info_i[11];
  assign N2812 = decode_info_i[3] & decode_info_i[12];
  assign N1613 = ~N1612;
  assign N1614 = ~decode_info_i[9];
  assign N1615 = ~N1666;
  assign N1616 = decode_info_i[12] | N2813;
  assign N2813 = decode_info_i[8] & decode_info_i[11];
  assign N1617 = ~N1616;
  assign N1618 = N2814 & N1614;
  assign N2814 = ~decode_info_i[7];
  assign N1619 = N2815 | decode_info_i[12];
  assign N2815 = decode_info_i[11] & decode_info_i[6];
  assign N1620 = ~N1619;
  assign N1621 = N1642 | N2727;
  assign N1643 = N2816 | N2707;
  assign N2816 = ~N1642;
  assign N1649 = N2819 | N2820;
  assign N2819 = N2817 | N2818;
  assign N2817 = ~N1646;
  assign N2818 = ~N1647;
  assign N2820 = ~N1648;
  assign N1651 = ~N1650;
  assign N1656 = ~N1655;
  assign N1662 = ~N1661;
  assign N1663 = ~decode_info_i[1];
  assign N1664 = ~decode_info_i[0];
  assign N1665 = decode_info_i[11] & decode_info_i[6];
  assign N1666 = decode_info_i[11] | decode_info_i[12];
  assign N1667 = N2688 | N1649;
  assign N1668 = N2690 | N1667;
  assign N1669 = N2692 | N1668;
  assign N1670 = N2694 | N1669;
  assign N1671 = N2697 | N1670;
  assign N1672 = N2700 | N1671;
  assign N1673 = N2703 | N1672;
  assign N1674 = ~N1673;
  assign N1873 = ~N1872;
  assign N1879 = N1876 | N1878;
  assign N1893 = N2822 | N1892;
  assign N2822 = N2821 | N1891;
  assign N2821 = N1885 | N1888;
  assign N1900 = N2824 | N1899;
  assign N2824 = N2823 | N1898;
  assign N2823 = N1895 | N1897;
  assign N1908 = N2826 | N1907;
  assign N2826 = N2825 | N1906;
  assign N2825 = N1903 | N1904;
  assign N1913 = N2828 | N1912;
  assign N2828 = N2827 | N1911;
  assign N2827 = N1909 | N1910;
  assign N1921 = N1918 | N1920;
  assign N1927 = N1924 | N1926;
  assign N1935 = N1931 | N1934;
  assign N1938 = N1936 | N1937;
  assign N1945 = N1941 | N1944;
  assign N1952 = N1948 | N1951;
  assign N1955 = N1953 | N1954;
  assign N1960 = N1957 | N1959;
  assign N1965 = N1962 | N1964;
  assign N1968 = N1966 | N1967;
  assign N1972 = N1970 | N1971;
  assign N1980 = N1977 | N1979;
  assign N1985 = N1981 | N1984;
  assign N1990 = N1988 | N1989;
  assign N1993 = N1991 | N1992;
  assign N2001 = N1997 | N2000;
  assign N2034 = N2004 | N2852;
  assign N2852 = N2007 | N2851;
  assign N2851 = N2008 | N2850;
  assign N2850 = N2009 | N2849;
  assign N2849 = N2010 | N2848;
  assign N2848 = N2012 | N2847;
  assign N2847 = N2013 | N2846;
  assign N2846 = N2014 | N2845;
  assign N2845 = N2015 | N2844;
  assign N2844 = N2016 | N2843;
  assign N2843 = N2017 | N2842;
  assign N2842 = N2019 | N2841;
  assign N2841 = N2020 | N2840;
  assign N2840 = N2021 | N2839;
  assign N2839 = N2024 | N2838;
  assign N2838 = N2025 | N2837;
  assign N2837 = N682 | N2836;
  assign N2836 = N2459 | N2835;
  assign N2835 = N2026 | N2834;
  assign N2834 = N2028 | N2833;
  assign N2833 = N2029 | N2832;
  assign N2832 = N2030 | N2831;
  assign N2831 = N2031 | N2830;
  assign N2830 = N2032 | N2829;
  assign N2829 = N2033 | N662;
  assign N2257 = ~N1879;
  assign N2258 = N2257;
  assign N2289 = ~N2288;
  assign N2292 = ~N2291;
  assign N2294 = ~N2293;
  assign N2302 = ~decode_info_i[2];
  assign N2334 = ~N2333;
  assign N2338 = ~N2337;
  assign N2367 = N2457 | N2861;
  assign N2861 = N2458 | N2860;
  assign N2860 = N2459 | N2859;
  assign N2859 = N2460 | N2858;
  assign N2858 = N2461 | N2857;
  assign N2857 = N2462 | N2856;
  assign N2856 = N2464 | N2855;
  assign N2855 = N2465 | N2854;
  assign N2854 = N2466 | N2853;
  assign N2853 = N2467 | N2468;
  assign N2407 = N2863 | N2406;
  assign N2863 = N2862 | N2403;
  assign N2862 = N2392 | N2397;
  assign N2412 = N2409 | N2411;
  assign N2430 = N2867 | N2429;
  assign N2867 = N2866 | N2427;
  assign N2866 = N2865 | N2424;
  assign N2865 = N2864 | N2422;
  assign N2864 = N2416 | N2419;
  assign N2456 = N2875 | N2455;
  assign N2875 = N2874 | N2453;
  assign N2874 = N2873 | N2450;
  assign N2873 = N2872 | N2448;
  assign N2872 = N2871 | N2444;
  assign N2871 = N2870 | N2442;
  assign N2870 = N2869 | N2439;
  assign N2869 = N2868 | N2437;
  assign N2868 = N2432 | N2434;
  assign N2469 = preissue_pkt_i[16] | N2893;
  assign N2893 = N2304 | N2892;
  assign N2892 = preissue_pkt_i[8] | N2891;
  assign N2891 = N1328 | N2890;
  assign N2890 = preissue_pkt_i[6] | N2889;
  assign N2889 = N1329 | N2888;
  assign N2888 = N1330 | N2887;
  assign N2887 = N395 | N2886;
  assign N2886 = N396 | N2885;
  assign N2885 = N2457 | N2884;
  assign N2884 = N2458 | N2883;
  assign N2883 = N2459 | N2882;
  assign N2882 = N2460 | N2881;
  assign N2881 = N2461 | N2880;
  assign N2880 = N2462 | N2879;
  assign N2879 = N2464 | N2878;
  assign N2878 = N2465 | N2877;
  assign N2877 = N2466 | N2876;
  assign N2876 = N2467 | N2468;
  assign N2485 = ~N234;
  assign N2486 = N2485;
  assign N2490 = ~N178;
  assign N2491 = N2490;
  assign N2502 = N222;
  assign N2505 = N219;
  assign N2510 = ~N196;
  assign N2511 = N2510;
  assign N2514 = N199;
  assign N2522 = N210;
  assign N2524 = N226;
  assign N2547 = N2894 | N2895;
  assign N2894 = ~N2544;
  assign N2895 = ~N2546;
  assign N2552 = ~N2551;
  assign N2555 = ~N2554;
  assign N2559 = N2896 | N2897;
  assign N2896 = ~N2557;
  assign N2897 = ~N2558;
  assign N2570 = N2903 | N2904;
  assign N2903 = N2901 | N2902;
  assign N2901 = N2899 | N2900;
  assign N2899 = N2898 | N2563;
  assign N2898 = ~N2560;
  assign N2900 = ~N2564;
  assign N2902 = ~N2567;
  assign N2904 = ~N2569;
  assign N2578 = N240 | N2908;
  assign N2908 = N2572 | N2907;
  assign N2907 = N241 | N2906;
  assign N2906 = N2574 | N2905;
  assign N2905 = N2576 | N2577;
  assign N2649 = N2645 | N2648;
  assign N2657 = N2654 | N2656;
  assign N2665 = N2661 | N2664;
  assign N2679 = N2674 | N2678;
  assign N2680 = N2657 | N2649;
  assign N2681 = N2665 | N2680;
  assign N2682 = N2679 | N2681;
  assign N2683 = ~N2682;
  assign N2684 = ~preissue_pkt_i[28];
  assign N2685 = ~preissue_pkt_i[26];
  assign N2686 = ~preissue_pkt_i[25];
  assign N2687 = ~N1649;
  assign N2688 = N1651 & N2687;
  assign N2689 = N2687 & N1650;
  assign N2690 = N1656 & N2689;
  assign N2691 = N2689 & N1655;
  assign N2692 = N1662 & N2691;
  assign N2693 = N2691 & N1661;
  assign N2694 = N2445 & N2693;
  assign N2695 = ~N2445;
  assign N2696 = N2693 & N2695;
  assign N2697 = N1986 & N2696;
  assign N2698 = ~N1986;
  assign N2699 = N2696 & N2698;
  assign N2700 = N2005 & N2699;
  assign N2701 = ~N2005;
  assign N2702 = N2699 & N2701;
  assign N2703 = N2457 & N2702;

endmodule



module bp_be_issue_queue
(
  clk_i,
  reset_i,
  en_i,
  clr_i,
  roll_i,
  read_i,
  read_cnt_i,
  read_size_i,
  cmt_i,
  cmt_cnt_i,
  cmt_size_i,
  fe_queue_i,
  fe_queue_v_i,
  fe_queue_ready_and_o,
  decode_info_i,
  preissue_pkt_o,
  issue_pkt_o
);

  input [3:0] read_cnt_i;
  input [3:0] read_size_i;
  input [3:0] cmt_cnt_i;
  input [3:0] cmt_size_i;
  input [173:0] fe_queue_i;
  input [12:0] decode_info_i;
  output [38:0] preissue_pkt_o;
  output [263:0] issue_pkt_o;
  input clk_i;
  input reset_i;
  input en_i;
  input clr_i;
  input roll_i;
  input read_i;
  input cmt_i;
  input fe_queue_v_i;
  output fe_queue_ready_and_o;
  wire [38:0] preissue_pkt_o;
  wire [263:0] issue_pkt_o;
  wire fe_queue_ready_and_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,
  N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,
  N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,ack,empty,empty_n,N69,N70,full,
  N71,N72,N73,N74,read_catchup,N75,N76,N77,N78,deq_catchup,N79,N80,N81,N82,N83,N84,
  N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,
  N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,
  N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,
  N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,
  N152,preissue_v,bypass_preissue,_0_net_,_2_net_,N153,queue_instr_raw_4__15_,
  queue_instr_raw_4__14_,queue_instr_raw_4__13_,queue_instr_raw_4__12_,
  queue_instr_raw_4__11_,queue_instr_raw_4__10_,queue_instr_raw_4__9_,queue_instr_raw_4__8_,
  queue_instr_raw_4__7_,queue_instr_raw_4__6_,queue_instr_raw_4__5_,
  queue_instr_raw_4__4_,queue_instr_raw_4__3_,queue_instr_raw_4__2_,queue_instr_raw_4__1_,
  queue_instr_raw_4__0_,queue_instr_raw_3__15_,queue_instr_raw_3__14_,queue_instr_raw_3__13_,
  queue_instr_raw_3__12_,queue_instr_raw_3__11_,queue_instr_raw_3__10_,
  queue_instr_raw_3__9_,queue_instr_raw_3__8_,queue_instr_raw_3__7_,queue_instr_raw_3__6_,
  queue_instr_raw_3__5_,queue_instr_raw_3__4_,queue_instr_raw_3__3_,
  queue_instr_raw_3__2_,queue_instr_raw_3__1_,queue_instr_raw_3__0_,queue_instr_raw_2__15_,
  queue_instr_raw_2__14_,queue_instr_raw_2__13_,queue_instr_raw_2__12_,
  queue_instr_raw_2__11_,queue_instr_raw_2__10_,queue_instr_raw_2__9_,queue_instr_raw_2__8_,
  queue_instr_raw_2__7_,queue_instr_raw_2__6_,queue_instr_raw_2__5_,queue_instr_raw_2__4_,
  queue_instr_raw_2__3_,queue_instr_raw_2__2_,queue_instr_raw_2__1_,
  queue_instr_raw_2__0_,queue_instr_raw_1__15_,queue_instr_raw_1__14_,queue_instr_raw_1__13_,
  queue_instr_raw_1__12_,queue_instr_raw_1__11_,queue_instr_raw_1__10_,
  queue_instr_raw_1__9_,queue_instr_raw_1__8_,queue_instr_raw_1__7_,queue_instr_raw_1__6_,
  queue_instr_raw_1__5_,queue_instr_raw_1__4_,queue_instr_raw_1__3_,queue_instr_raw_1__2_,
  queue_instr_raw_1__1_,queue_instr_raw_1__0_,queue_instr_raw_0__15_,
  queue_instr_raw_0__14_,queue_instr_raw_0__13_,queue_instr_raw_0__12_,queue_instr_raw_0__11_,
  queue_instr_raw_0__10_,queue_instr_raw_0__9_,queue_instr_raw_0__8_,
  queue_instr_raw_0__7_,queue_instr_raw_0__6_,queue_instr_raw_0__5_,queue_instr_raw_0__4_,
  queue_instr_raw_0__3_,queue_instr_raw_0__2_,queue_instr_raw_0__1_,
  queue_instr_raw_0__0_,N154,preissue_size_4__1_,preissue_size_4__0_,preissue_size_3__1_,
  preissue_size_3__0_,preissue_size_2__1_,preissue_size_2__0_,preissue_size_1__1_,
  preissue_size_1__0_,preissue_size_0__1_,preissue_size_0__0_,N155,N156,N157,N158,N159,N160,
  N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,
  N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,
  N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,
  N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,
  N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,
  N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,
  N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,
  N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
  N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,
  N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
  N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,
  N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,
  N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,
  N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,
  N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,
  N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,
  N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,
  N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,
  N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,
  N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,
  N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,
  N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,
  N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,
  N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,
  N593,N594,N595,N596,N597,N598,N599,preissue_pkt_r_irs1_v_,preissue_pkt_r_irs2_v_,
  preissue_pkt_r_frs1_v_,preissue_pkt_r_frs2_v_,preissue_pkt_r_frs3_v_,
  preissue_pkt_r_size__1_,preissue_pkt_r_size__0_,bypass_issue,_4_net_,_6_net_,
  fe_queue_lo_pc__38_,fe_queue_lo_pc__37_,fe_queue_lo_pc__36_,fe_queue_lo_pc__35_,
  fe_queue_lo_pc__34_,fe_queue_lo_pc__33_,fe_queue_lo_pc__32_,fe_queue_lo_pc__31_,
  fe_queue_lo_pc__30_,fe_queue_lo_pc__29_,fe_queue_lo_pc__28_,fe_queue_lo_pc__27_,
  fe_queue_lo_pc__26_,fe_queue_lo_pc__25_,fe_queue_lo_pc__24_,fe_queue_lo_pc__23_,
  fe_queue_lo_pc__22_,fe_queue_lo_pc__21_,fe_queue_lo_pc__20_,fe_queue_lo_pc__19_,
  fe_queue_lo_pc__18_,fe_queue_lo_pc__17_,fe_queue_lo_pc__16_,fe_queue_lo_pc__15_,
  fe_queue_lo_pc__14_,fe_queue_lo_pc__13_,fe_queue_lo_pc__12_,fe_queue_lo_pc__11_,
  fe_queue_lo_pc__10_,fe_queue_lo_pc__9_,fe_queue_lo_pc__8_,fe_queue_lo_pc__7_,fe_queue_lo_pc__6_,
  fe_queue_lo_pc__5_,fe_queue_lo_pc__4_,fe_queue_lo_pc__3_,fe_queue_lo_pc__2_,
  fe_queue_lo_pc__1_,fe_queue_lo_pc__0_,fe_queue_lo_instr__79_,fe_queue_lo_instr__78_,
  fe_queue_lo_instr__77_,fe_queue_lo_instr__76_,fe_queue_lo_instr__75_,
  fe_queue_lo_instr__74_,fe_queue_lo_instr__73_,fe_queue_lo_instr__72_,
  fe_queue_lo_instr__71_,fe_queue_lo_instr__70_,fe_queue_lo_instr__69_,fe_queue_lo_instr__68_,
  fe_queue_lo_instr__67_,fe_queue_lo_instr__66_,fe_queue_lo_instr__65_,
  fe_queue_lo_instr__64_,fe_queue_lo_instr__63_,fe_queue_lo_instr__62_,fe_queue_lo_instr__61_,
  fe_queue_lo_instr__60_,fe_queue_lo_instr__59_,fe_queue_lo_instr__58_,
  fe_queue_lo_instr__57_,fe_queue_lo_instr__56_,fe_queue_lo_instr__55_,fe_queue_lo_instr__54_,
  fe_queue_lo_instr__53_,fe_queue_lo_instr__52_,fe_queue_lo_instr__51_,
  fe_queue_lo_instr__50_,fe_queue_lo_instr__49_,fe_queue_lo_instr__48_,fe_queue_lo_instr__47_,
  fe_queue_lo_instr__46_,fe_queue_lo_instr__45_,fe_queue_lo_instr__44_,
  fe_queue_lo_instr__43_,fe_queue_lo_instr__42_,fe_queue_lo_instr__41_,fe_queue_lo_instr__40_,
  fe_queue_lo_instr__39_,fe_queue_lo_instr__38_,fe_queue_lo_instr__37_,
  fe_queue_lo_instr__36_,fe_queue_lo_instr__35_,fe_queue_lo_instr__34_,fe_queue_lo_instr__33_,
  fe_queue_lo_instr__32_,fe_queue_lo_instr__31_,fe_queue_lo_instr__30_,
  fe_queue_lo_instr__29_,fe_queue_lo_instr__28_,fe_queue_lo_instr__27_,fe_queue_lo_instr__26_,
  fe_queue_lo_instr__25_,fe_queue_lo_instr__24_,fe_queue_lo_instr__23_,
  fe_queue_lo_instr__22_,fe_queue_lo_instr__21_,fe_queue_lo_instr__20_,fe_queue_lo_instr__19_,
  fe_queue_lo_instr__18_,fe_queue_lo_instr__17_,fe_queue_lo_instr__16_,
  fe_queue_lo_instr__15_,fe_queue_lo_instr__14_,fe_queue_lo_instr__13_,fe_queue_lo_instr__12_,
  fe_queue_lo_instr__11_,fe_queue_lo_instr__10_,fe_queue_lo_instr__9_,
  fe_queue_lo_instr__8_,fe_queue_lo_instr__7_,fe_queue_lo_instr__6_,fe_queue_lo_instr__5_,
  fe_queue_lo_instr__4_,fe_queue_lo_instr__3_,fe_queue_lo_instr__2_,
  fe_queue_lo_instr__1_,fe_queue_lo_instr__0_,fe_queue_lo_msg_type__2_,fe_queue_lo_msg_type__1_,
  fe_queue_lo_msg_type__0_,N600,illegal_instr_lo,N601,N602,N604,N605,N606,N608,N609,
  N610,N612,N613,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,
  N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,
  N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,
  N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,
  N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,
  N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,
  N708,N709,N710,N711,N712,N713,N714;
  wire [6:0] rptr_r,wptr_r,rptr_n,wptr_n,cptr_r,cptr_n,rptr_jmp,wptr_jmp,cptr_jmp;
  wire [3:0] enq,read,deq;
  wire [79:0] queue_instr_n;
  wire [2:0] preissue_entry_sel;
  wire [31:0] \e_0_.instr ,\e_1_.instr ,\e_2_.instr ,\e_3_.instr ,\e_4_.instr ;
  wire [159:0] preissue_instr;
  assign issue_pkt_o[113] = 1'b0;
  assign issue_pkt_o[114] = 1'b0;
  assign empty = rptr_r == wptr_r;
  assign empty_n = rptr_n == wptr_n;
  assign N69 = cptr_r[5:3] == wptr_r[5:3];
  assign N70 = cptr_r[6] ^ wptr_r[6];
  assign read_catchup = { N74, N73, N72, N71 } >= read_cnt_i;
  assign deq_catchup = { N78, N77, N76, N75 } >= cmt_cnt_i;

  bsg_circular_ptr_slots_p128_max_add_p127
  cptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(cptr_jmp),
    .o(cptr_r),
    .n_o(cptr_n)
  );


  bsg_circular_ptr_slots_p128_max_add_p127
  wptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(wptr_jmp),
    .o(wptr_r),
    .n_o(wptr_n)
  );


  bsg_circular_ptr_slots_p128_max_add_p127
  rptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(rptr_jmp),
    .o(rptr_r),
    .n_o(rptr_n)
  );

  assign bypass_preissue = wptr_r == rptr_n;

  bsg_mem_1r1w_00000050_00000008
  preissue_fifo_mem
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(_0_net_),
    .w_addr_i(wptr_r[5:3]),
    .w_data_i(fe_queue_i[134:55]),
    .r_v_i(_2_net_),
    .r_addr_i(rptr_n[5:3]),
    .r_data_o(queue_instr_n)
  );


  bp_be_expander
  \e_0_.expander 
  (
    .cinstr_i({ queue_instr_raw_0__15_, queue_instr_raw_0__14_, queue_instr_raw_0__13_, queue_instr_raw_0__12_, queue_instr_raw_0__11_, queue_instr_raw_0__10_, queue_instr_raw_0__9_, queue_instr_raw_0__8_, queue_instr_raw_0__7_, queue_instr_raw_0__6_, queue_instr_raw_0__5_, queue_instr_raw_0__4_, queue_instr_raw_0__3_, queue_instr_raw_0__2_, queue_instr_raw_0__1_, queue_instr_raw_0__0_ }),
    .instr_o(\e_0_.instr )
  );


  bp_be_expander
  \e_1_.expander 
  (
    .cinstr_i({ queue_instr_raw_1__15_, queue_instr_raw_1__14_, queue_instr_raw_1__13_, queue_instr_raw_1__12_, queue_instr_raw_1__11_, queue_instr_raw_1__10_, queue_instr_raw_1__9_, queue_instr_raw_1__8_, queue_instr_raw_1__7_, queue_instr_raw_1__6_, queue_instr_raw_1__5_, queue_instr_raw_1__4_, queue_instr_raw_1__3_, queue_instr_raw_1__2_, queue_instr_raw_1__1_, queue_instr_raw_1__0_ }),
    .instr_o(\e_1_.instr )
  );


  bp_be_expander
  \e_2_.expander 
  (
    .cinstr_i({ queue_instr_raw_2__15_, queue_instr_raw_2__14_, queue_instr_raw_2__13_, queue_instr_raw_2__12_, queue_instr_raw_2__11_, queue_instr_raw_2__10_, queue_instr_raw_2__9_, queue_instr_raw_2__8_, queue_instr_raw_2__7_, queue_instr_raw_2__6_, queue_instr_raw_2__5_, queue_instr_raw_2__4_, queue_instr_raw_2__3_, queue_instr_raw_2__2_, queue_instr_raw_2__1_, queue_instr_raw_2__0_ }),
    .instr_o(\e_2_.instr )
  );


  bp_be_expander
  \e_3_.expander 
  (
    .cinstr_i({ queue_instr_raw_3__15_, queue_instr_raw_3__14_, queue_instr_raw_3__13_, queue_instr_raw_3__12_, queue_instr_raw_3__11_, queue_instr_raw_3__10_, queue_instr_raw_3__9_, queue_instr_raw_3__8_, queue_instr_raw_3__7_, queue_instr_raw_3__6_, queue_instr_raw_3__5_, queue_instr_raw_3__4_, queue_instr_raw_3__3_, queue_instr_raw_3__2_, queue_instr_raw_3__1_, queue_instr_raw_3__0_ }),
    .instr_o(\e_3_.instr )
  );


  bp_be_expander
  \e_4_.expander 
  (
    .cinstr_i({ queue_instr_raw_4__15_, queue_instr_raw_4__14_, queue_instr_raw_4__13_, queue_instr_raw_4__12_, queue_instr_raw_4__11_, queue_instr_raw_4__10_, queue_instr_raw_4__9_, queue_instr_raw_4__8_, queue_instr_raw_4__7_, queue_instr_raw_4__6_, queue_instr_raw_4__5_, queue_instr_raw_4__4_, queue_instr_raw_4__3_, queue_instr_raw_4__2_, queue_instr_raw_4__1_, queue_instr_raw_4__0_ }),
    .instr_o(\e_4_.instr )
  );

  assign N183 = N178 | N179;
  assign N184 = N173 | N174;
  assign N185 = N180 | N181;
  assign N186 = N183 | N184;
  assign N187 = N185 | N182;
  assign N188 = N186 | N187;
  assign N189 = N171 | N172;
  assign N190 = N175 | N181;
  assign N191 = N189 | N184;
  assign N192 = N190 | N182;
  assign N193 = N191 | N192;
  assign N195 = N194 | N174;
  assign N196 = N189 | N195;
  assign N197 = N196 | N192;
  assign N199 = N194 | N198;
  assign N200 = N189 | N199;
  assign N201 = N200 | N192;
  assign N202 = N183 | N195;
  assign N203 = N202 | N192;
  assign N205 = N186 | N192;
  assign N206 = N171 | N179;
  assign N207 = N206 | N184;
  assign N208 = N207 | N192;
  assign N209 = N206 | N195;
  assign N210 = N209 | N192;
  assign N211 = N206 | N199;
  assign N212 = N211 | N192;
  assign N213 = N173 | N198;
  assign N214 = N206 | N213;
  assign N215 = N214 | N187;
  assign N217 = N189 | N213;
  assign N218 = N217 | N187;
  assign N220 = N191 | N187;
  assign N222 = N207 | N187;
  assign N224 = N178 | N172;
  assign N225 = N224 | N195;
  assign N226 = N225 | N192;
  assign N228 = N224 | N184;
  assign N229 = N228 | N192;
  assign N230 = N228 | N187;
  assign N231 = N224 | N213;
  assign N232 = N231 | N192;
  assign N233 = N231 | N187;
  assign N235 = N171 & N172;
  assign N236 = N235 & N174;
  assign N237 = N172 & N194;
  assign N238 = N174 & N180;
  assign N239 = N237 & N238;
  assign N240 = N171 & N173;
  assign N241 = N240 & N174;
  assign N242 = N173 & N175;
  assign N243 = N178 & N194;
  assign N244 = N243 & N238;
  assign N265 = N246 & N247;
  assign N266 = N248 & N249;
  assign N267 = N250 & N251;
  assign N268 = N252 & N253;
  assign N269 = N254 & N255;
  assign N270 = preissue_pkt_o[15] & N256;
  assign N271 = N257 & N258;
  assign N272 = N259 & N260;
  assign N273 = N261 & N262;
  assign N274 = N263 & N264;
  assign N275 = preissue_pkt_o[5] & preissue_pkt_o[4];
  assign N276 = preissue_pkt_o[3] & preissue_pkt_o[2];
  assign N277 = N265 & N266;
  assign N278 = N267 & N268;
  assign N279 = N269 & N270;
  assign N280 = N271 & N272;
  assign N281 = N273 & N274;
  assign N282 = N275 & N276;
  assign N283 = N277 & N278;
  assign N284 = N279 & N280;
  assign N285 = N281 & N282;
  assign N286 = N283 & N284;
  assign N287 = N286 & N285;
  assign N290 = preissue_pkt_o[24] & N288;
  assign N291 = N290 & N289;
  assign N294 = N292 & N293;
  assign N295 = N294 & preissue_pkt_o[22];
  assign N299 = N296 & N297;
  assign N300 = N299 & N298;
  assign N303 = N301 & preissue_pkt_o[23];
  assign N304 = N303 & N302;
  assign N320 = preissue_pkt_o[32] & N312;
  assign N321 = N313 & N314;
  assign N322 = N315 & N316;
  assign N323 = preissue_pkt_o[8] & N317;
  assign N324 = preissue_pkt_o[6] & N318;
  assign N325 = N319 & preissue_pkt_o[3];
  assign N326 = N320 & N321;
  assign N327 = N322 & N323;
  assign N328 = N324 & N325;
  assign N329 = N326 & N327;
  assign N330 = N328 & preissue_pkt_o[2];
  assign N331 = N329 & N330;
  assign N338 = preissue_pkt_o[33] & N333;
  assign N339 = N334 & N335;
  assign N340 = N336 & N337;
  assign N341 = N338 & N339;
  assign N342 = N341 & N340;
  assign N347 = preissue_pkt_o[33] & N343;
  assign N348 = N344 & N345;
  assign N349 = N346 & preissue_pkt_o[22];
  assign N350 = N347 & N348;
  assign N351 = N350 & N349;
  assign N356 = preissue_pkt_o[33] & N352;
  assign N357 = N353 & N354;
  assign N358 = preissue_pkt_o[23] & N355;
  assign N359 = N356 & N357;
  assign N360 = N359 & N358;
  assign N364 = preissue_pkt_o[33] & N361;
  assign N365 = N362 & N363;
  assign N366 = preissue_pkt_o[23] & preissue_pkt_o[22];
  assign N367 = N364 & N365;
  assign N368 = N367 & N366;
  assign N373 = preissue_pkt_o[33] & N369;
  assign N374 = N370 & preissue_pkt_o[27];
  assign N375 = N371 & N372;
  assign N376 = N373 & N374;
  assign N377 = N376 & N375;
  assign N381 = preissue_pkt_o[33] & N378;
  assign N382 = N379 & preissue_pkt_o[27];
  assign N383 = N380 & preissue_pkt_o[22];
  assign N384 = N381 & N382;
  assign N385 = N384 & N383;
  assign N389 = preissue_pkt_o[33] & N386;
  assign N390 = N387 & preissue_pkt_o[27];
  assign N391 = preissue_pkt_o[23] & N388;
  assign N392 = N389 & N390;
  assign N393 = N392 & N391;
  assign N396 = preissue_pkt_o[33] & N394;
  assign N397 = N395 & preissue_pkt_o[27];
  assign N398 = preissue_pkt_o[23] & preissue_pkt_o[22];
  assign N399 = N396 & N397;
  assign N400 = N399 & N398;
  assign N406 = N401 & N402;
  assign N407 = N403 & N404;
  assign N408 = N405 & preissue_pkt_o[22];
  assign N409 = N406 & N407;
  assign N410 = N409 & N408;
  assign N416 = N411 & N412;
  assign N417 = N413 & preissue_pkt_o[27];
  assign N418 = N414 & N415;
  assign N419 = N416 & N417;
  assign N420 = N419 & N418;
  assign N428 = preissue_pkt_o[33] & preissue_pkt_o[31];
  assign N429 = N421 & N422;
  assign N430 = N423 & N424;
  assign N431 = N425 & N426;
  assign N432 = N428 & N429;
  assign N433 = N430 & N431;
  assign N434 = N432 & N433;
  assign N435 = N434 & N427;
  assign N442 = preissue_pkt_o[33] & preissue_pkt_o[31];
  assign N443 = N436 & preissue_pkt_o[27];
  assign N444 = N437 & N438;
  assign N445 = N439 & N440;
  assign N446 = N442 & N443;
  assign N447 = N444 & N445;
  assign N448 = N446 & N447;
  assign N449 = N448 & N441;
  assign N456 = preissue_pkt_o[33] & preissue_pkt_o[31];
  assign N457 = N450 & N451;
  assign N458 = N452 & N453;
  assign N459 = N454 & N455;
  assign N460 = N456 & N457;
  assign N461 = N458 & N459;
  assign N462 = N460 & N461;
  assign N463 = N462 & preissue_pkt_o[14];
  assign N469 = preissue_pkt_o[33] & preissue_pkt_o[31];
  assign N470 = N464 & preissue_pkt_o[27];
  assign N471 = N465 & N466;
  assign N472 = N467 & N468;
  assign N473 = N469 & N470;
  assign N474 = N471 & N472;
  assign N475 = N473 & N474;
  assign N476 = N475 & preissue_pkt_o[14];
  assign N482 = preissue_pkt_o[33] & N478;
  assign N483 = preissue_pkt_o[30] & N479;
  assign N484 = N480 & N481;
  assign N485 = N482 & N483;
  assign N486 = N485 & N484;
  assign N490 = preissue_pkt_o[33] & N487;
  assign N491 = preissue_pkt_o[30] & N488;
  assign N492 = N489 & preissue_pkt_o[22];
  assign N493 = N490 & N491;
  assign N494 = N493 & N492;
  assign N498 = preissue_pkt_o[33] & N495;
  assign N499 = preissue_pkt_o[30] & N496;
  assign N500 = preissue_pkt_o[23] & N497;
  assign N501 = N498 & N499;
  assign N502 = N501 & N500;
  assign N505 = preissue_pkt_o[33] & N503;
  assign N506 = preissue_pkt_o[30] & N504;
  assign N507 = preissue_pkt_o[23] & preissue_pkt_o[22];
  assign N508 = N505 & N506;
  assign N509 = N508 & N507;
  assign N513 = preissue_pkt_o[33] & N510;
  assign N514 = preissue_pkt_o[30] & preissue_pkt_o[27];
  assign N515 = N511 & N512;
  assign N516 = N513 & N514;
  assign N517 = N516 & N515;
  assign N520 = preissue_pkt_o[33] & N518;
  assign N521 = preissue_pkt_o[30] & preissue_pkt_o[27];
  assign N522 = N519 & preissue_pkt_o[22];
  assign N523 = N520 & N521;
  assign N524 = N523 & N522;
  assign N527 = preissue_pkt_o[33] & N525;
  assign N528 = preissue_pkt_o[30] & preissue_pkt_o[27];
  assign N529 = preissue_pkt_o[23] & N526;
  assign N530 = N527 & N528;
  assign N531 = N530 & N529;
  assign N533 = preissue_pkt_o[33] & N532;
  assign N534 = preissue_pkt_o[30] & preissue_pkt_o[27];
  assign N535 = preissue_pkt_o[23] & preissue_pkt_o[22];
  assign N536 = N533 & N534;
  assign N537 = N536 & N535;
  assign N544 = preissue_pkt_o[33] & preissue_pkt_o[31];
  assign N545 = preissue_pkt_o[30] & N538;
  assign N546 = N539 & N540;
  assign N547 = N541 & N542;
  assign N548 = N544 & N545;
  assign N549 = N546 & N547;
  assign N550 = N548 & N549;
  assign N551 = N550 & N543;
  assign N557 = preissue_pkt_o[33] & preissue_pkt_o[31];
  assign N558 = preissue_pkt_o[30] & preissue_pkt_o[27];
  assign N559 = N552 & N553;
  assign N560 = N554 & N555;
  assign N561 = N557 & N558;
  assign N562 = N559 & N560;
  assign N563 = N561 & N562;
  assign N564 = N563 & N556;
  assign N567 = N566 & preissue_pkt_o[27];
  assign N568 = N567 & preissue_pkt_o[22];
  assign N570 = N569 & preissue_pkt_o[31];
  assign N571 = N570 & preissue_pkt_o[27];
  assign N572 = preissue_pkt_o[31] & preissue_pkt_o[22];
  assign N574 = N573 & preissue_pkt_o[23];
  assign N576 = N575 & preissue_pkt_o[30];
  assign N580 = N577 & N578;
  assign N581 = N580 & N579;
  assign N582 = preissue_pkt_o[31] & preissue_pkt_o[30];
  assign N583 = N582 & preissue_pkt_o[14];
  assign N584 = preissue_pkt_o[31] & preissue_pkt_o[23];
  assign N585 = preissue_pkt_o[31] & preissue_pkt_o[16];
  assign N586 = preissue_pkt_o[31] & preissue_pkt_o[15];

  bsg_dff_reset_en_width_p39
  issue_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(preissue_v),
    .data_i(preissue_pkt_o),
    .data_o({ preissue_pkt_r_irs1_v_, preissue_pkt_r_irs2_v_, preissue_pkt_r_frs1_v_, preissue_pkt_r_frs2_v_, preissue_pkt_r_frs3_v_, issue_pkt_o[205:174], preissue_pkt_r_size__1_, preissue_pkt_r_size__0_ })
  );

  assign bypass_issue = wptr_r[5:3] == rptr_r[5:3];

  bsg_mem_1r1w_000000ae_00000008
  queue_fifo_mem
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(_4_net_),
    .w_addr_i(wptr_r[5:3]),
    .w_data_i(fe_queue_i),
    .r_v_i(_6_net_),
    .r_addr_i(rptr_r[5:3]),
    .r_data_o({ fe_queue_lo_pc__38_, fe_queue_lo_pc__37_, fe_queue_lo_pc__36_, fe_queue_lo_pc__35_, fe_queue_lo_pc__34_, fe_queue_lo_pc__33_, fe_queue_lo_pc__32_, fe_queue_lo_pc__31_, fe_queue_lo_pc__30_, fe_queue_lo_pc__29_, fe_queue_lo_pc__28_, fe_queue_lo_pc__27_, fe_queue_lo_pc__26_, fe_queue_lo_pc__25_, fe_queue_lo_pc__24_, fe_queue_lo_pc__23_, fe_queue_lo_pc__22_, fe_queue_lo_pc__21_, fe_queue_lo_pc__20_, fe_queue_lo_pc__19_, fe_queue_lo_pc__18_, fe_queue_lo_pc__17_, fe_queue_lo_pc__16_, fe_queue_lo_pc__15_, fe_queue_lo_pc__14_, fe_queue_lo_pc__13_, fe_queue_lo_pc__12_, fe_queue_lo_pc__11_, fe_queue_lo_pc__10_, fe_queue_lo_pc__9_, fe_queue_lo_pc__8_, fe_queue_lo_pc__7_, fe_queue_lo_pc__6_, fe_queue_lo_pc__5_, fe_queue_lo_pc__4_, fe_queue_lo_pc__3_, fe_queue_lo_pc__2_, fe_queue_lo_pc__1_, fe_queue_lo_pc__0_, fe_queue_lo_instr__79_, fe_queue_lo_instr__78_, fe_queue_lo_instr__77_, fe_queue_lo_instr__76_, fe_queue_lo_instr__75_, fe_queue_lo_instr__74_, fe_queue_lo_instr__73_, fe_queue_lo_instr__72_, fe_queue_lo_instr__71_, fe_queue_lo_instr__70_, fe_queue_lo_instr__69_, fe_queue_lo_instr__68_, fe_queue_lo_instr__67_, fe_queue_lo_instr__66_, fe_queue_lo_instr__65_, fe_queue_lo_instr__64_, fe_queue_lo_instr__63_, fe_queue_lo_instr__62_, fe_queue_lo_instr__61_, fe_queue_lo_instr__60_, fe_queue_lo_instr__59_, fe_queue_lo_instr__58_, fe_queue_lo_instr__57_, fe_queue_lo_instr__56_, fe_queue_lo_instr__55_, fe_queue_lo_instr__54_, fe_queue_lo_instr__53_, fe_queue_lo_instr__52_, fe_queue_lo_instr__51_, fe_queue_lo_instr__50_, fe_queue_lo_instr__49_, fe_queue_lo_instr__48_, fe_queue_lo_instr__47_, fe_queue_lo_instr__46_, fe_queue_lo_instr__45_, fe_queue_lo_instr__44_, fe_queue_lo_instr__43_, fe_queue_lo_instr__42_, fe_queue_lo_instr__41_, fe_queue_lo_instr__40_, fe_queue_lo_instr__39_, fe_queue_lo_instr__38_, fe_queue_lo_instr__37_, fe_queue_lo_instr__36_, fe_queue_lo_instr__35_, fe_queue_lo_instr__34_, fe_queue_lo_instr__33_, fe_queue_lo_instr__32_, fe_queue_lo_instr__31_, fe_queue_lo_instr__30_, fe_queue_lo_instr__29_, fe_queue_lo_instr__28_, fe_queue_lo_instr__27_, fe_queue_lo_instr__26_, fe_queue_lo_instr__25_, fe_queue_lo_instr__24_, fe_queue_lo_instr__23_, fe_queue_lo_instr__22_, fe_queue_lo_instr__21_, fe_queue_lo_instr__20_, fe_queue_lo_instr__19_, fe_queue_lo_instr__18_, fe_queue_lo_instr__17_, fe_queue_lo_instr__16_, fe_queue_lo_instr__15_, fe_queue_lo_instr__14_, fe_queue_lo_instr__13_, fe_queue_lo_instr__12_, fe_queue_lo_instr__11_, fe_queue_lo_instr__10_, fe_queue_lo_instr__9_, fe_queue_lo_instr__8_, fe_queue_lo_instr__7_, fe_queue_lo_instr__6_, fe_queue_lo_instr__5_, fe_queue_lo_instr__4_, fe_queue_lo_instr__3_, fe_queue_lo_instr__2_, fe_queue_lo_instr__1_, fe_queue_lo_instr__0_, issue_pkt_o[48:0], issue_pkt_o[173:171], fe_queue_lo_msg_type__2_, fe_queue_lo_msg_type__1_, fe_queue_lo_msg_type__0_ })
  );


  bp_be_instr_decoder_00
  instr_decoder
  (
    .preissue_pkt_i({ preissue_pkt_r_irs1_v_, preissue_pkt_r_irs2_v_, preissue_pkt_r_frs1_v_, preissue_pkt_r_frs2_v_, preissue_pkt_r_frs3_v_, issue_pkt_o[205:174], preissue_pkt_r_size__1_, preissue_pkt_r_size__0_ }),
    .decode_info_i(decode_info_i),
    .decode_o(issue_pkt_o[168:115]),
    .illegal_instr_o(illegal_instr_lo),
    .ecall_m_o(issue_pkt_o[256]),
    .ecall_s_o(issue_pkt_o[255]),
    .ecall_u_o(issue_pkt_o[254]),
    .ebreak_o(issue_pkt_o[253]),
    .dbreak_o(issue_pkt_o[252]),
    .dret_o(issue_pkt_o[251]),
    .mret_o(issue_pkt_o[250]),
    .sret_o(issue_pkt_o[249]),
    .wfi_o(issue_pkt_o[248]),
    .sfence_vma_o(issue_pkt_o[247]),
    .fencei_o(issue_pkt_o[246]),
    .csrw_o(issue_pkt_o[245]),
    .imm_o(issue_pkt_o[112:49])
  );

  assign N601 = fe_queue_lo_msg_type__1_ | fe_queue_lo_msg_type__2_;
  assign N602 = fe_queue_lo_msg_type__0_ | N601;
  assign issue_pkt_o[261] = ~N602;
  assign N604 = ~fe_queue_lo_msg_type__1_;
  assign N605 = N604 | fe_queue_lo_msg_type__2_;
  assign N606 = fe_queue_lo_msg_type__0_ | N605;
  assign issue_pkt_o[260] = ~N606;
  assign N608 = ~fe_queue_lo_msg_type__0_;
  assign N609 = fe_queue_lo_msg_type__1_ | fe_queue_lo_msg_type__2_;
  assign N610 = N608 | N609;
  assign issue_pkt_o[259] = ~N610;
  assign N612 = N604 | fe_queue_lo_msg_type__2_;
  assign N613 = N608 | N612;
  assign issue_pkt_o[258] = ~N613;
  assign N615 = ~fe_queue_lo_msg_type__2_;
  assign N616 = fe_queue_lo_msg_type__1_ | N615;
  assign N617 = fe_queue_lo_msg_type__0_ | N616;
  assign N618 = ~N617;
  assign N619 = fe_queue_lo_msg_type__1_ | N615;
  assign N620 = fe_queue_lo_msg_type__0_ | N619;
  assign N621 = ~N620;
  assign N622 = ~preissue_size_0__0_;
  assign N623 = N622 | preissue_size_0__1_;
  assign N624 = ~N623;
  assign N625 = ~preissue_size_1__0_;
  assign N626 = N625 | preissue_size_1__1_;
  assign N627 = ~N626;
  assign N628 = ~preissue_size_2__0_;
  assign N629 = N628 | preissue_size_2__1_;
  assign N630 = ~N629;
  assign N631 = ~preissue_size_3__0_;
  assign N632 = N631 | preissue_size_3__1_;
  assign N633 = ~N632;
  assign N634 = ~preissue_size_4__0_;
  assign N635 = N634 | preissue_size_4__1_;
  assign N636 = ~N635;
  assign { N78, N77, N76, N75 } = cptr_r[2:0] + cmt_size_i;
  assign { N74, N73, N72, N71 } = rptr_r[2:0] + read_size_i;
  assign issue_pkt_o[244:206] = { fe_queue_lo_pc__38_, fe_queue_lo_pc__37_, fe_queue_lo_pc__36_, fe_queue_lo_pc__35_, fe_queue_lo_pc__34_, fe_queue_lo_pc__33_, fe_queue_lo_pc__32_, fe_queue_lo_pc__31_, fe_queue_lo_pc__30_, fe_queue_lo_pc__29_, fe_queue_lo_pc__28_, fe_queue_lo_pc__27_, fe_queue_lo_pc__26_, fe_queue_lo_pc__25_, fe_queue_lo_pc__24_, fe_queue_lo_pc__23_, fe_queue_lo_pc__22_, fe_queue_lo_pc__21_, fe_queue_lo_pc__20_, fe_queue_lo_pc__19_, fe_queue_lo_pc__18_, fe_queue_lo_pc__17_, fe_queue_lo_pc__16_, fe_queue_lo_pc__15_, fe_queue_lo_pc__14_, fe_queue_lo_pc__13_, fe_queue_lo_pc__12_, fe_queue_lo_pc__11_, fe_queue_lo_pc__10_, fe_queue_lo_pc__9_, fe_queue_lo_pc__8_, fe_queue_lo_pc__7_, fe_queue_lo_pc__6_, fe_queue_lo_pc__5_, fe_queue_lo_pc__4_, fe_queue_lo_pc__3_, fe_queue_lo_pc__2_, fe_queue_lo_pc__1_, fe_queue_lo_pc__0_ } + { rptr_r[2:0], 1'b0 };
  assign { N152, N151, N150, N149, N148, N147, N146 } = 1'b0 - cptr_r;
  assign { N145, N144, N143, N142, N141, N140, N139 } = 1'b0 - wptr_r;
  assign { N120, N119, N118, N117, N116, N115, N114 } = 1'b0 - rptr_r;
  assign { N107, N106, N105, N104 } = { 1'b1, 1'b0, 1'b0, 1'b0 } - cptr_r[2:0];
  assign { N96, N95, N94, N93 } = { 1'b1, 1'b0, 1'b0, 1'b0 } - rptr_r[2:0];
  assign { N128, N127, N126, N125, N124, N123, N122 } = cptr_r - rptr_r;
  assign { N135, N134, N133, N132, N131, N130, N129 } = { N128, N127, N126, N125, N124, N123, N122 } + deq;
  assign { N85, N84, N83, N82 } = { 1'b1, 1'b0, 1'b0, 1'b0 } - wptr_r[2:0];
  assign N159 = N0 & N1 & N2;
  assign N0 = ~preissue_entry_sel[2];
  assign N1 = ~preissue_entry_sel[0];
  assign N2 = ~preissue_entry_sel[1];
  assign N160 = preissue_entry_sel[0] & N3;
  assign N3 = ~preissue_entry_sel[1];
  assign N161 = N4 & preissue_entry_sel[1];
  assign N4 = ~preissue_entry_sel[0];
  assign N162 = preissue_entry_sel[0] & preissue_entry_sel[1];
  assign N163 = N5 & N6 & N7;
  assign N5 = ~preissue_entry_sel[2];
  assign N6 = ~preissue_entry_sel[0];
  assign N7 = ~preissue_entry_sel[1];
  assign N164 = preissue_entry_sel[0] & N8;
  assign N8 = ~preissue_entry_sel[1];
  assign N165 = N9 & preissue_entry_sel[1];
  assign N9 = ~preissue_entry_sel[0];
  assign N166 = preissue_entry_sel[0] & preissue_entry_sel[1];
  assign N167 = N10 & N11 & N12;
  assign N10 = ~preissue_entry_sel[2];
  assign N11 = ~preissue_entry_sel[0];
  assign N12 = ~preissue_entry_sel[1];
  assign N168 = preissue_entry_sel[0] & N13;
  assign N13 = ~preissue_entry_sel[1];
  assign N169 = N14 & preissue_entry_sel[1];
  assign N14 = ~preissue_entry_sel[0];
  assign N170 = preissue_entry_sel[0] & preissue_entry_sel[1];
  assign { N89, N88, N87, N86 } = (N15)? { N85, N84, N83, N82 } : 
                                  (N16)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = 1'b1;
  assign N16 = N81;
  assign enq = (N17)? { N89, N88, N87, N86 } : 
               (N18)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N17 = ack;
  assign N18 = N79;
  assign { N100, N99, N98, N97 } = (N19)? { N96, N95, N94, N93 } : 
                                   (N20)? read_size_i : 1'b0;
  assign N19 = read_catchup;
  assign N20 = N92;
  assign read = (N21)? { N100, N99, N98, N97 } : 
                (N22)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N21 = read_i;
  assign N22 = N90;
  assign { N111, N110, N109, N108 } = (N23)? { N107, N106, N105, N104 } : 
                                      (N24)? cmt_size_i : 1'b0;
  assign N23 = deq_catchup;
  assign N24 = N103;
  assign deq = (N25)? { N111, N110, N109, N108 } : 
               (N26)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N25 = cmt_i;
  assign N26 = N101;
  assign rptr_jmp = (N27)? { N120, N119, N118, N117, N116, N115, N114 } : 
                    (N137)? { N135, N134, N133, N132, N131, N130, N129 } : 
                    (N113)? { 1'b0, 1'b0, 1'b0, read } : 1'b0;
  assign N27 = clr_i;
  assign wptr_jmp = (N27)? { N145, N144, N143, N142, N141, N140, N139 } : 
                    (N28)? { 1'b0, 1'b0, 1'b0, enq } : 1'b0;
  assign N28 = N138;
  assign cptr_jmp = (N27)? { N152, N151, N150, N149, N148, N147, N146 } : 
                    (N28)? { 1'b0, 1'b0, 1'b0, deq } : 1'b0;
  assign preissue_entry_sel = (N29)? wptr_r[2:0] : 
                              (N30)? rptr_n[2:0] : 1'b0;
  assign N29 = bypass_preissue;
  assign N30 = N153;
  assign { queue_instr_raw_4__15_, queue_instr_raw_4__14_, queue_instr_raw_4__13_, queue_instr_raw_4__12_, queue_instr_raw_4__11_, queue_instr_raw_4__10_, queue_instr_raw_4__9_, queue_instr_raw_4__8_, queue_instr_raw_4__7_, queue_instr_raw_4__6_, queue_instr_raw_4__5_, queue_instr_raw_4__4_, queue_instr_raw_4__3_, queue_instr_raw_4__2_, queue_instr_raw_4__1_, queue_instr_raw_4__0_, queue_instr_raw_3__15_, queue_instr_raw_3__14_, queue_instr_raw_3__13_, queue_instr_raw_3__12_, queue_instr_raw_3__11_, queue_instr_raw_3__10_, queue_instr_raw_3__9_, queue_instr_raw_3__8_, queue_instr_raw_3__7_, queue_instr_raw_3__6_, queue_instr_raw_3__5_, queue_instr_raw_3__4_, queue_instr_raw_3__3_, queue_instr_raw_3__2_, queue_instr_raw_3__1_, queue_instr_raw_3__0_, queue_instr_raw_2__15_, queue_instr_raw_2__14_, queue_instr_raw_2__13_, queue_instr_raw_2__12_, queue_instr_raw_2__11_, queue_instr_raw_2__10_, queue_instr_raw_2__9_, queue_instr_raw_2__8_, queue_instr_raw_2__7_, queue_instr_raw_2__6_, queue_instr_raw_2__5_, queue_instr_raw_2__4_, queue_instr_raw_2__3_, queue_instr_raw_2__2_, queue_instr_raw_2__1_, queue_instr_raw_2__0_, queue_instr_raw_1__15_, queue_instr_raw_1__14_, queue_instr_raw_1__13_, queue_instr_raw_1__12_, queue_instr_raw_1__11_, queue_instr_raw_1__10_, queue_instr_raw_1__9_, queue_instr_raw_1__8_, queue_instr_raw_1__7_, queue_instr_raw_1__6_, queue_instr_raw_1__5_, queue_instr_raw_1__4_, queue_instr_raw_1__3_, queue_instr_raw_1__2_, queue_instr_raw_1__1_, queue_instr_raw_1__0_, queue_instr_raw_0__15_, queue_instr_raw_0__14_, queue_instr_raw_0__13_, queue_instr_raw_0__12_, queue_instr_raw_0__11_, queue_instr_raw_0__10_, queue_instr_raw_0__9_, queue_instr_raw_0__8_, queue_instr_raw_0__7_, queue_instr_raw_0__6_, queue_instr_raw_0__5_, queue_instr_raw_0__4_, queue_instr_raw_0__3_, queue_instr_raw_0__2_, queue_instr_raw_0__1_, queue_instr_raw_0__0_ } = (N29)? fe_queue_i[134:55] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (N30)? queue_instr_n : 1'b0;
  assign preissue_size_0__1_ = ~preissue_size_0__0_;
  assign preissue_instr[31:0] = (N31)? \e_0_.instr  : 
                                (N32)? { queue_instr_raw_1__15_, queue_instr_raw_1__14_, queue_instr_raw_1__13_, queue_instr_raw_1__12_, queue_instr_raw_1__11_, queue_instr_raw_1__10_, queue_instr_raw_1__9_, queue_instr_raw_1__8_, queue_instr_raw_1__7_, queue_instr_raw_1__6_, queue_instr_raw_1__5_, queue_instr_raw_1__4_, queue_instr_raw_1__3_, queue_instr_raw_1__2_, queue_instr_raw_1__1_, queue_instr_raw_1__0_, queue_instr_raw_0__15_, queue_instr_raw_0__14_, queue_instr_raw_0__13_, queue_instr_raw_0__12_, queue_instr_raw_0__11_, queue_instr_raw_0__10_, queue_instr_raw_0__9_, queue_instr_raw_0__8_, queue_instr_raw_0__7_, queue_instr_raw_0__6_, queue_instr_raw_0__5_, queue_instr_raw_0__4_, queue_instr_raw_0__3_, queue_instr_raw_0__2_, queue_instr_raw_0__1_, queue_instr_raw_0__0_ } : 1'b0;
  assign N31 = N624;
  assign N32 = N623;
  assign preissue_size_1__1_ = ~preissue_size_1__0_;
  assign preissue_instr[63:32] = (N33)? \e_1_.instr  : 
                                 (N34)? { queue_instr_raw_2__15_, queue_instr_raw_2__14_, queue_instr_raw_2__13_, queue_instr_raw_2__12_, queue_instr_raw_2__11_, queue_instr_raw_2__10_, queue_instr_raw_2__9_, queue_instr_raw_2__8_, queue_instr_raw_2__7_, queue_instr_raw_2__6_, queue_instr_raw_2__5_, queue_instr_raw_2__4_, queue_instr_raw_2__3_, queue_instr_raw_2__2_, queue_instr_raw_2__1_, queue_instr_raw_2__0_, queue_instr_raw_1__15_, queue_instr_raw_1__14_, queue_instr_raw_1__13_, queue_instr_raw_1__12_, queue_instr_raw_1__11_, queue_instr_raw_1__10_, queue_instr_raw_1__9_, queue_instr_raw_1__8_, queue_instr_raw_1__7_, queue_instr_raw_1__6_, queue_instr_raw_1__5_, queue_instr_raw_1__4_, queue_instr_raw_1__3_, queue_instr_raw_1__2_, queue_instr_raw_1__1_, queue_instr_raw_1__0_ } : 1'b0;
  assign N33 = N627;
  assign N34 = N626;
  assign preissue_size_2__1_ = ~preissue_size_2__0_;
  assign preissue_instr[95:64] = (N35)? \e_2_.instr  : 
                                 (N36)? { queue_instr_raw_3__15_, queue_instr_raw_3__14_, queue_instr_raw_3__13_, queue_instr_raw_3__12_, queue_instr_raw_3__11_, queue_instr_raw_3__10_, queue_instr_raw_3__9_, queue_instr_raw_3__8_, queue_instr_raw_3__7_, queue_instr_raw_3__6_, queue_instr_raw_3__5_, queue_instr_raw_3__4_, queue_instr_raw_3__3_, queue_instr_raw_3__2_, queue_instr_raw_3__1_, queue_instr_raw_3__0_, queue_instr_raw_2__15_, queue_instr_raw_2__14_, queue_instr_raw_2__13_, queue_instr_raw_2__12_, queue_instr_raw_2__11_, queue_instr_raw_2__10_, queue_instr_raw_2__9_, queue_instr_raw_2__8_, queue_instr_raw_2__7_, queue_instr_raw_2__6_, queue_instr_raw_2__5_, queue_instr_raw_2__4_, queue_instr_raw_2__3_, queue_instr_raw_2__2_, queue_instr_raw_2__1_, queue_instr_raw_2__0_ } : 1'b0;
  assign N35 = N630;
  assign N36 = N629;
  assign preissue_size_3__1_ = ~preissue_size_3__0_;
  assign preissue_instr[127:96] = (N37)? \e_3_.instr  : 
                                  (N38)? { queue_instr_raw_4__15_, queue_instr_raw_4__14_, queue_instr_raw_4__13_, queue_instr_raw_4__12_, queue_instr_raw_4__11_, queue_instr_raw_4__10_, queue_instr_raw_4__9_, queue_instr_raw_4__8_, queue_instr_raw_4__7_, queue_instr_raw_4__6_, queue_instr_raw_4__5_, queue_instr_raw_4__4_, queue_instr_raw_4__3_, queue_instr_raw_4__2_, queue_instr_raw_4__1_, queue_instr_raw_4__0_, queue_instr_raw_3__15_, queue_instr_raw_3__14_, queue_instr_raw_3__13_, queue_instr_raw_3__12_, queue_instr_raw_3__11_, queue_instr_raw_3__10_, queue_instr_raw_3__9_, queue_instr_raw_3__8_, queue_instr_raw_3__7_, queue_instr_raw_3__6_, queue_instr_raw_3__5_, queue_instr_raw_3__4_, queue_instr_raw_3__3_, queue_instr_raw_3__2_, queue_instr_raw_3__1_, queue_instr_raw_3__0_ } : 1'b0;
  assign N37 = N633;
  assign N38 = N632;
  assign preissue_size_4__1_ = ~preissue_size_4__0_;
  assign preissue_instr[159:128] = (N39)? \e_4_.instr  : 
                                   (N40)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, queue_instr_raw_4__15_, queue_instr_raw_4__14_, queue_instr_raw_4__13_, queue_instr_raw_4__12_, queue_instr_raw_4__11_, queue_instr_raw_4__10_, queue_instr_raw_4__9_, queue_instr_raw_4__8_, queue_instr_raw_4__7_, queue_instr_raw_4__6_, queue_instr_raw_4__5_, queue_instr_raw_4__4_, queue_instr_raw_4__3_, queue_instr_raw_4__2_, queue_instr_raw_4__1_, queue_instr_raw_4__0_ } : 1'b0;
  assign N39 = N636;
  assign N40 = N635;
  assign { N308, N307 } = (N41)? { preissue_v, preissue_v } : 
                          (N306)? { 1'b0, 1'b0 } : 1'b0;
  assign N41 = N305;
  assign { N311, N310 } = (N42)? { N308, N307 } : 
                          (N309)? { 1'b0, 1'b0 } : 1'b0;
  assign N42 = N287;
  assign N590 = (N43)? preissue_v : 
                (N589)? 1'b0 : 1'b0;
  assign N43 = N587;
  assign N591 = (N44)? preissue_v : 
                (N45)? 1'b0 : 
                (N43)? preissue_v : 1'b0;
  assign N44 = N477;
  assign N45 = N565;
  assign N594 = (N45)? preissue_v : 
                (N593)? 1'b0 : 1'b0;
  assign { N597, N596, N595 } = (N46)? { N594, N591, N590 } : 
                                (N332)? { 1'b0, preissue_v, preissue_v } : 1'b0;
  assign N46 = N331;
  assign preissue_pkt_o[34] = (N47)? preissue_v : 
                              (N599)? 1'b0 : 1'b0;
  assign N47 = N234;
  assign preissue_pkt_o[38:35] = (N48)? { preissue_v, 1'b0, 1'b0, 1'b0 } : 
                                 (N49)? { preissue_v, preissue_v, 1'b0, 1'b0 } : 
                                 (N50)? { N311, N310, 1'b0, 1'b0 } : 
                                 (N51)? { preissue_v, 1'b0, 1'b0, 1'b0 } : 
                                 (N52)? { preissue_v, 1'b0, 1'b0, preissue_v } : 
                                 (N53)? { N597, 1'b0, N596, N595 } : 
                                 (N47)? { 1'b0, 1'b0, preissue_v, preissue_v } : 
                                 (N54)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N48 = N204;
  assign N49 = N216;
  assign N50 = N219;
  assign N51 = N221;
  assign N52 = N223;
  assign N53 = N227;
  assign N54 = N245;
  assign issue_pkt_o[170:169] = (N55)? { preissue_pkt_r_size__1_, preissue_pkt_r_size__0_ } : 
                                (N600)? { 1'b1, 1'b1 } : 1'b0;
  assign N55 = issue_pkt_o[262];
  assign preissue_pkt_o[0] = (N56)? preissue_size_0__0_ : 
                             (N57)? preissue_size_1__0_ : 
                             (N58)? preissue_size_2__0_ : 
                             (N59)? preissue_size_3__0_ : 
                             (N60)? preissue_size_4__0_ : 1'b0;
  assign N56 = N159;
  assign N57 = N160;
  assign N58 = N161;
  assign N59 = N162;
  assign N60 = preissue_entry_sel[2];
  assign preissue_pkt_o[1] = (N56)? preissue_size_0__1_ : 
                             (N57)? preissue_size_1__1_ : 
                             (N58)? preissue_size_2__1_ : 
                             (N59)? preissue_size_3__1_ : 
                             (N60)? preissue_size_4__1_ : 1'b0;
  assign preissue_pkt_o[2] = (N61)? preissue_instr[0] : 
                             (N62)? preissue_instr[32] : 
                             (N63)? preissue_instr[64] : 
                             (N64)? preissue_instr[96] : 
                             (N60)? preissue_instr[128] : 1'b0;
  assign N61 = N163;
  assign N62 = N164;
  assign N63 = N165;
  assign N64 = N166;
  assign N177 = (N65)? preissue_instr[0] : 
                (N66)? preissue_instr[32] : 
                (N67)? preissue_instr[64] : 
                (N68)? preissue_instr[96] : 
                (N60)? preissue_instr[128] : 1'b0;
  assign N65 = N167;
  assign N66 = N168;
  assign N67 = N169;
  assign N68 = N170;
  assign preissue_pkt_o[3] = (N61)? preissue_instr[1] : 
                             (N62)? preissue_instr[33] : 
                             (N63)? preissue_instr[65] : 
                             (N64)? preissue_instr[97] : 
                             (N60)? preissue_instr[129] : 1'b0;
  assign N176 = (N65)? preissue_instr[1] : 
                (N66)? preissue_instr[33] : 
                (N67)? preissue_instr[65] : 
                (N68)? preissue_instr[97] : 
                (N60)? preissue_instr[129] : 1'b0;
  assign preissue_pkt_o[4] = (N61)? preissue_instr[2] : 
                             (N62)? preissue_instr[34] : 
                             (N63)? preissue_instr[66] : 
                             (N64)? preissue_instr[98] : 
                             (N60)? preissue_instr[130] : 1'b0;
  assign N175 = (N65)? preissue_instr[2] : 
                (N66)? preissue_instr[34] : 
                (N67)? preissue_instr[66] : 
                (N68)? preissue_instr[98] : 
                (N60)? preissue_instr[130] : 1'b0;
  assign preissue_pkt_o[5] = (N61)? preissue_instr[3] : 
                             (N62)? preissue_instr[35] : 
                             (N63)? preissue_instr[67] : 
                             (N64)? preissue_instr[99] : 
                             (N60)? preissue_instr[131] : 1'b0;
  assign N174 = (N65)? preissue_instr[3] : 
                (N66)? preissue_instr[35] : 
                (N67)? preissue_instr[67] : 
                (N68)? preissue_instr[99] : 
                (N60)? preissue_instr[131] : 1'b0;
  assign preissue_pkt_o[6] = (N61)? preissue_instr[4] : 
                             (N62)? preissue_instr[36] : 
                             (N63)? preissue_instr[68] : 
                             (N64)? preissue_instr[100] : 
                             (N60)? preissue_instr[132] : 1'b0;
  assign N173 = (N65)? preissue_instr[4] : 
                (N66)? preissue_instr[36] : 
                (N67)? preissue_instr[68] : 
                (N68)? preissue_instr[100] : 
                (N60)? preissue_instr[132] : 1'b0;
  assign preissue_pkt_o[7] = (N61)? preissue_instr[5] : 
                             (N62)? preissue_instr[37] : 
                             (N63)? preissue_instr[69] : 
                             (N64)? preissue_instr[101] : 
                             (N60)? preissue_instr[133] : 1'b0;
  assign N172 = (N65)? preissue_instr[5] : 
                (N66)? preissue_instr[37] : 
                (N67)? preissue_instr[69] : 
                (N68)? preissue_instr[101] : 
                (N60)? preissue_instr[133] : 1'b0;
  assign preissue_pkt_o[8] = (N61)? preissue_instr[6] : 
                             (N62)? preissue_instr[38] : 
                             (N63)? preissue_instr[70] : 
                             (N64)? preissue_instr[102] : 
                             (N60)? preissue_instr[134] : 1'b0;
  assign N171 = (N65)? preissue_instr[6] : 
                (N66)? preissue_instr[38] : 
                (N67)? preissue_instr[70] : 
                (N68)? preissue_instr[102] : 
                (N60)? preissue_instr[134] : 1'b0;
  assign preissue_pkt_o[9] = (N61)? preissue_instr[7] : 
                             (N62)? preissue_instr[39] : 
                             (N63)? preissue_instr[71] : 
                             (N64)? preissue_instr[103] : 
                             (N60)? preissue_instr[135] : 1'b0;
  assign preissue_pkt_o[10] = (N61)? preissue_instr[8] : 
                              (N62)? preissue_instr[40] : 
                              (N63)? preissue_instr[72] : 
                              (N64)? preissue_instr[104] : 
                              (N60)? preissue_instr[136] : 1'b0;
  assign preissue_pkt_o[11] = (N61)? preissue_instr[9] : 
                              (N62)? preissue_instr[41] : 
                              (N63)? preissue_instr[73] : 
                              (N64)? preissue_instr[105] : 
                              (N60)? preissue_instr[137] : 1'b0;
  assign preissue_pkt_o[12] = (N61)? preissue_instr[10] : 
                              (N62)? preissue_instr[42] : 
                              (N63)? preissue_instr[74] : 
                              (N64)? preissue_instr[106] : 
                              (N60)? preissue_instr[138] : 1'b0;
  assign preissue_pkt_o[13] = (N61)? preissue_instr[11] : 
                              (N62)? preissue_instr[43] : 
                              (N63)? preissue_instr[75] : 
                              (N64)? preissue_instr[107] : 
                              (N60)? preissue_instr[139] : 1'b0;
  assign preissue_pkt_o[14] = (N61)? preissue_instr[12] : 
                              (N62)? preissue_instr[44] : 
                              (N63)? preissue_instr[76] : 
                              (N64)? preissue_instr[108] : 
                              (N60)? preissue_instr[140] : 1'b0;
  assign preissue_pkt_o[15] = (N61)? preissue_instr[13] : 
                              (N62)? preissue_instr[45] : 
                              (N63)? preissue_instr[77] : 
                              (N64)? preissue_instr[109] : 
                              (N60)? preissue_instr[141] : 1'b0;
  assign preissue_pkt_o[16] = (N61)? preissue_instr[14] : 
                              (N62)? preissue_instr[46] : 
                              (N63)? preissue_instr[78] : 
                              (N64)? preissue_instr[110] : 
                              (N60)? preissue_instr[142] : 1'b0;
  assign preissue_pkt_o[17] = (N61)? preissue_instr[15] : 
                              (N62)? preissue_instr[47] : 
                              (N63)? preissue_instr[79] : 
                              (N64)? preissue_instr[111] : 
                              (N60)? preissue_instr[143] : 1'b0;
  assign preissue_pkt_o[18] = (N61)? preissue_instr[16] : 
                              (N62)? preissue_instr[48] : 
                              (N63)? preissue_instr[80] : 
                              (N64)? preissue_instr[112] : 
                              (N60)? preissue_instr[144] : 1'b0;
  assign preissue_pkt_o[19] = (N61)? preissue_instr[17] : 
                              (N62)? preissue_instr[49] : 
                              (N63)? preissue_instr[81] : 
                              (N64)? preissue_instr[113] : 
                              (N60)? preissue_instr[145] : 1'b0;
  assign preissue_pkt_o[20] = (N61)? preissue_instr[18] : 
                              (N62)? preissue_instr[50] : 
                              (N63)? preissue_instr[82] : 
                              (N64)? preissue_instr[114] : 
                              (N60)? preissue_instr[146] : 1'b0;
  assign preissue_pkt_o[21] = (N61)? preissue_instr[19] : 
                              (N62)? preissue_instr[51] : 
                              (N63)? preissue_instr[83] : 
                              (N64)? preissue_instr[115] : 
                              (N60)? preissue_instr[147] : 1'b0;
  assign preissue_pkt_o[22] = (N61)? preissue_instr[20] : 
                              (N62)? preissue_instr[52] : 
                              (N63)? preissue_instr[84] : 
                              (N64)? preissue_instr[116] : 
                              (N60)? preissue_instr[148] : 1'b0;
  assign preissue_pkt_o[23] = (N61)? preissue_instr[21] : 
                              (N62)? preissue_instr[53] : 
                              (N63)? preissue_instr[85] : 
                              (N64)? preissue_instr[117] : 
                              (N60)? preissue_instr[149] : 1'b0;
  assign preissue_pkt_o[24] = (N61)? preissue_instr[22] : 
                              (N62)? preissue_instr[54] : 
                              (N63)? preissue_instr[86] : 
                              (N64)? preissue_instr[118] : 
                              (N60)? preissue_instr[150] : 1'b0;
  assign preissue_pkt_o[25] = (N61)? preissue_instr[23] : 
                              (N62)? preissue_instr[55] : 
                              (N63)? preissue_instr[87] : 
                              (N64)? preissue_instr[119] : 
                              (N60)? preissue_instr[151] : 1'b0;
  assign preissue_pkt_o[26] = (N61)? preissue_instr[24] : 
                              (N62)? preissue_instr[56] : 
                              (N63)? preissue_instr[88] : 
                              (N64)? preissue_instr[120] : 
                              (N60)? preissue_instr[152] : 1'b0;
  assign preissue_pkt_o[27] = (N61)? preissue_instr[25] : 
                              (N62)? preissue_instr[57] : 
                              (N63)? preissue_instr[89] : 
                              (N64)? preissue_instr[121] : 
                              (N60)? preissue_instr[153] : 1'b0;
  assign preissue_pkt_o[28] = (N61)? preissue_instr[26] : 
                              (N62)? preissue_instr[58] : 
                              (N63)? preissue_instr[90] : 
                              (N64)? preissue_instr[122] : 
                              (N60)? preissue_instr[154] : 1'b0;
  assign preissue_pkt_o[29] = (N61)? preissue_instr[27] : 
                              (N62)? preissue_instr[59] : 
                              (N63)? preissue_instr[91] : 
                              (N64)? preissue_instr[123] : 
                              (N60)? preissue_instr[155] : 1'b0;
  assign preissue_pkt_o[30] = (N61)? preissue_instr[28] : 
                              (N62)? preissue_instr[60] : 
                              (N63)? preissue_instr[92] : 
                              (N64)? preissue_instr[124] : 
                              (N60)? preissue_instr[156] : 1'b0;
  assign preissue_pkt_o[31] = (N61)? preissue_instr[29] : 
                              (N62)? preissue_instr[61] : 
                              (N63)? preissue_instr[93] : 
                              (N64)? preissue_instr[125] : 
                              (N60)? preissue_instr[157] : 1'b0;
  assign preissue_pkt_o[32] = (N61)? preissue_instr[30] : 
                              (N62)? preissue_instr[62] : 
                              (N63)? preissue_instr[94] : 
                              (N64)? preissue_instr[126] : 
                              (N60)? preissue_instr[158] : 1'b0;
  assign preissue_pkt_o[33] = (N61)? preissue_instr[31] : 
                              (N62)? preissue_instr[63] : 
                              (N63)? preissue_instr[95] : 
                              (N64)? preissue_instr[127] : 
                              (N60)? preissue_instr[159] : 1'b0;
  assign ack = fe_queue_ready_and_o & fe_queue_v_i;
  assign full = N69 & N70;
  assign N79 = ~ack;
  assign N80 = ack;
  assign N81 = ~1'b1;
  assign N90 = ~read_i;
  assign N91 = read_i;
  assign N92 = ~read_catchup;
  assign N101 = ~cmt_i;
  assign N102 = cmt_i;
  assign N103 = ~deq_catchup;
  assign N112 = roll_i | clr_i;
  assign N113 = ~N112;
  assign N121 = N137;
  assign N136 = ~clr_i;
  assign N137 = roll_i & N136;
  assign N138 = ~clr_i;
  assign preissue_v = N642 | N646;
  assign N642 = N641 | roll_i;
  assign N641 = N639 & N640;
  assign N639 = N638 | read[0];
  assign N638 = N637 | read[1];
  assign N637 = read[3] | read[2];
  assign N640 = ~empty_n;
  assign N646 = N645 & empty;
  assign N645 = N644 | enq[0];
  assign N644 = N643 | enq[1];
  assign N643 = enq[3] | enq[2];
  assign _2_net_ = ~bypass_preissue;
  assign _0_net_ = N648 | enq[0];
  assign N648 = N647 | enq[1];
  assign N647 = enq[3] | enq[2];
  assign N153 = ~bypass_preissue;
  assign N154 = ~N649;
  assign N649 = queue_instr_raw_0__1_ & queue_instr_raw_0__0_;
  assign preissue_size_0__0_ = N154;
  assign N155 = ~N650;
  assign N650 = queue_instr_raw_1__1_ & queue_instr_raw_1__0_;
  assign preissue_size_1__0_ = N155;
  assign N156 = ~N651;
  assign N651 = queue_instr_raw_2__1_ & queue_instr_raw_2__0_;
  assign preissue_size_2__0_ = N156;
  assign N157 = ~N652;
  assign N652 = queue_instr_raw_3__1_ & queue_instr_raw_3__0_;
  assign preissue_size_3__0_ = N157;
  assign N158 = ~N653;
  assign N653 = queue_instr_raw_4__1_ & queue_instr_raw_4__0_;
  assign preissue_size_4__0_ = N158;
  assign N178 = ~N171;
  assign N179 = ~N172;
  assign N180 = ~N175;
  assign N181 = ~N176;
  assign N182 = ~N177;
  assign N194 = ~N173;
  assign N198 = ~N174;
  assign N204 = N660 | N661;
  assign N660 = N658 | N659;
  assign N658 = N656 | N657;
  assign N656 = N654 | N655;
  assign N654 = ~N188;
  assign N655 = ~N193;
  assign N657 = ~N197;
  assign N659 = ~N201;
  assign N661 = ~N203;
  assign N216 = N668 | N669;
  assign N668 = N666 | N667;
  assign N666 = N664 | N665;
  assign N664 = N662 | N663;
  assign N662 = ~N205;
  assign N663 = ~N208;
  assign N665 = ~N210;
  assign N667 = ~N212;
  assign N669 = ~N215;
  assign N219 = ~N218;
  assign N221 = ~N220;
  assign N223 = ~N222;
  assign N227 = ~N226;
  assign N234 = N674 | N675;
  assign N674 = N672 | N673;
  assign N672 = N670 | N671;
  assign N670 = ~N229;
  assign N671 = ~N230;
  assign N673 = ~N232;
  assign N675 = ~N233;
  assign N245 = N181 | N680;
  assign N680 = N182 | N679;
  assign N679 = N236 | N678;
  assign N678 = N239 | N677;
  assign N677 = N241 | N676;
  assign N676 = N242 | N244;
  assign N246 = ~preissue_pkt_o[33];
  assign N247 = ~preissue_pkt_o[32];
  assign N248 = ~preissue_pkt_o[31];
  assign N249 = ~preissue_pkt_o[30];
  assign N250 = ~preissue_pkt_o[29];
  assign N251 = ~preissue_pkt_o[28];
  assign N252 = ~preissue_pkt_o[27];
  assign N253 = ~preissue_pkt_o[26];
  assign N254 = ~preissue_pkt_o[25];
  assign N255 = ~preissue_pkt_o[16];
  assign N256 = ~preissue_pkt_o[14];
  assign N257 = ~preissue_pkt_o[13];
  assign N258 = ~preissue_pkt_o[12];
  assign N259 = ~preissue_pkt_o[11];
  assign N260 = ~preissue_pkt_o[10];
  assign N261 = ~preissue_pkt_o[9];
  assign N262 = ~preissue_pkt_o[8];
  assign N263 = ~preissue_pkt_o[7];
  assign N264 = ~preissue_pkt_o[6];
  assign N288 = ~preissue_pkt_o[23];
  assign N289 = ~preissue_pkt_o[22];
  assign N292 = ~preissue_pkt_o[24];
  assign N293 = ~preissue_pkt_o[23];
  assign N296 = ~preissue_pkt_o[24];
  assign N297 = ~preissue_pkt_o[23];
  assign N298 = ~preissue_pkt_o[22];
  assign N301 = ~preissue_pkt_o[24];
  assign N302 = ~preissue_pkt_o[22];
  assign N305 = N682 | N304;
  assign N682 = N681 | N300;
  assign N681 = N291 | N295;
  assign N306 = ~N305;
  assign N309 = ~N287;
  assign N312 = ~preissue_pkt_o[29];
  assign N313 = ~preissue_pkt_o[28];
  assign N314 = ~preissue_pkt_o[26];
  assign N315 = ~preissue_pkt_o[25];
  assign N316 = ~preissue_pkt_o[24];
  assign N317 = ~preissue_pkt_o[7];
  assign N318 = ~preissue_pkt_o[5];
  assign N319 = ~preissue_pkt_o[4];
  assign N332 = ~N331;
  assign N333 = ~preissue_pkt_o[31];
  assign N334 = ~preissue_pkt_o[30];
  assign N335 = ~preissue_pkt_o[27];
  assign N336 = ~preissue_pkt_o[23];
  assign N337 = ~preissue_pkt_o[22];
  assign N343 = ~preissue_pkt_o[31];
  assign N344 = ~preissue_pkt_o[30];
  assign N345 = ~preissue_pkt_o[27];
  assign N346 = ~preissue_pkt_o[23];
  assign N352 = ~preissue_pkt_o[31];
  assign N353 = ~preissue_pkt_o[30];
  assign N354 = ~preissue_pkt_o[27];
  assign N355 = ~preissue_pkt_o[22];
  assign N361 = ~preissue_pkt_o[31];
  assign N362 = ~preissue_pkt_o[30];
  assign N363 = ~preissue_pkt_o[27];
  assign N369 = ~preissue_pkt_o[31];
  assign N370 = ~preissue_pkt_o[30];
  assign N371 = ~preissue_pkt_o[23];
  assign N372 = ~preissue_pkt_o[22];
  assign N378 = ~preissue_pkt_o[31];
  assign N379 = ~preissue_pkt_o[30];
  assign N380 = ~preissue_pkt_o[23];
  assign N386 = ~preissue_pkt_o[31];
  assign N387 = ~preissue_pkt_o[30];
  assign N388 = ~preissue_pkt_o[22];
  assign N394 = ~preissue_pkt_o[31];
  assign N395 = ~preissue_pkt_o[30];
  assign N401 = ~preissue_pkt_o[33];
  assign N402 = ~preissue_pkt_o[31];
  assign N403 = ~preissue_pkt_o[30];
  assign N404 = ~preissue_pkt_o[27];
  assign N405 = ~preissue_pkt_o[23];
  assign N411 = ~preissue_pkt_o[33];
  assign N412 = ~preissue_pkt_o[31];
  assign N413 = ~preissue_pkt_o[30];
  assign N414 = ~preissue_pkt_o[23];
  assign N415 = ~preissue_pkt_o[22];
  assign N421 = ~preissue_pkt_o[30];
  assign N422 = ~preissue_pkt_o[27];
  assign N423 = ~preissue_pkt_o[23];
  assign N424 = ~preissue_pkt_o[22];
  assign N425 = ~preissue_pkt_o[16];
  assign N426 = ~preissue_pkt_o[15];
  assign N427 = ~preissue_pkt_o[14];
  assign N436 = ~preissue_pkt_o[30];
  assign N437 = ~preissue_pkt_o[23];
  assign N438 = ~preissue_pkt_o[22];
  assign N439 = ~preissue_pkt_o[16];
  assign N440 = ~preissue_pkt_o[15];
  assign N441 = ~preissue_pkt_o[14];
  assign N450 = ~preissue_pkt_o[30];
  assign N451 = ~preissue_pkt_o[27];
  assign N452 = ~preissue_pkt_o[23];
  assign N453 = ~preissue_pkt_o[22];
  assign N454 = ~preissue_pkt_o[16];
  assign N455 = ~preissue_pkt_o[15];
  assign N464 = ~preissue_pkt_o[30];
  assign N465 = ~preissue_pkt_o[23];
  assign N466 = ~preissue_pkt_o[22];
  assign N467 = ~preissue_pkt_o[16];
  assign N468 = ~preissue_pkt_o[15];
  assign N477 = N694 | N476;
  assign N694 = N693 | N463;
  assign N693 = N692 | N449;
  assign N692 = N691 | N435;
  assign N691 = N690 | N420;
  assign N690 = N689 | N410;
  assign N689 = N688 | N400;
  assign N688 = N687 | N393;
  assign N687 = N686 | N385;
  assign N686 = N685 | N377;
  assign N685 = N684 | N368;
  assign N684 = N683 | N360;
  assign N683 = N342 | N351;
  assign N478 = ~preissue_pkt_o[31];
  assign N479 = ~preissue_pkt_o[27];
  assign N480 = ~preissue_pkt_o[23];
  assign N481 = ~preissue_pkt_o[22];
  assign N487 = ~preissue_pkt_o[31];
  assign N488 = ~preissue_pkt_o[27];
  assign N489 = ~preissue_pkt_o[23];
  assign N495 = ~preissue_pkt_o[31];
  assign N496 = ~preissue_pkt_o[27];
  assign N497 = ~preissue_pkt_o[22];
  assign N503 = ~preissue_pkt_o[31];
  assign N504 = ~preissue_pkt_o[27];
  assign N510 = ~preissue_pkt_o[31];
  assign N511 = ~preissue_pkt_o[23];
  assign N512 = ~preissue_pkt_o[22];
  assign N518 = ~preissue_pkt_o[31];
  assign N519 = ~preissue_pkt_o[23];
  assign N525 = ~preissue_pkt_o[31];
  assign N526 = ~preissue_pkt_o[22];
  assign N532 = ~preissue_pkt_o[31];
  assign N538 = ~preissue_pkt_o[27];
  assign N539 = ~preissue_pkt_o[23];
  assign N540 = ~preissue_pkt_o[22];
  assign N541 = ~preissue_pkt_o[16];
  assign N542 = ~preissue_pkt_o[15];
  assign N543 = ~preissue_pkt_o[14];
  assign N552 = ~preissue_pkt_o[23];
  assign N553 = ~preissue_pkt_o[22];
  assign N554 = ~preissue_pkt_o[16];
  assign N555 = ~preissue_pkt_o[15];
  assign N556 = ~preissue_pkt_o[14];
  assign N565 = N702 | N564;
  assign N702 = N701 | N551;
  assign N701 = N700 | N537;
  assign N700 = N699 | N531;
  assign N699 = N698 | N524;
  assign N698 = N697 | N517;
  assign N697 = N696 | N509;
  assign N696 = N695 | N502;
  assign N695 = N486 | N494;
  assign N566 = ~preissue_pkt_o[33];
  assign N569 = ~preissue_pkt_o[33];
  assign N573 = ~preissue_pkt_o[33];
  assign N575 = ~preissue_pkt_o[33];
  assign N577 = ~preissue_pkt_o[33];
  assign N578 = ~preissue_pkt_o[27];
  assign N579 = ~preissue_pkt_o[22];
  assign N587 = N568 | N710;
  assign N710 = N571 | N709;
  assign N709 = N572 | N708;
  assign N708 = N574 | N707;
  assign N707 = N576 | N706;
  assign N706 = N581 | N705;
  assign N705 = N583 | N704;
  assign N704 = N584 | N703;
  assign N703 = N585 | N586;
  assign N588 = ~N587;
  assign N589 = N588;
  assign N592 = ~N565;
  assign N593 = N592;
  assign N598 = ~N234;
  assign N599 = N598;
  assign _6_net_ = ~bypass_issue;
  assign _4_net_ = N712 | enq[0];
  assign N712 = N711 | enq[1];
  assign N711 = enq[3] | enq[2];
  assign fe_queue_ready_and_o = ~full;
  assign N600 = ~issue_pkt_o[262];
  assign issue_pkt_o[263] = en_i & N713;
  assign N713 = ~empty;
  assign issue_pkt_o[262] = N621 & N714;
  assign N714 = ~illegal_instr_lo;
  assign issue_pkt_o[257] = N618 & illegal_instr_lo;

endmodule

